module NyGPU(
SREG_0,
SREG_1,
SREG_10,
SREG_11,
SREG_12,
SREG_13,
SREG_14,
SREG_15,
SREG_16,
SREG_17,
SREG_18,
SREG_19,
SREG_2,
SREG_20,
SREG_21,
SREG_22,
SREG_23,
SREG_24,
SREG_25,
SREG_26,
SREG_27,
SREG_28,
SREG_29,
SREG_3,
SREG_30,
SREG_31,
SREG_4,
SREG_5,
SREG_6,
SREG_7,
SREG_8,
SREG_9,
VREG_0_0,
VREG_0_1,
VREG_0_10,
VREG_0_11,
VREG_0_12,
VREG_0_13,
VREG_0_14,
VREG_0_15,
VREG_0_2,
VREG_0_3,
VREG_0_4,
VREG_0_5,
VREG_0_6,
VREG_0_7,
VREG_0_8,
VREG_0_9,
VREG_10_0,
VREG_10_1,
VREG_10_10,
VREG_10_11,
VREG_10_12,
VREG_10_13,
VREG_10_14,
VREG_10_15,
VREG_10_2,
VREG_10_3,
VREG_10_4,
VREG_10_5,
VREG_10_6,
VREG_10_7,
VREG_10_8,
VREG_10_9,
VREG_11_0,
VREG_11_1,
VREG_11_10,
VREG_11_11,
VREG_11_12,
VREG_11_13,
VREG_11_14,
VREG_11_15,
VREG_11_2,
VREG_11_3,
VREG_11_4,
VREG_11_5,
VREG_11_6,
VREG_11_7,
VREG_11_8,
VREG_11_9,
VREG_12_0,
VREG_12_1,
VREG_12_10,
VREG_12_11,
VREG_12_12,
VREG_12_13,
VREG_12_14,
VREG_12_15,
VREG_12_2,
VREG_12_3,
VREG_12_4,
VREG_12_5,
VREG_12_6,
VREG_12_7,
VREG_12_8,
VREG_12_9,
VREG_13_0,
VREG_13_1,
VREG_13_10,
VREG_13_11,
VREG_13_12,
VREG_13_13,
VREG_13_14,
VREG_13_15,
VREG_13_2,
VREG_13_3,
VREG_13_4,
VREG_13_5,
VREG_13_6,
VREG_13_7,
VREG_13_8,
VREG_13_9,
VREG_14_0,
VREG_14_1,
VREG_14_10,
VREG_14_11,
VREG_14_12,
VREG_14_13,
VREG_14_14,
VREG_14_15,
VREG_14_2,
VREG_14_3,
VREG_14_4,
VREG_14_5,
VREG_14_6,
VREG_14_7,
VREG_14_8,
VREG_14_9,
VREG_15_0,
VREG_15_1,
VREG_15_10,
VREG_15_11,
VREG_15_12,
VREG_15_13,
VREG_15_14,
VREG_15_15,
VREG_15_2,
VREG_15_3,
VREG_15_4,
VREG_15_5,
VREG_15_6,
VREG_15_7,
VREG_15_8,
VREG_15_9,
VREG_16_0,
VREG_16_1,
VREG_16_10,
VREG_16_11,
VREG_16_12,
VREG_16_13,
VREG_16_14,
VREG_16_15,
VREG_16_2,
VREG_16_3,
VREG_16_4,
VREG_16_5,
VREG_16_6,
VREG_16_7,
VREG_16_8,
VREG_16_9,
VREG_17_0,
VREG_17_1,
VREG_17_10,
VREG_17_11,
VREG_17_12,
VREG_17_13,
VREG_17_14,
VREG_17_15,
VREG_17_2,
VREG_17_3,
VREG_17_4,
VREG_17_5,
VREG_17_6,
VREG_17_7,
VREG_17_8,
VREG_17_9,
VREG_18_0,
VREG_18_1,
VREG_18_10,
VREG_18_11,
VREG_18_12,
VREG_18_13,
VREG_18_14,
VREG_18_15,
VREG_18_2,
VREG_18_3,
VREG_18_4,
VREG_18_5,
VREG_18_6,
VREG_18_7,
VREG_18_8,
VREG_18_9,
VREG_19_0,
VREG_19_1,
VREG_19_10,
VREG_19_11,
VREG_19_12,
VREG_19_13,
VREG_19_14,
VREG_19_15,
VREG_19_2,
VREG_19_3,
VREG_19_4,
VREG_19_5,
VREG_19_6,
VREG_19_7,
VREG_19_8,
VREG_19_9,
VREG_1_0,
VREG_1_1,
VREG_1_10,
VREG_1_11,
VREG_1_12,
VREG_1_13,
VREG_1_14,
VREG_1_15,
VREG_1_2,
VREG_1_3,
VREG_1_4,
VREG_1_5,
VREG_1_6,
VREG_1_7,
VREG_1_8,
VREG_1_9,
VREG_20_0,
VREG_20_1,
VREG_20_10,
VREG_20_11,
VREG_20_12,
VREG_20_13,
VREG_20_14,
VREG_20_15,
VREG_20_2,
VREG_20_3,
VREG_20_4,
VREG_20_5,
VREG_20_6,
VREG_20_7,
VREG_20_8,
VREG_20_9,
VREG_21_0,
VREG_21_1,
VREG_21_10,
VREG_21_11,
VREG_21_12,
VREG_21_13,
VREG_21_14,
VREG_21_15,
VREG_21_2,
VREG_21_3,
VREG_21_4,
VREG_21_5,
VREG_21_6,
VREG_21_7,
VREG_21_8,
VREG_21_9,
VREG_22_0,
VREG_22_1,
VREG_22_10,
VREG_22_11,
VREG_22_12,
VREG_22_13,
VREG_22_14,
VREG_22_15,
VREG_22_2,
VREG_22_3,
VREG_22_4,
VREG_22_5,
VREG_22_6,
VREG_22_7,
VREG_22_8,
VREG_22_9,
VREG_23_0,
VREG_23_1,
VREG_23_10,
VREG_23_11,
VREG_23_12,
VREG_23_13,
VREG_23_14,
VREG_23_15,
VREG_23_2,
VREG_23_3,
VREG_23_4,
VREG_23_5,
VREG_23_6,
VREG_23_7,
VREG_23_8,
VREG_23_9,
VREG_24_0,
VREG_24_1,
VREG_24_10,
VREG_24_11,
VREG_24_12,
VREG_24_13,
VREG_24_14,
VREG_24_15,
VREG_24_2,
VREG_24_3,
VREG_24_4,
VREG_24_5,
VREG_24_6,
VREG_24_7,
VREG_24_8,
VREG_24_9,
VREG_25_0,
VREG_25_1,
VREG_25_10,
VREG_25_11,
VREG_25_12,
VREG_25_13,
VREG_25_14,
VREG_25_15,
VREG_25_2,
VREG_25_3,
VREG_25_4,
VREG_25_5,
VREG_25_6,
VREG_25_7,
VREG_25_8,
VREG_25_9,
VREG_26_0,
VREG_26_1,
VREG_26_10,
VREG_26_11,
VREG_26_12,
VREG_26_13,
VREG_26_14,
VREG_26_15,
VREG_26_2,
VREG_26_3,
VREG_26_4,
VREG_26_5,
VREG_26_6,
VREG_26_7,
VREG_26_8,
VREG_26_9,
VREG_27_0,
VREG_27_1,
VREG_27_10,
VREG_27_11,
VREG_27_12,
VREG_27_13,
VREG_27_14,
VREG_27_15,
VREG_27_2,
VREG_27_3,
VREG_27_4,
VREG_27_5,
VREG_27_6,
VREG_27_7,
VREG_27_8,
VREG_27_9,
VREG_28_0,
VREG_28_1,
VREG_28_10,
VREG_28_11,
VREG_28_12,
VREG_28_13,
VREG_28_14,
VREG_28_15,
VREG_28_2,
VREG_28_3,
VREG_28_4,
VREG_28_5,
VREG_28_6,
VREG_28_7,
VREG_28_8,
VREG_28_9,
VREG_29_0,
VREG_29_1,
VREG_29_10,
VREG_29_11,
VREG_29_12,
VREG_29_13,
VREG_29_14,
VREG_29_15,
VREG_29_2,
VREG_29_3,
VREG_29_4,
VREG_29_5,
VREG_29_6,
VREG_29_7,
VREG_29_8,
VREG_29_9,
VREG_2_0,
VREG_2_1,
VREG_2_10,
VREG_2_11,
VREG_2_12,
VREG_2_13,
VREG_2_14,
VREG_2_15,
VREG_2_2,
VREG_2_3,
VREG_2_4,
VREG_2_5,
VREG_2_6,
VREG_2_7,
VREG_2_8,
VREG_2_9,
VREG_30_0,
VREG_30_1,
VREG_30_10,
VREG_30_11,
VREG_30_12,
VREG_30_13,
VREG_30_14,
VREG_30_15,
VREG_30_2,
VREG_30_3,
VREG_30_4,
VREG_30_5,
VREG_30_6,
VREG_30_7,
VREG_30_8,
VREG_30_9,
VREG_31_0,
VREG_31_1,
VREG_31_10,
VREG_31_11,
VREG_31_12,
VREG_31_13,
VREG_31_14,
VREG_31_15,
VREG_31_2,
VREG_31_3,
VREG_31_4,
VREG_31_5,
VREG_31_6,
VREG_31_7,
VREG_31_8,
VREG_31_9,
VREG_3_0,
VREG_3_1,
VREG_3_10,
VREG_3_11,
VREG_3_12,
VREG_3_13,
VREG_3_14,
VREG_3_15,
VREG_3_2,
VREG_3_3,
VREG_3_4,
VREG_3_5,
VREG_3_6,
VREG_3_7,
VREG_3_8,
VREG_3_9,
VREG_4_0,
VREG_4_1,
VREG_4_10,
VREG_4_11,
VREG_4_12,
VREG_4_13,
VREG_4_14,
VREG_4_15,
VREG_4_2,
VREG_4_3,
VREG_4_4,
VREG_4_5,
VREG_4_6,
VREG_4_7,
VREG_4_8,
VREG_4_9,
VREG_5_0,
VREG_5_1,
VREG_5_10,
VREG_5_11,
VREG_5_12,
VREG_5_13,
VREG_5_14,
VREG_5_15,
VREG_5_2,
VREG_5_3,
VREG_5_4,
VREG_5_5,
VREG_5_6,
VREG_5_7,
VREG_5_8,
VREG_5_9,
VREG_6_0,
VREG_6_1,
VREG_6_10,
VREG_6_11,
VREG_6_12,
VREG_6_13,
VREG_6_14,
VREG_6_15,
VREG_6_2,
VREG_6_3,
VREG_6_4,
VREG_6_5,
VREG_6_6,
VREG_6_7,
VREG_6_8,
VREG_6_9,
VREG_7_0,
VREG_7_1,
VREG_7_10,
VREG_7_11,
VREG_7_12,
VREG_7_13,
VREG_7_14,
VREG_7_15,
VREG_7_2,
VREG_7_3,
VREG_7_4,
VREG_7_5,
VREG_7_6,
VREG_7_7,
VREG_7_8,
VREG_7_9,
VREG_8_0,
VREG_8_1,
VREG_8_10,
VREG_8_11,
VREG_8_12,
VREG_8_13,
VREG_8_14,
VREG_8_15,
VREG_8_2,
VREG_8_3,
VREG_8_4,
VREG_8_5,
VREG_8_6,
VREG_8_7,
VREG_8_8,
VREG_8_9,
VREG_9_0,
VREG_9_1,
VREG_9_10,
VREG_9_11,
VREG_9_12,
VREG_9_13,
VREG_9_14,
VREG_9_15,
VREG_9_2,
VREG_9_3,
VREG_9_4,
VREG_9_5,
VREG_9_6,
VREG_9_7,
VREG_9_8,
VREG_9_9,
imem_raddr_ila,
imem_rdata_ila,
pc,
vector_mask_register,
clk,rst,
step
);
input clk;
input rst;
input step;
input [31:0] imem_rdata_ila;
output [31:0] imem_raddr_ila;
output     [31:0] SREG_0;
output     [31:0] SREG_1;
output     [31:0] SREG_10;
output     [31:0] SREG_11;
output     [31:0] SREG_12;
output     [31:0] SREG_13;
output     [31:0] SREG_14;
output     [31:0] SREG_15;
output     [31:0] SREG_16;
output     [31:0] SREG_17;
output     [31:0] SREG_18;
output     [31:0] SREG_19;
output     [31:0] SREG_2;
output     [31:0] SREG_20;
output     [31:0] SREG_21;
output     [31:0] SREG_22;
output     [31:0] SREG_23;
output     [31:0] SREG_24;
output     [31:0] SREG_25;
output     [31:0] SREG_26;
output     [31:0] SREG_27;
output     [31:0] SREG_28;
output     [31:0] SREG_29;
output     [31:0] SREG_3;
output     [31:0] SREG_30;
output     [31:0] SREG_31;
output     [31:0] SREG_4;
output     [31:0] SREG_5;
output     [31:0] SREG_6;
output     [31:0] SREG_7;
output     [31:0] SREG_8;
output     [31:0] SREG_9;
output     [31:0] VREG_0_0;
output     [31:0] VREG_0_1;
output     [31:0] VREG_0_10;
output     [31:0] VREG_0_11;
output     [31:0] VREG_0_12;
output     [31:0] VREG_0_13;
output     [31:0] VREG_0_14;
output     [31:0] VREG_0_15;
output     [31:0] VREG_0_2;
output     [31:0] VREG_0_3;
output     [31:0] VREG_0_4;
output     [31:0] VREG_0_5;
output     [31:0] VREG_0_6;
output     [31:0] VREG_0_7;
output     [31:0] VREG_0_8;
output     [31:0] VREG_0_9;
output     [31:0] VREG_10_0;
output     [31:0] VREG_10_1;
output     [31:0] VREG_10_10;
output     [31:0] VREG_10_11;
output     [31:0] VREG_10_12;
output     [31:0] VREG_10_13;
output     [31:0] VREG_10_14;
output     [31:0] VREG_10_15;
output     [31:0] VREG_10_2;
output     [31:0] VREG_10_3;
output     [31:0] VREG_10_4;
output     [31:0] VREG_10_5;
output     [31:0] VREG_10_6;
output     [31:0] VREG_10_7;
output     [31:0] VREG_10_8;
output     [31:0] VREG_10_9;
output     [31:0] VREG_11_0;
output     [31:0] VREG_11_1;
output     [31:0] VREG_11_10;
output     [31:0] VREG_11_11;
output     [31:0] VREG_11_12;
output     [31:0] VREG_11_13;
output     [31:0] VREG_11_14;
output     [31:0] VREG_11_15;
output     [31:0] VREG_11_2;
output     [31:0] VREG_11_3;
output     [31:0] VREG_11_4;
output     [31:0] VREG_11_5;
output     [31:0] VREG_11_6;
output     [31:0] VREG_11_7;
output     [31:0] VREG_11_8;
output     [31:0] VREG_11_9;
output     [31:0] VREG_12_0;
output     [31:0] VREG_12_1;
output     [31:0] VREG_12_10;
output     [31:0] VREG_12_11;
output     [31:0] VREG_12_12;
output     [31:0] VREG_12_13;
output     [31:0] VREG_12_14;
output     [31:0] VREG_12_15;
output     [31:0] VREG_12_2;
output     [31:0] VREG_12_3;
output     [31:0] VREG_12_4;
output     [31:0] VREG_12_5;
output     [31:0] VREG_12_6;
output     [31:0] VREG_12_7;
output     [31:0] VREG_12_8;
output     [31:0] VREG_12_9;
output     [31:0] VREG_13_0;
output     [31:0] VREG_13_1;
output     [31:0] VREG_13_10;
output     [31:0] VREG_13_11;
output     [31:0] VREG_13_12;
output     [31:0] VREG_13_13;
output     [31:0] VREG_13_14;
output     [31:0] VREG_13_15;
output     [31:0] VREG_13_2;
output     [31:0] VREG_13_3;
output     [31:0] VREG_13_4;
output     [31:0] VREG_13_5;
output     [31:0] VREG_13_6;
output     [31:0] VREG_13_7;
output     [31:0] VREG_13_8;
output     [31:0] VREG_13_9;
output     [31:0] VREG_14_0;
output     [31:0] VREG_14_1;
output     [31:0] VREG_14_10;
output     [31:0] VREG_14_11;
output     [31:0] VREG_14_12;
output     [31:0] VREG_14_13;
output     [31:0] VREG_14_14;
output     [31:0] VREG_14_15;
output     [31:0] VREG_14_2;
output     [31:0] VREG_14_3;
output     [31:0] VREG_14_4;
output     [31:0] VREG_14_5;
output     [31:0] VREG_14_6;
output     [31:0] VREG_14_7;
output     [31:0] VREG_14_8;
output     [31:0] VREG_14_9;
output     [31:0] VREG_15_0;
output     [31:0] VREG_15_1;
output     [31:0] VREG_15_10;
output     [31:0] VREG_15_11;
output     [31:0] VREG_15_12;
output     [31:0] VREG_15_13;
output     [31:0] VREG_15_14;
output     [31:0] VREG_15_15;
output     [31:0] VREG_15_2;
output     [31:0] VREG_15_3;
output     [31:0] VREG_15_4;
output     [31:0] VREG_15_5;
output     [31:0] VREG_15_6;
output     [31:0] VREG_15_7;
output     [31:0] VREG_15_8;
output     [31:0] VREG_15_9;
output     [31:0] VREG_16_0;
output     [31:0] VREG_16_1;
output     [31:0] VREG_16_10;
output     [31:0] VREG_16_11;
output     [31:0] VREG_16_12;
output     [31:0] VREG_16_13;
output     [31:0] VREG_16_14;
output     [31:0] VREG_16_15;
output     [31:0] VREG_16_2;
output     [31:0] VREG_16_3;
output     [31:0] VREG_16_4;
output     [31:0] VREG_16_5;
output     [31:0] VREG_16_6;
output     [31:0] VREG_16_7;
output     [31:0] VREG_16_8;
output     [31:0] VREG_16_9;
output     [31:0] VREG_17_0;
output     [31:0] VREG_17_1;
output     [31:0] VREG_17_10;
output     [31:0] VREG_17_11;
output     [31:0] VREG_17_12;
output     [31:0] VREG_17_13;
output     [31:0] VREG_17_14;
output     [31:0] VREG_17_15;
output     [31:0] VREG_17_2;
output     [31:0] VREG_17_3;
output     [31:0] VREG_17_4;
output     [31:0] VREG_17_5;
output     [31:0] VREG_17_6;
output     [31:0] VREG_17_7;
output     [31:0] VREG_17_8;
output     [31:0] VREG_17_9;
output     [31:0] VREG_18_0;
output     [31:0] VREG_18_1;
output     [31:0] VREG_18_10;
output     [31:0] VREG_18_11;
output     [31:0] VREG_18_12;
output     [31:0] VREG_18_13;
output     [31:0] VREG_18_14;
output     [31:0] VREG_18_15;
output     [31:0] VREG_18_2;
output     [31:0] VREG_18_3;
output     [31:0] VREG_18_4;
output     [31:0] VREG_18_5;
output     [31:0] VREG_18_6;
output     [31:0] VREG_18_7;
output     [31:0] VREG_18_8;
output     [31:0] VREG_18_9;
output     [31:0] VREG_19_0;
output     [31:0] VREG_19_1;
output     [31:0] VREG_19_10;
output     [31:0] VREG_19_11;
output     [31:0] VREG_19_12;
output     [31:0] VREG_19_13;
output     [31:0] VREG_19_14;
output     [31:0] VREG_19_15;
output     [31:0] VREG_19_2;
output     [31:0] VREG_19_3;
output     [31:0] VREG_19_4;
output     [31:0] VREG_19_5;
output     [31:0] VREG_19_6;
output     [31:0] VREG_19_7;
output     [31:0] VREG_19_8;
output     [31:0] VREG_19_9;
output     [31:0] VREG_1_0;
output     [31:0] VREG_1_1;
output     [31:0] VREG_1_10;
output     [31:0] VREG_1_11;
output     [31:0] VREG_1_12;
output     [31:0] VREG_1_13;
output     [31:0] VREG_1_14;
output     [31:0] VREG_1_15;
output     [31:0] VREG_1_2;
output     [31:0] VREG_1_3;
output     [31:0] VREG_1_4;
output     [31:0] VREG_1_5;
output     [31:0] VREG_1_6;
output     [31:0] VREG_1_7;
output     [31:0] VREG_1_8;
output     [31:0] VREG_1_9;
output     [31:0] VREG_20_0;
output     [31:0] VREG_20_1;
output     [31:0] VREG_20_10;
output     [31:0] VREG_20_11;
output     [31:0] VREG_20_12;
output     [31:0] VREG_20_13;
output     [31:0] VREG_20_14;
output     [31:0] VREG_20_15;
output     [31:0] VREG_20_2;
output     [31:0] VREG_20_3;
output     [31:0] VREG_20_4;
output     [31:0] VREG_20_5;
output     [31:0] VREG_20_6;
output     [31:0] VREG_20_7;
output     [31:0] VREG_20_8;
output     [31:0] VREG_20_9;
output     [31:0] VREG_21_0;
output     [31:0] VREG_21_1;
output     [31:0] VREG_21_10;
output     [31:0] VREG_21_11;
output     [31:0] VREG_21_12;
output     [31:0] VREG_21_13;
output     [31:0] VREG_21_14;
output     [31:0] VREG_21_15;
output     [31:0] VREG_21_2;
output     [31:0] VREG_21_3;
output     [31:0] VREG_21_4;
output     [31:0] VREG_21_5;
output     [31:0] VREG_21_6;
output     [31:0] VREG_21_7;
output     [31:0] VREG_21_8;
output     [31:0] VREG_21_9;
output     [31:0] VREG_22_0;
output     [31:0] VREG_22_1;
output     [31:0] VREG_22_10;
output     [31:0] VREG_22_11;
output     [31:0] VREG_22_12;
output     [31:0] VREG_22_13;
output     [31:0] VREG_22_14;
output     [31:0] VREG_22_15;
output     [31:0] VREG_22_2;
output     [31:0] VREG_22_3;
output     [31:0] VREG_22_4;
output     [31:0] VREG_22_5;
output     [31:0] VREG_22_6;
output     [31:0] VREG_22_7;
output     [31:0] VREG_22_8;
output     [31:0] VREG_22_9;
output     [31:0] VREG_23_0;
output     [31:0] VREG_23_1;
output     [31:0] VREG_23_10;
output     [31:0] VREG_23_11;
output     [31:0] VREG_23_12;
output     [31:0] VREG_23_13;
output     [31:0] VREG_23_14;
output     [31:0] VREG_23_15;
output     [31:0] VREG_23_2;
output     [31:0] VREG_23_3;
output     [31:0] VREG_23_4;
output     [31:0] VREG_23_5;
output     [31:0] VREG_23_6;
output     [31:0] VREG_23_7;
output     [31:0] VREG_23_8;
output     [31:0] VREG_23_9;
output     [31:0] VREG_24_0;
output     [31:0] VREG_24_1;
output     [31:0] VREG_24_10;
output     [31:0] VREG_24_11;
output     [31:0] VREG_24_12;
output     [31:0] VREG_24_13;
output     [31:0] VREG_24_14;
output     [31:0] VREG_24_15;
output     [31:0] VREG_24_2;
output     [31:0] VREG_24_3;
output     [31:0] VREG_24_4;
output     [31:0] VREG_24_5;
output     [31:0] VREG_24_6;
output     [31:0] VREG_24_7;
output     [31:0] VREG_24_8;
output     [31:0] VREG_24_9;
output     [31:0] VREG_25_0;
output     [31:0] VREG_25_1;
output     [31:0] VREG_25_10;
output     [31:0] VREG_25_11;
output     [31:0] VREG_25_12;
output     [31:0] VREG_25_13;
output     [31:0] VREG_25_14;
output     [31:0] VREG_25_15;
output     [31:0] VREG_25_2;
output     [31:0] VREG_25_3;
output     [31:0] VREG_25_4;
output     [31:0] VREG_25_5;
output     [31:0] VREG_25_6;
output     [31:0] VREG_25_7;
output     [31:0] VREG_25_8;
output     [31:0] VREG_25_9;
output     [31:0] VREG_26_0;
output     [31:0] VREG_26_1;
output     [31:0] VREG_26_10;
output     [31:0] VREG_26_11;
output     [31:0] VREG_26_12;
output     [31:0] VREG_26_13;
output     [31:0] VREG_26_14;
output     [31:0] VREG_26_15;
output     [31:0] VREG_26_2;
output     [31:0] VREG_26_3;
output     [31:0] VREG_26_4;
output     [31:0] VREG_26_5;
output     [31:0] VREG_26_6;
output     [31:0] VREG_26_7;
output     [31:0] VREG_26_8;
output     [31:0] VREG_26_9;
output     [31:0] VREG_27_0;
output     [31:0] VREG_27_1;
output     [31:0] VREG_27_10;
output     [31:0] VREG_27_11;
output     [31:0] VREG_27_12;
output     [31:0] VREG_27_13;
output     [31:0] VREG_27_14;
output     [31:0] VREG_27_15;
output     [31:0] VREG_27_2;
output     [31:0] VREG_27_3;
output     [31:0] VREG_27_4;
output     [31:0] VREG_27_5;
output     [31:0] VREG_27_6;
output     [31:0] VREG_27_7;
output     [31:0] VREG_27_8;
output     [31:0] VREG_27_9;
output     [31:0] VREG_28_0;
output     [31:0] VREG_28_1;
output     [31:0] VREG_28_10;
output     [31:0] VREG_28_11;
output     [31:0] VREG_28_12;
output     [31:0] VREG_28_13;
output     [31:0] VREG_28_14;
output     [31:0] VREG_28_15;
output     [31:0] VREG_28_2;
output     [31:0] VREG_28_3;
output     [31:0] VREG_28_4;
output     [31:0] VREG_28_5;
output     [31:0] VREG_28_6;
output     [31:0] VREG_28_7;
output     [31:0] VREG_28_8;
output     [31:0] VREG_28_9;
output     [31:0] VREG_29_0;
output     [31:0] VREG_29_1;
output     [31:0] VREG_29_10;
output     [31:0] VREG_29_11;
output     [31:0] VREG_29_12;
output     [31:0] VREG_29_13;
output     [31:0] VREG_29_14;
output     [31:0] VREG_29_15;
output     [31:0] VREG_29_2;
output     [31:0] VREG_29_3;
output     [31:0] VREG_29_4;
output     [31:0] VREG_29_5;
output     [31:0] VREG_29_6;
output     [31:0] VREG_29_7;
output     [31:0] VREG_29_8;
output     [31:0] VREG_29_9;
output     [31:0] VREG_2_0;
output     [31:0] VREG_2_1;
output     [31:0] VREG_2_10;
output     [31:0] VREG_2_11;
output     [31:0] VREG_2_12;
output     [31:0] VREG_2_13;
output     [31:0] VREG_2_14;
output     [31:0] VREG_2_15;
output     [31:0] VREG_2_2;
output     [31:0] VREG_2_3;
output     [31:0] VREG_2_4;
output     [31:0] VREG_2_5;
output     [31:0] VREG_2_6;
output     [31:0] VREG_2_7;
output     [31:0] VREG_2_8;
output     [31:0] VREG_2_9;
output     [31:0] VREG_30_0;
output     [31:0] VREG_30_1;
output     [31:0] VREG_30_10;
output     [31:0] VREG_30_11;
output     [31:0] VREG_30_12;
output     [31:0] VREG_30_13;
output     [31:0] VREG_30_14;
output     [31:0] VREG_30_15;
output     [31:0] VREG_30_2;
output     [31:0] VREG_30_3;
output     [31:0] VREG_30_4;
output     [31:0] VREG_30_5;
output     [31:0] VREG_30_6;
output     [31:0] VREG_30_7;
output     [31:0] VREG_30_8;
output     [31:0] VREG_30_9;
output     [31:0] VREG_31_0;
output     [31:0] VREG_31_1;
output     [31:0] VREG_31_10;
output     [31:0] VREG_31_11;
output     [31:0] VREG_31_12;
output     [31:0] VREG_31_13;
output     [31:0] VREG_31_14;
output     [31:0] VREG_31_15;
output     [31:0] VREG_31_2;
output     [31:0] VREG_31_3;
output     [31:0] VREG_31_4;
output     [31:0] VREG_31_5;
output     [31:0] VREG_31_6;
output     [31:0] VREG_31_7;
output     [31:0] VREG_31_8;
output     [31:0] VREG_31_9;
output     [31:0] VREG_3_0;
output     [31:0] VREG_3_1;
output     [31:0] VREG_3_10;
output     [31:0] VREG_3_11;
output     [31:0] VREG_3_12;
output     [31:0] VREG_3_13;
output     [31:0] VREG_3_14;
output     [31:0] VREG_3_15;
output     [31:0] VREG_3_2;
output     [31:0] VREG_3_3;
output     [31:0] VREG_3_4;
output     [31:0] VREG_3_5;
output     [31:0] VREG_3_6;
output     [31:0] VREG_3_7;
output     [31:0] VREG_3_8;
output     [31:0] VREG_3_9;
output     [31:0] VREG_4_0;
output     [31:0] VREG_4_1;
output     [31:0] VREG_4_10;
output     [31:0] VREG_4_11;
output     [31:0] VREG_4_12;
output     [31:0] VREG_4_13;
output     [31:0] VREG_4_14;
output     [31:0] VREG_4_15;
output     [31:0] VREG_4_2;
output     [31:0] VREG_4_3;
output     [31:0] VREG_4_4;
output     [31:0] VREG_4_5;
output     [31:0] VREG_4_6;
output     [31:0] VREG_4_7;
output     [31:0] VREG_4_8;
output     [31:0] VREG_4_9;
output     [31:0] VREG_5_0;
output     [31:0] VREG_5_1;
output     [31:0] VREG_5_10;
output     [31:0] VREG_5_11;
output     [31:0] VREG_5_12;
output     [31:0] VREG_5_13;
output     [31:0] VREG_5_14;
output     [31:0] VREG_5_15;
output     [31:0] VREG_5_2;
output     [31:0] VREG_5_3;
output     [31:0] VREG_5_4;
output     [31:0] VREG_5_5;
output     [31:0] VREG_5_6;
output     [31:0] VREG_5_7;
output     [31:0] VREG_5_8;
output     [31:0] VREG_5_9;
output     [31:0] VREG_6_0;
output     [31:0] VREG_6_1;
output     [31:0] VREG_6_10;
output     [31:0] VREG_6_11;
output     [31:0] VREG_6_12;
output     [31:0] VREG_6_13;
output     [31:0] VREG_6_14;
output     [31:0] VREG_6_15;
output     [31:0] VREG_6_2;
output     [31:0] VREG_6_3;
output     [31:0] VREG_6_4;
output     [31:0] VREG_6_5;
output     [31:0] VREG_6_6;
output     [31:0] VREG_6_7;
output     [31:0] VREG_6_8;
output     [31:0] VREG_6_9;
output     [31:0] VREG_7_0;
output     [31:0] VREG_7_1;
output     [31:0] VREG_7_10;
output     [31:0] VREG_7_11;
output     [31:0] VREG_7_12;
output     [31:0] VREG_7_13;
output     [31:0] VREG_7_14;
output     [31:0] VREG_7_15;
output     [31:0] VREG_7_2;
output     [31:0] VREG_7_3;
output     [31:0] VREG_7_4;
output     [31:0] VREG_7_5;
output     [31:0] VREG_7_6;
output     [31:0] VREG_7_7;
output     [31:0] VREG_7_8;
output     [31:0] VREG_7_9;
output     [31:0] VREG_8_0;
output     [31:0] VREG_8_1;
output     [31:0] VREG_8_10;
output     [31:0] VREG_8_11;
output     [31:0] VREG_8_12;
output     [31:0] VREG_8_13;
output     [31:0] VREG_8_14;
output     [31:0] VREG_8_15;
output     [31:0] VREG_8_2;
output     [31:0] VREG_8_3;
output     [31:0] VREG_8_4;
output     [31:0] VREG_8_5;
output     [31:0] VREG_8_6;
output     [31:0] VREG_8_7;
output     [31:0] VREG_8_8;
output     [31:0] VREG_8_9;
output     [31:0] VREG_9_0;
output     [31:0] VREG_9_1;
output     [31:0] VREG_9_10;
output     [31:0] VREG_9_11;
output     [31:0] VREG_9_12;
output     [31:0] VREG_9_13;
output     [31:0] VREG_9_14;
output     [31:0] VREG_9_15;
output     [31:0] VREG_9_2;
output     [31:0] VREG_9_3;
output     [31:0] VREG_9_4;
output     [31:0] VREG_9_5;
output     [31:0] VREG_9_6;
output     [31:0] VREG_9_7;
output     [31:0] VREG_9_8;
output     [31:0] VREG_9_9;
output     [31:0] pc;
output     [31:0] vector_mask_register;
reg     [31:0] SREG_0;
reg     [31:0] SREG_1;
reg     [31:0] SREG_10;
reg     [31:0] SREG_11;
reg     [31:0] SREG_12;
reg     [31:0] SREG_13;
reg     [31:0] SREG_14;
reg     [31:0] SREG_15;
reg     [31:0] SREG_16;
reg     [31:0] SREG_17;
reg     [31:0] SREG_18;
reg     [31:0] SREG_19;
reg     [31:0] SREG_2;
reg     [31:0] SREG_20;
reg     [31:0] SREG_21;
reg     [31:0] SREG_22;
reg     [31:0] SREG_23;
reg     [31:0] SREG_24;
reg     [31:0] SREG_25;
reg     [31:0] SREG_26;
reg     [31:0] SREG_27;
reg     [31:0] SREG_28;
reg     [31:0] SREG_29;
reg     [31:0] SREG_3;
reg     [31:0] SREG_30;
reg     [31:0] SREG_31;
reg     [31:0] SREG_4;
reg     [31:0] SREG_5;
reg     [31:0] SREG_6;
reg     [31:0] SREG_7;
reg     [31:0] SREG_8;
reg     [31:0] SREG_9;
reg     [31:0] VREG_0_0;
reg     [31:0] VREG_0_1;
reg     [31:0] VREG_0_10;
reg     [31:0] VREG_0_11;
reg     [31:0] VREG_0_12;
reg     [31:0] VREG_0_13;
reg     [31:0] VREG_0_14;
reg     [31:0] VREG_0_15;
reg     [31:0] VREG_0_2;
reg     [31:0] VREG_0_3;
reg     [31:0] VREG_0_4;
reg     [31:0] VREG_0_5;
reg     [31:0] VREG_0_6;
reg     [31:0] VREG_0_7;
reg     [31:0] VREG_0_8;
reg     [31:0] VREG_0_9;
reg     [31:0] VREG_10_0;
reg     [31:0] VREG_10_1;
reg     [31:0] VREG_10_10;
reg     [31:0] VREG_10_11;
reg     [31:0] VREG_10_12;
reg     [31:0] VREG_10_13;
reg     [31:0] VREG_10_14;
reg     [31:0] VREG_10_15;
reg     [31:0] VREG_10_2;
reg     [31:0] VREG_10_3;
reg     [31:0] VREG_10_4;
reg     [31:0] VREG_10_5;
reg     [31:0] VREG_10_6;
reg     [31:0] VREG_10_7;
reg     [31:0] VREG_10_8;
reg     [31:0] VREG_10_9;
reg     [31:0] VREG_11_0;
reg     [31:0] VREG_11_1;
reg     [31:0] VREG_11_10;
reg     [31:0] VREG_11_11;
reg     [31:0] VREG_11_12;
reg     [31:0] VREG_11_13;
reg     [31:0] VREG_11_14;
reg     [31:0] VREG_11_15;
reg     [31:0] VREG_11_2;
reg     [31:0] VREG_11_3;
reg     [31:0] VREG_11_4;
reg     [31:0] VREG_11_5;
reg     [31:0] VREG_11_6;
reg     [31:0] VREG_11_7;
reg     [31:0] VREG_11_8;
reg     [31:0] VREG_11_9;
reg     [31:0] VREG_12_0;
reg     [31:0] VREG_12_1;
reg     [31:0] VREG_12_10;
reg     [31:0] VREG_12_11;
reg     [31:0] VREG_12_12;
reg     [31:0] VREG_12_13;
reg     [31:0] VREG_12_14;
reg     [31:0] VREG_12_15;
reg     [31:0] VREG_12_2;
reg     [31:0] VREG_12_3;
reg     [31:0] VREG_12_4;
reg     [31:0] VREG_12_5;
reg     [31:0] VREG_12_6;
reg     [31:0] VREG_12_7;
reg     [31:0] VREG_12_8;
reg     [31:0] VREG_12_9;
reg     [31:0] VREG_13_0;
reg     [31:0] VREG_13_1;
reg     [31:0] VREG_13_10;
reg     [31:0] VREG_13_11;
reg     [31:0] VREG_13_12;
reg     [31:0] VREG_13_13;
reg     [31:0] VREG_13_14;
reg     [31:0] VREG_13_15;
reg     [31:0] VREG_13_2;
reg     [31:0] VREG_13_3;
reg     [31:0] VREG_13_4;
reg     [31:0] VREG_13_5;
reg     [31:0] VREG_13_6;
reg     [31:0] VREG_13_7;
reg     [31:0] VREG_13_8;
reg     [31:0] VREG_13_9;
reg     [31:0] VREG_14_0;
reg     [31:0] VREG_14_1;
reg     [31:0] VREG_14_10;
reg     [31:0] VREG_14_11;
reg     [31:0] VREG_14_12;
reg     [31:0] VREG_14_13;
reg     [31:0] VREG_14_14;
reg     [31:0] VREG_14_15;
reg     [31:0] VREG_14_2;
reg     [31:0] VREG_14_3;
reg     [31:0] VREG_14_4;
reg     [31:0] VREG_14_5;
reg     [31:0] VREG_14_6;
reg     [31:0] VREG_14_7;
reg     [31:0] VREG_14_8;
reg     [31:0] VREG_14_9;
reg     [31:0] VREG_15_0;
reg     [31:0] VREG_15_1;
reg     [31:0] VREG_15_10;
reg     [31:0] VREG_15_11;
reg     [31:0] VREG_15_12;
reg     [31:0] VREG_15_13;
reg     [31:0] VREG_15_14;
reg     [31:0] VREG_15_15;
reg     [31:0] VREG_15_2;
reg     [31:0] VREG_15_3;
reg     [31:0] VREG_15_4;
reg     [31:0] VREG_15_5;
reg     [31:0] VREG_15_6;
reg     [31:0] VREG_15_7;
reg     [31:0] VREG_15_8;
reg     [31:0] VREG_15_9;
reg     [31:0] VREG_16_0;
reg     [31:0] VREG_16_1;
reg     [31:0] VREG_16_10;
reg     [31:0] VREG_16_11;
reg     [31:0] VREG_16_12;
reg     [31:0] VREG_16_13;
reg     [31:0] VREG_16_14;
reg     [31:0] VREG_16_15;
reg     [31:0] VREG_16_2;
reg     [31:0] VREG_16_3;
reg     [31:0] VREG_16_4;
reg     [31:0] VREG_16_5;
reg     [31:0] VREG_16_6;
reg     [31:0] VREG_16_7;
reg     [31:0] VREG_16_8;
reg     [31:0] VREG_16_9;
reg     [31:0] VREG_17_0;
reg     [31:0] VREG_17_1;
reg     [31:0] VREG_17_10;
reg     [31:0] VREG_17_11;
reg     [31:0] VREG_17_12;
reg     [31:0] VREG_17_13;
reg     [31:0] VREG_17_14;
reg     [31:0] VREG_17_15;
reg     [31:0] VREG_17_2;
reg     [31:0] VREG_17_3;
reg     [31:0] VREG_17_4;
reg     [31:0] VREG_17_5;
reg     [31:0] VREG_17_6;
reg     [31:0] VREG_17_7;
reg     [31:0] VREG_17_8;
reg     [31:0] VREG_17_9;
reg     [31:0] VREG_18_0;
reg     [31:0] VREG_18_1;
reg     [31:0] VREG_18_10;
reg     [31:0] VREG_18_11;
reg     [31:0] VREG_18_12;
reg     [31:0] VREG_18_13;
reg     [31:0] VREG_18_14;
reg     [31:0] VREG_18_15;
reg     [31:0] VREG_18_2;
reg     [31:0] VREG_18_3;
reg     [31:0] VREG_18_4;
reg     [31:0] VREG_18_5;
reg     [31:0] VREG_18_6;
reg     [31:0] VREG_18_7;
reg     [31:0] VREG_18_8;
reg     [31:0] VREG_18_9;
reg     [31:0] VREG_19_0;
reg     [31:0] VREG_19_1;
reg     [31:0] VREG_19_10;
reg     [31:0] VREG_19_11;
reg     [31:0] VREG_19_12;
reg     [31:0] VREG_19_13;
reg     [31:0] VREG_19_14;
reg     [31:0] VREG_19_15;
reg     [31:0] VREG_19_2;
reg     [31:0] VREG_19_3;
reg     [31:0] VREG_19_4;
reg     [31:0] VREG_19_5;
reg     [31:0] VREG_19_6;
reg     [31:0] VREG_19_7;
reg     [31:0] VREG_19_8;
reg     [31:0] VREG_19_9;
reg     [31:0] VREG_1_0;
reg     [31:0] VREG_1_1;
reg     [31:0] VREG_1_10;
reg     [31:0] VREG_1_11;
reg     [31:0] VREG_1_12;
reg     [31:0] VREG_1_13;
reg     [31:0] VREG_1_14;
reg     [31:0] VREG_1_15;
reg     [31:0] VREG_1_2;
reg     [31:0] VREG_1_3;
reg     [31:0] VREG_1_4;
reg     [31:0] VREG_1_5;
reg     [31:0] VREG_1_6;
reg     [31:0] VREG_1_7;
reg     [31:0] VREG_1_8;
reg     [31:0] VREG_1_9;
reg     [31:0] VREG_20_0;
reg     [31:0] VREG_20_1;
reg     [31:0] VREG_20_10;
reg     [31:0] VREG_20_11;
reg     [31:0] VREG_20_12;
reg     [31:0] VREG_20_13;
reg     [31:0] VREG_20_14;
reg     [31:0] VREG_20_15;
reg     [31:0] VREG_20_2;
reg     [31:0] VREG_20_3;
reg     [31:0] VREG_20_4;
reg     [31:0] VREG_20_5;
reg     [31:0] VREG_20_6;
reg     [31:0] VREG_20_7;
reg     [31:0] VREG_20_8;
reg     [31:0] VREG_20_9;
reg     [31:0] VREG_21_0;
reg     [31:0] VREG_21_1;
reg     [31:0] VREG_21_10;
reg     [31:0] VREG_21_11;
reg     [31:0] VREG_21_12;
reg     [31:0] VREG_21_13;
reg     [31:0] VREG_21_14;
reg     [31:0] VREG_21_15;
reg     [31:0] VREG_21_2;
reg     [31:0] VREG_21_3;
reg     [31:0] VREG_21_4;
reg     [31:0] VREG_21_5;
reg     [31:0] VREG_21_6;
reg     [31:0] VREG_21_7;
reg     [31:0] VREG_21_8;
reg     [31:0] VREG_21_9;
reg     [31:0] VREG_22_0;
reg     [31:0] VREG_22_1;
reg     [31:0] VREG_22_10;
reg     [31:0] VREG_22_11;
reg     [31:0] VREG_22_12;
reg     [31:0] VREG_22_13;
reg     [31:0] VREG_22_14;
reg     [31:0] VREG_22_15;
reg     [31:0] VREG_22_2;
reg     [31:0] VREG_22_3;
reg     [31:0] VREG_22_4;
reg     [31:0] VREG_22_5;
reg     [31:0] VREG_22_6;
reg     [31:0] VREG_22_7;
reg     [31:0] VREG_22_8;
reg     [31:0] VREG_22_9;
reg     [31:0] VREG_23_0;
reg     [31:0] VREG_23_1;
reg     [31:0] VREG_23_10;
reg     [31:0] VREG_23_11;
reg     [31:0] VREG_23_12;
reg     [31:0] VREG_23_13;
reg     [31:0] VREG_23_14;
reg     [31:0] VREG_23_15;
reg     [31:0] VREG_23_2;
reg     [31:0] VREG_23_3;
reg     [31:0] VREG_23_4;
reg     [31:0] VREG_23_5;
reg     [31:0] VREG_23_6;
reg     [31:0] VREG_23_7;
reg     [31:0] VREG_23_8;
reg     [31:0] VREG_23_9;
reg     [31:0] VREG_24_0;
reg     [31:0] VREG_24_1;
reg     [31:0] VREG_24_10;
reg     [31:0] VREG_24_11;
reg     [31:0] VREG_24_12;
reg     [31:0] VREG_24_13;
reg     [31:0] VREG_24_14;
reg     [31:0] VREG_24_15;
reg     [31:0] VREG_24_2;
reg     [31:0] VREG_24_3;
reg     [31:0] VREG_24_4;
reg     [31:0] VREG_24_5;
reg     [31:0] VREG_24_6;
reg     [31:0] VREG_24_7;
reg     [31:0] VREG_24_8;
reg     [31:0] VREG_24_9;
reg     [31:0] VREG_25_0;
reg     [31:0] VREG_25_1;
reg     [31:0] VREG_25_10;
reg     [31:0] VREG_25_11;
reg     [31:0] VREG_25_12;
reg     [31:0] VREG_25_13;
reg     [31:0] VREG_25_14;
reg     [31:0] VREG_25_15;
reg     [31:0] VREG_25_2;
reg     [31:0] VREG_25_3;
reg     [31:0] VREG_25_4;
reg     [31:0] VREG_25_5;
reg     [31:0] VREG_25_6;
reg     [31:0] VREG_25_7;
reg     [31:0] VREG_25_8;
reg     [31:0] VREG_25_9;
reg     [31:0] VREG_26_0;
reg     [31:0] VREG_26_1;
reg     [31:0] VREG_26_10;
reg     [31:0] VREG_26_11;
reg     [31:0] VREG_26_12;
reg     [31:0] VREG_26_13;
reg     [31:0] VREG_26_14;
reg     [31:0] VREG_26_15;
reg     [31:0] VREG_26_2;
reg     [31:0] VREG_26_3;
reg     [31:0] VREG_26_4;
reg     [31:0] VREG_26_5;
reg     [31:0] VREG_26_6;
reg     [31:0] VREG_26_7;
reg     [31:0] VREG_26_8;
reg     [31:0] VREG_26_9;
reg     [31:0] VREG_27_0;
reg     [31:0] VREG_27_1;
reg     [31:0] VREG_27_10;
reg     [31:0] VREG_27_11;
reg     [31:0] VREG_27_12;
reg     [31:0] VREG_27_13;
reg     [31:0] VREG_27_14;
reg     [31:0] VREG_27_15;
reg     [31:0] VREG_27_2;
reg     [31:0] VREG_27_3;
reg     [31:0] VREG_27_4;
reg     [31:0] VREG_27_5;
reg     [31:0] VREG_27_6;
reg     [31:0] VREG_27_7;
reg     [31:0] VREG_27_8;
reg     [31:0] VREG_27_9;
reg     [31:0] VREG_28_0;
reg     [31:0] VREG_28_1;
reg     [31:0] VREG_28_10;
reg     [31:0] VREG_28_11;
reg     [31:0] VREG_28_12;
reg     [31:0] VREG_28_13;
reg     [31:0] VREG_28_14;
reg     [31:0] VREG_28_15;
reg     [31:0] VREG_28_2;
reg     [31:0] VREG_28_3;
reg     [31:0] VREG_28_4;
reg     [31:0] VREG_28_5;
reg     [31:0] VREG_28_6;
reg     [31:0] VREG_28_7;
reg     [31:0] VREG_28_8;
reg     [31:0] VREG_28_9;
reg     [31:0] VREG_29_0;
reg     [31:0] VREG_29_1;
reg     [31:0] VREG_29_10;
reg     [31:0] VREG_29_11;
reg     [31:0] VREG_29_12;
reg     [31:0] VREG_29_13;
reg     [31:0] VREG_29_14;
reg     [31:0] VREG_29_15;
reg     [31:0] VREG_29_2;
reg     [31:0] VREG_29_3;
reg     [31:0] VREG_29_4;
reg     [31:0] VREG_29_5;
reg     [31:0] VREG_29_6;
reg     [31:0] VREG_29_7;
reg     [31:0] VREG_29_8;
reg     [31:0] VREG_29_9;
reg     [31:0] VREG_2_0;
reg     [31:0] VREG_2_1;
reg     [31:0] VREG_2_10;
reg     [31:0] VREG_2_11;
reg     [31:0] VREG_2_12;
reg     [31:0] VREG_2_13;
reg     [31:0] VREG_2_14;
reg     [31:0] VREG_2_15;
reg     [31:0] VREG_2_2;
reg     [31:0] VREG_2_3;
reg     [31:0] VREG_2_4;
reg     [31:0] VREG_2_5;
reg     [31:0] VREG_2_6;
reg     [31:0] VREG_2_7;
reg     [31:0] VREG_2_8;
reg     [31:0] VREG_2_9;
reg     [31:0] VREG_30_0;
reg     [31:0] VREG_30_1;
reg     [31:0] VREG_30_10;
reg     [31:0] VREG_30_11;
reg     [31:0] VREG_30_12;
reg     [31:0] VREG_30_13;
reg     [31:0] VREG_30_14;
reg     [31:0] VREG_30_15;
reg     [31:0] VREG_30_2;
reg     [31:0] VREG_30_3;
reg     [31:0] VREG_30_4;
reg     [31:0] VREG_30_5;
reg     [31:0] VREG_30_6;
reg     [31:0] VREG_30_7;
reg     [31:0] VREG_30_8;
reg     [31:0] VREG_30_9;
reg     [31:0] VREG_31_0;
reg     [31:0] VREG_31_1;
reg     [31:0] VREG_31_10;
reg     [31:0] VREG_31_11;
reg     [31:0] VREG_31_12;
reg     [31:0] VREG_31_13;
reg     [31:0] VREG_31_14;
reg     [31:0] VREG_31_15;
reg     [31:0] VREG_31_2;
reg     [31:0] VREG_31_3;
reg     [31:0] VREG_31_4;
reg     [31:0] VREG_31_5;
reg     [31:0] VREG_31_6;
reg     [31:0] VREG_31_7;
reg     [31:0] VREG_31_8;
reg     [31:0] VREG_31_9;
reg     [31:0] VREG_3_0;
reg     [31:0] VREG_3_1;
reg     [31:0] VREG_3_10;
reg     [31:0] VREG_3_11;
reg     [31:0] VREG_3_12;
reg     [31:0] VREG_3_13;
reg     [31:0] VREG_3_14;
reg     [31:0] VREG_3_15;
reg     [31:0] VREG_3_2;
reg     [31:0] VREG_3_3;
reg     [31:0] VREG_3_4;
reg     [31:0] VREG_3_5;
reg     [31:0] VREG_3_6;
reg     [31:0] VREG_3_7;
reg     [31:0] VREG_3_8;
reg     [31:0] VREG_3_9;
reg     [31:0] VREG_4_0;
reg     [31:0] VREG_4_1;
reg     [31:0] VREG_4_10;
reg     [31:0] VREG_4_11;
reg     [31:0] VREG_4_12;
reg     [31:0] VREG_4_13;
reg     [31:0] VREG_4_14;
reg     [31:0] VREG_4_15;
reg     [31:0] VREG_4_2;
reg     [31:0] VREG_4_3;
reg     [31:0] VREG_4_4;
reg     [31:0] VREG_4_5;
reg     [31:0] VREG_4_6;
reg     [31:0] VREG_4_7;
reg     [31:0] VREG_4_8;
reg     [31:0] VREG_4_9;
reg     [31:0] VREG_5_0;
reg     [31:0] VREG_5_1;
reg     [31:0] VREG_5_10;
reg     [31:0] VREG_5_11;
reg     [31:0] VREG_5_12;
reg     [31:0] VREG_5_13;
reg     [31:0] VREG_5_14;
reg     [31:0] VREG_5_15;
reg     [31:0] VREG_5_2;
reg     [31:0] VREG_5_3;
reg     [31:0] VREG_5_4;
reg     [31:0] VREG_5_5;
reg     [31:0] VREG_5_6;
reg     [31:0] VREG_5_7;
reg     [31:0] VREG_5_8;
reg     [31:0] VREG_5_9;
reg     [31:0] VREG_6_0;
reg     [31:0] VREG_6_1;
reg     [31:0] VREG_6_10;
reg     [31:0] VREG_6_11;
reg     [31:0] VREG_6_12;
reg     [31:0] VREG_6_13;
reg     [31:0] VREG_6_14;
reg     [31:0] VREG_6_15;
reg     [31:0] VREG_6_2;
reg     [31:0] VREG_6_3;
reg     [31:0] VREG_6_4;
reg     [31:0] VREG_6_5;
reg     [31:0] VREG_6_6;
reg     [31:0] VREG_6_7;
reg     [31:0] VREG_6_8;
reg     [31:0] VREG_6_9;
reg     [31:0] VREG_7_0;
reg     [31:0] VREG_7_1;
reg     [31:0] VREG_7_10;
reg     [31:0] VREG_7_11;
reg     [31:0] VREG_7_12;
reg     [31:0] VREG_7_13;
reg     [31:0] VREG_7_14;
reg     [31:0] VREG_7_15;
reg     [31:0] VREG_7_2;
reg     [31:0] VREG_7_3;
reg     [31:0] VREG_7_4;
reg     [31:0] VREG_7_5;
reg     [31:0] VREG_7_6;
reg     [31:0] VREG_7_7;
reg     [31:0] VREG_7_8;
reg     [31:0] VREG_7_9;
reg     [31:0] VREG_8_0;
reg     [31:0] VREG_8_1;
reg     [31:0] VREG_8_10;
reg     [31:0] VREG_8_11;
reg     [31:0] VREG_8_12;
reg     [31:0] VREG_8_13;
reg     [31:0] VREG_8_14;
reg     [31:0] VREG_8_15;
reg     [31:0] VREG_8_2;
reg     [31:0] VREG_8_3;
reg     [31:0] VREG_8_4;
reg     [31:0] VREG_8_5;
reg     [31:0] VREG_8_6;
reg     [31:0] VREG_8_7;
reg     [31:0] VREG_8_8;
reg     [31:0] VREG_8_9;
reg     [31:0] VREG_9_0;
reg     [31:0] VREG_9_1;
reg     [31:0] VREG_9_10;
reg     [31:0] VREG_9_11;
reg     [31:0] VREG_9_12;
reg     [31:0] VREG_9_13;
reg     [31:0] VREG_9_14;
reg     [31:0] VREG_9_15;
reg     [31:0] VREG_9_2;
reg     [31:0] VREG_9_3;
reg     [31:0] VREG_9_4;
reg     [31:0] VREG_9_5;
reg     [31:0] VREG_9_6;
reg     [31:0] VREG_9_7;
reg     [31:0] VREG_9_8;
reg     [31:0] VREG_9_9;
reg     [31:0] pc;
reg     [31:0] vector_mask_register;
wire     [29:0] n0;
wire     [31:0] n1;
wire     [31:0] n2;
wire      [4:0] n3;
wire            n4;
wire      [2:0] n5;
wire            n6;
wire      [2:0] n7;
wire            n8;
wire      [5:0] n9;
wire            n10;
wire      [4:0] n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire     [31:0] n44;
wire     [31:0] n45;
wire     [31:0] n46;
wire     [31:0] n47;
wire     [31:0] n48;
wire     [31:0] n49;
wire     [31:0] n50;
wire     [31:0] n51;
wire     [31:0] n52;
wire     [31:0] n53;
wire     [31:0] n54;
wire     [31:0] n55;
wire     [31:0] n56;
wire     [31:0] n57;
wire     [31:0] n58;
wire     [31:0] n59;
wire     [31:0] n60;
wire     [31:0] n61;
wire     [31:0] n62;
wire     [31:0] n63;
wire     [31:0] n64;
wire     [31:0] n65;
wire     [31:0] n66;
wire     [31:0] n67;
wire     [31:0] n68;
wire     [31:0] n69;
wire     [31:0] n70;
wire     [31:0] n71;
wire     [31:0] n72;
wire     [31:0] n73;
wire     [31:0] n74;
wire     [31:0] n75;
wire      [4:0] n76;
wire            n77;
wire            n78;
wire            n79;
wire            n80;
wire            n81;
wire            n82;
wire            n83;
wire            n84;
wire            n85;
wire            n86;
wire            n87;
wire            n88;
wire            n89;
wire            n90;
wire            n91;
wire            n92;
wire            n93;
wire            n94;
wire            n95;
wire            n96;
wire            n97;
wire            n98;
wire            n99;
wire            n100;
wire            n101;
wire            n102;
wire            n103;
wire            n104;
wire            n105;
wire            n106;
wire            n107;
wire            n108;
wire     [31:0] n109;
wire     [31:0] n110;
wire     [31:0] n111;
wire     [31:0] n112;
wire     [31:0] n113;
wire     [31:0] n114;
wire     [31:0] n115;
wire     [31:0] n116;
wire     [31:0] n117;
wire     [31:0] n118;
wire     [31:0] n119;
wire     [31:0] n120;
wire     [31:0] n121;
wire     [31:0] n122;
wire     [31:0] n123;
wire     [31:0] n124;
wire     [31:0] n125;
wire     [31:0] n126;
wire     [31:0] n127;
wire     [31:0] n128;
wire     [31:0] n129;
wire     [31:0] n130;
wire     [31:0] n131;
wire     [31:0] n132;
wire     [31:0] n133;
wire     [31:0] n134;
wire     [31:0] n135;
wire     [31:0] n136;
wire     [31:0] n137;
wire     [31:0] n138;
wire     [31:0] n139;
wire     [31:0] n140;
wire     [31:0] n141;
wire            n142;
wire     [31:0] n143;
wire            n144;
wire     [31:0] n145;
wire            n146;
wire     [31:0] n147;
wire            n148;
wire     [31:0] n149;
wire     [31:0] n150;
wire     [31:0] n151;
wire     [31:0] n152;
wire     [31:0] n153;
wire     [31:0] n154;
wire     [31:0] n155;
wire            n156;
wire            n157;
wire      [1:0] n158;
wire            n159;
wire      [4:0] n160;
wire      [5:0] n161;
wire            n162;
wire     [13:0] n163;
wire     [31:0] n164;
wire     [31:0] n165;
wire            n166;
wire     [31:0] n167;
wire            n168;
wire     [31:0] n169;
wire            n170;
wire     [31:0] n171;
wire            n172;
wire     [31:0] n173;
wire     [31:0] n174;
wire     [31:0] n175;
wire     [31:0] n176;
wire     [31:0] n177;
wire            n178;
wire      [8:0] n179;
wire     [31:0] n180;
wire     [31:0] n181;
wire     [31:0] n182;
wire     [31:0] n183;
wire     [31:0] n184;
wire     [31:0] n185;
wire     [31:0] n186;
wire     [31:0] n187;
wire     [31:0] n188;
wire     [31:0] n189;
wire     [31:0] n190;
wire            n191;
wire            n192;
wire     [31:0] n193;
wire     [31:0] n194;
wire     [31:0] n195;
wire     [31:0] n196;
wire            n197;
wire     [31:0] n198;
wire     [31:0] n199;
wire     [31:0] n200;
wire     [31:0] n201;
wire     [31:0] n202;
wire     [31:0] n203;
wire     [31:0] n204;
wire     [31:0] n205;
wire     [31:0] n206;
wire     [31:0] n207;
wire     [31:0] n208;
wire     [31:0] n209;
wire     [31:0] n210;
wire     [31:0] n211;
wire     [31:0] n212;
wire     [31:0] n213;
wire     [31:0] n214;
wire     [31:0] n215;
wire     [31:0] n216;
wire     [31:0] n217;
wire     [31:0] n218;
wire            n219;
wire     [31:0] n220;
wire     [31:0] n221;
wire     [31:0] n222;
wire     [31:0] n223;
wire     [31:0] n224;
wire     [31:0] n225;
wire     [31:0] n226;
wire     [31:0] n227;
wire     [31:0] n228;
wire     [31:0] n229;
wire     [31:0] n230;
wire     [31:0] n231;
wire     [31:0] n232;
wire     [31:0] n233;
wire     [31:0] n234;
wire     [31:0] n235;
wire     [31:0] n236;
wire     [31:0] n237;
wire     [31:0] n238;
wire     [31:0] n239;
wire     [31:0] n240;
wire            n241;
wire     [31:0] n242;
wire     [31:0] n243;
wire     [31:0] n244;
wire     [31:0] n245;
wire     [31:0] n246;
wire     [31:0] n247;
wire     [31:0] n248;
wire     [31:0] n249;
wire     [31:0] n250;
wire     [31:0] n251;
wire     [31:0] n252;
wire     [31:0] n253;
wire     [31:0] n254;
wire     [31:0] n255;
wire     [31:0] n256;
wire     [31:0] n257;
wire     [31:0] n258;
wire     [31:0] n259;
wire     [31:0] n260;
wire     [31:0] n261;
wire     [31:0] n262;
wire            n263;
wire     [31:0] n264;
wire     [31:0] n265;
wire     [31:0] n266;
wire     [31:0] n267;
wire     [31:0] n268;
wire     [31:0] n269;
wire     [31:0] n270;
wire     [31:0] n271;
wire     [31:0] n272;
wire     [31:0] n273;
wire     [31:0] n274;
wire     [31:0] n275;
wire     [31:0] n276;
wire     [31:0] n277;
wire     [31:0] n278;
wire     [31:0] n279;
wire     [31:0] n280;
wire     [31:0] n281;
wire     [31:0] n282;
wire     [31:0] n283;
wire     [31:0] n284;
wire            n285;
wire     [31:0] n286;
wire     [31:0] n287;
wire     [31:0] n288;
wire     [31:0] n289;
wire     [31:0] n290;
wire     [31:0] n291;
wire     [31:0] n292;
wire     [31:0] n293;
wire     [31:0] n294;
wire     [31:0] n295;
wire     [31:0] n296;
wire     [31:0] n297;
wire     [31:0] n298;
wire     [31:0] n299;
wire     [31:0] n300;
wire     [31:0] n301;
wire     [31:0] n302;
wire     [31:0] n303;
wire     [31:0] n304;
wire     [31:0] n305;
wire     [31:0] n306;
wire            n307;
wire     [31:0] n308;
wire     [31:0] n309;
wire     [31:0] n310;
wire     [31:0] n311;
wire     [31:0] n312;
wire     [31:0] n313;
wire     [31:0] n314;
wire     [31:0] n315;
wire     [31:0] n316;
wire     [31:0] n317;
wire     [31:0] n318;
wire     [31:0] n319;
wire     [31:0] n320;
wire     [31:0] n321;
wire     [31:0] n322;
wire     [31:0] n323;
wire     [31:0] n324;
wire     [31:0] n325;
wire     [31:0] n326;
wire     [31:0] n327;
wire     [31:0] n328;
wire            n329;
wire     [31:0] n330;
wire     [31:0] n331;
wire     [31:0] n332;
wire     [31:0] n333;
wire     [31:0] n334;
wire     [31:0] n335;
wire     [31:0] n336;
wire     [31:0] n337;
wire     [31:0] n338;
wire     [31:0] n339;
wire     [31:0] n340;
wire     [31:0] n341;
wire     [31:0] n342;
wire     [31:0] n343;
wire     [31:0] n344;
wire     [31:0] n345;
wire     [31:0] n346;
wire     [31:0] n347;
wire     [31:0] n348;
wire     [31:0] n349;
wire     [31:0] n350;
wire            n351;
wire     [31:0] n352;
wire     [31:0] n353;
wire     [31:0] n354;
wire     [31:0] n355;
wire     [31:0] n356;
wire     [31:0] n357;
wire     [31:0] n358;
wire     [31:0] n359;
wire     [31:0] n360;
wire     [31:0] n361;
wire     [31:0] n362;
wire     [31:0] n363;
wire     [31:0] n364;
wire     [31:0] n365;
wire     [31:0] n366;
wire     [31:0] n367;
wire     [31:0] n368;
wire     [31:0] n369;
wire     [31:0] n370;
wire     [31:0] n371;
wire     [31:0] n372;
wire            n373;
wire     [31:0] n374;
wire     [31:0] n375;
wire     [31:0] n376;
wire     [31:0] n377;
wire     [31:0] n378;
wire     [31:0] n379;
wire     [31:0] n380;
wire     [31:0] n381;
wire     [31:0] n382;
wire     [31:0] n383;
wire     [31:0] n384;
wire     [31:0] n385;
wire     [31:0] n386;
wire     [31:0] n387;
wire     [31:0] n388;
wire     [31:0] n389;
wire     [31:0] n390;
wire     [31:0] n391;
wire     [31:0] n392;
wire     [31:0] n393;
wire     [31:0] n394;
wire            n395;
wire     [31:0] n396;
wire     [31:0] n397;
wire     [31:0] n398;
wire     [31:0] n399;
wire     [31:0] n400;
wire     [31:0] n401;
wire     [31:0] n402;
wire     [31:0] n403;
wire     [31:0] n404;
wire     [31:0] n405;
wire     [31:0] n406;
wire     [31:0] n407;
wire     [31:0] n408;
wire     [31:0] n409;
wire     [31:0] n410;
wire     [31:0] n411;
wire     [31:0] n412;
wire     [31:0] n413;
wire     [31:0] n414;
wire     [31:0] n415;
wire     [31:0] n416;
wire            n417;
wire     [31:0] n418;
wire     [31:0] n419;
wire     [31:0] n420;
wire     [31:0] n421;
wire     [31:0] n422;
wire     [31:0] n423;
wire     [31:0] n424;
wire     [31:0] n425;
wire     [31:0] n426;
wire     [31:0] n427;
wire     [31:0] n428;
wire     [31:0] n429;
wire     [31:0] n430;
wire     [31:0] n431;
wire     [31:0] n432;
wire     [31:0] n433;
wire     [31:0] n434;
wire     [31:0] n435;
wire     [31:0] n436;
wire     [31:0] n437;
wire     [31:0] n438;
wire            n439;
wire     [31:0] n440;
wire     [31:0] n441;
wire     [31:0] n442;
wire     [31:0] n443;
wire     [31:0] n444;
wire     [31:0] n445;
wire     [31:0] n446;
wire     [31:0] n447;
wire     [31:0] n448;
wire     [31:0] n449;
wire     [31:0] n450;
wire     [31:0] n451;
wire     [31:0] n452;
wire     [31:0] n453;
wire     [31:0] n454;
wire     [31:0] n455;
wire     [31:0] n456;
wire     [31:0] n457;
wire     [31:0] n458;
wire     [31:0] n459;
wire     [31:0] n460;
wire            n461;
wire     [31:0] n462;
wire     [31:0] n463;
wire     [31:0] n464;
wire     [31:0] n465;
wire     [31:0] n466;
wire     [31:0] n467;
wire     [31:0] n468;
wire     [31:0] n469;
wire     [31:0] n470;
wire     [31:0] n471;
wire     [31:0] n472;
wire     [31:0] n473;
wire     [31:0] n474;
wire     [31:0] n475;
wire     [31:0] n476;
wire     [31:0] n477;
wire     [31:0] n478;
wire     [31:0] n479;
wire     [31:0] n480;
wire     [31:0] n481;
wire     [31:0] n482;
wire            n483;
wire     [31:0] n484;
wire     [31:0] n485;
wire     [31:0] n486;
wire     [31:0] n487;
wire     [31:0] n488;
wire     [31:0] n489;
wire     [31:0] n490;
wire     [31:0] n491;
wire     [31:0] n492;
wire     [31:0] n493;
wire     [31:0] n494;
wire     [31:0] n495;
wire     [31:0] n496;
wire     [31:0] n497;
wire     [31:0] n498;
wire     [31:0] n499;
wire     [31:0] n500;
wire     [31:0] n501;
wire     [31:0] n502;
wire     [31:0] n503;
wire     [31:0] n504;
wire            n505;
wire     [31:0] n506;
wire     [31:0] n507;
wire     [31:0] n508;
wire     [31:0] n509;
wire     [31:0] n510;
wire     [31:0] n511;
wire     [31:0] n512;
wire     [31:0] n513;
wire     [31:0] n514;
wire     [31:0] n515;
wire     [31:0] n516;
wire     [31:0] n517;
wire     [31:0] n518;
wire     [31:0] n519;
wire     [31:0] n520;
wire     [31:0] n521;
wire     [31:0] n522;
wire     [31:0] n523;
wire     [31:0] n524;
wire     [31:0] n525;
wire     [31:0] n526;
wire            n527;
wire     [31:0] n528;
wire     [31:0] n529;
wire     [31:0] n530;
wire     [31:0] n531;
wire     [31:0] n532;
wire     [31:0] n533;
wire     [31:0] n534;
wire     [31:0] n535;
wire     [31:0] n536;
wire     [31:0] n537;
wire     [31:0] n538;
wire     [31:0] n539;
wire     [31:0] n540;
wire     [31:0] n541;
wire     [31:0] n542;
wire     [31:0] n543;
wire     [31:0] n544;
wire     [31:0] n545;
wire     [31:0] n546;
wire     [31:0] n547;
wire     [31:0] n548;
wire            n549;
wire     [31:0] n550;
wire     [31:0] n551;
wire     [31:0] n552;
wire     [31:0] n553;
wire     [31:0] n554;
wire     [31:0] n555;
wire     [31:0] n556;
wire     [31:0] n557;
wire     [31:0] n558;
wire     [31:0] n559;
wire     [31:0] n560;
wire     [31:0] n561;
wire     [31:0] n562;
wire     [31:0] n563;
wire     [31:0] n564;
wire     [31:0] n565;
wire     [31:0] n566;
wire     [31:0] n567;
wire     [31:0] n568;
wire     [31:0] n569;
wire     [31:0] n570;
wire            n571;
wire     [31:0] n572;
wire     [31:0] n573;
wire     [31:0] n574;
wire     [31:0] n575;
wire     [31:0] n576;
wire     [31:0] n577;
wire     [31:0] n578;
wire     [31:0] n579;
wire     [31:0] n580;
wire     [31:0] n581;
wire     [31:0] n582;
wire     [31:0] n583;
wire     [31:0] n584;
wire     [31:0] n585;
wire     [31:0] n586;
wire     [31:0] n587;
wire     [31:0] n588;
wire     [31:0] n589;
wire     [31:0] n590;
wire     [31:0] n591;
wire     [31:0] n592;
wire            n593;
wire     [31:0] n594;
wire     [31:0] n595;
wire     [31:0] n596;
wire     [31:0] n597;
wire     [31:0] n598;
wire     [31:0] n599;
wire     [31:0] n600;
wire     [31:0] n601;
wire     [31:0] n602;
wire     [31:0] n603;
wire     [31:0] n604;
wire     [31:0] n605;
wire     [31:0] n606;
wire     [31:0] n607;
wire     [31:0] n608;
wire     [31:0] n609;
wire     [31:0] n610;
wire     [31:0] n611;
wire     [31:0] n612;
wire     [31:0] n613;
wire     [31:0] n614;
wire            n615;
wire     [31:0] n616;
wire     [31:0] n617;
wire     [31:0] n618;
wire     [31:0] n619;
wire     [31:0] n620;
wire     [31:0] n621;
wire     [31:0] n622;
wire     [31:0] n623;
wire     [31:0] n624;
wire     [31:0] n625;
wire     [31:0] n626;
wire     [31:0] n627;
wire     [31:0] n628;
wire     [31:0] n629;
wire     [31:0] n630;
wire     [31:0] n631;
wire     [31:0] n632;
wire     [31:0] n633;
wire     [31:0] n634;
wire     [31:0] n635;
wire     [31:0] n636;
wire            n637;
wire     [31:0] n638;
wire     [31:0] n639;
wire     [31:0] n640;
wire     [31:0] n641;
wire     [31:0] n642;
wire     [31:0] n643;
wire     [31:0] n644;
wire     [31:0] n645;
wire     [31:0] n646;
wire     [31:0] n647;
wire     [31:0] n648;
wire     [31:0] n649;
wire     [31:0] n650;
wire     [31:0] n651;
wire     [31:0] n652;
wire     [31:0] n653;
wire     [31:0] n654;
wire     [31:0] n655;
wire     [31:0] n656;
wire     [31:0] n657;
wire     [31:0] n658;
wire            n659;
wire     [31:0] n660;
wire     [31:0] n661;
wire     [31:0] n662;
wire     [31:0] n663;
wire     [31:0] n664;
wire     [31:0] n665;
wire     [31:0] n666;
wire     [31:0] n667;
wire     [31:0] n668;
wire     [31:0] n669;
wire     [31:0] n670;
wire     [31:0] n671;
wire     [31:0] n672;
wire     [31:0] n673;
wire     [31:0] n674;
wire     [31:0] n675;
wire     [31:0] n676;
wire     [31:0] n677;
wire     [31:0] n678;
wire     [31:0] n679;
wire     [31:0] n680;
wire            n681;
wire     [31:0] n682;
wire     [31:0] n683;
wire     [31:0] n684;
wire     [31:0] n685;
wire     [31:0] n686;
wire     [31:0] n687;
wire     [31:0] n688;
wire     [31:0] n689;
wire     [31:0] n690;
wire     [31:0] n691;
wire     [31:0] n692;
wire     [31:0] n693;
wire     [31:0] n694;
wire     [31:0] n695;
wire     [31:0] n696;
wire     [31:0] n697;
wire     [31:0] n698;
wire     [31:0] n699;
wire     [31:0] n700;
wire     [31:0] n701;
wire     [31:0] n702;
wire            n703;
wire     [31:0] n704;
wire     [31:0] n705;
wire     [31:0] n706;
wire     [31:0] n707;
wire     [31:0] n708;
wire     [31:0] n709;
wire     [31:0] n710;
wire     [31:0] n711;
wire     [31:0] n712;
wire     [31:0] n713;
wire     [31:0] n714;
wire     [31:0] n715;
wire     [31:0] n716;
wire     [31:0] n717;
wire     [31:0] n718;
wire     [31:0] n719;
wire     [31:0] n720;
wire     [31:0] n721;
wire     [31:0] n722;
wire     [31:0] n723;
wire     [31:0] n724;
wire            n725;
wire     [31:0] n726;
wire     [31:0] n727;
wire     [31:0] n728;
wire     [31:0] n729;
wire     [31:0] n730;
wire     [31:0] n731;
wire     [31:0] n732;
wire     [31:0] n733;
wire     [31:0] n734;
wire     [31:0] n735;
wire     [31:0] n736;
wire     [31:0] n737;
wire     [31:0] n738;
wire     [31:0] n739;
wire     [31:0] n740;
wire     [31:0] n741;
wire     [31:0] n742;
wire     [31:0] n743;
wire     [31:0] n744;
wire     [31:0] n745;
wire     [31:0] n746;
wire            n747;
wire     [31:0] n748;
wire     [31:0] n749;
wire     [31:0] n750;
wire     [31:0] n751;
wire     [31:0] n752;
wire     [31:0] n753;
wire     [31:0] n754;
wire     [31:0] n755;
wire     [31:0] n756;
wire     [31:0] n757;
wire     [31:0] n758;
wire     [31:0] n759;
wire     [31:0] n760;
wire     [31:0] n761;
wire     [31:0] n762;
wire     [31:0] n763;
wire     [31:0] n764;
wire     [31:0] n765;
wire     [31:0] n766;
wire     [31:0] n767;
wire     [31:0] n768;
wire            n769;
wire     [31:0] n770;
wire     [31:0] n771;
wire     [31:0] n772;
wire     [31:0] n773;
wire     [31:0] n774;
wire     [31:0] n775;
wire     [31:0] n776;
wire     [31:0] n777;
wire     [31:0] n778;
wire     [31:0] n779;
wire     [31:0] n780;
wire     [31:0] n781;
wire     [31:0] n782;
wire     [31:0] n783;
wire     [31:0] n784;
wire     [31:0] n785;
wire     [31:0] n786;
wire     [31:0] n787;
wire     [31:0] n788;
wire     [31:0] n789;
wire     [31:0] n790;
wire            n791;
wire     [31:0] n792;
wire     [31:0] n793;
wire     [31:0] n794;
wire     [31:0] n795;
wire     [31:0] n796;
wire     [31:0] n797;
wire     [31:0] n798;
wire     [31:0] n799;
wire     [31:0] n800;
wire     [31:0] n801;
wire     [31:0] n802;
wire     [31:0] n803;
wire     [31:0] n804;
wire     [31:0] n805;
wire     [31:0] n806;
wire     [31:0] n807;
wire     [31:0] n808;
wire     [31:0] n809;
wire     [31:0] n810;
wire     [31:0] n811;
wire     [31:0] n812;
wire            n813;
wire     [31:0] n814;
wire     [31:0] n815;
wire     [31:0] n816;
wire     [31:0] n817;
wire     [31:0] n818;
wire     [31:0] n819;
wire     [31:0] n820;
wire     [31:0] n821;
wire     [31:0] n822;
wire     [31:0] n823;
wire     [31:0] n824;
wire     [31:0] n825;
wire     [31:0] n826;
wire     [31:0] n827;
wire     [31:0] n828;
wire     [31:0] n829;
wire     [31:0] n830;
wire     [31:0] n831;
wire     [31:0] n832;
wire     [31:0] n833;
wire     [31:0] n834;
wire            n835;
wire     [31:0] n836;
wire     [31:0] n837;
wire     [31:0] n838;
wire     [31:0] n839;
wire     [31:0] n840;
wire     [31:0] n841;
wire     [31:0] n842;
wire     [31:0] n843;
wire     [31:0] n844;
wire     [31:0] n845;
wire     [31:0] n846;
wire     [31:0] n847;
wire     [31:0] n848;
wire     [31:0] n849;
wire     [31:0] n850;
wire     [31:0] n851;
wire     [31:0] n852;
wire     [31:0] n853;
wire     [31:0] n854;
wire     [31:0] n855;
wire     [31:0] n856;
wire            n857;
wire     [31:0] n858;
wire     [31:0] n859;
wire     [31:0] n860;
wire     [31:0] n861;
wire     [31:0] n862;
wire     [31:0] n863;
wire     [31:0] n864;
wire     [31:0] n865;
wire     [31:0] n866;
wire     [31:0] n867;
wire     [31:0] n868;
wire     [31:0] n869;
wire     [31:0] n870;
wire     [31:0] n871;
wire     [31:0] n872;
wire     [31:0] n873;
wire     [31:0] n874;
wire     [31:0] n875;
wire     [31:0] n876;
wire     [31:0] n877;
wire     [31:0] n878;
wire            n879;
wire            n880;
wire            n881;
wire            n882;
wire            n883;
wire            n884;
wire            n885;
wire            n886;
wire            n887;
wire            n888;
wire            n889;
wire            n890;
wire            n891;
wire            n892;
wire            n893;
wire            n894;
wire            n895;
wire            n896;
wire            n897;
wire            n898;
wire            n899;
wire            n900;
wire            n901;
wire            n902;
wire            n903;
wire            n904;
wire            n905;
wire            n906;
wire            n907;
wire            n908;
wire            n909;
wire            n910;
wire            n911;
wire            n912;
wire            n913;
wire            n914;
wire            n915;
wire            n916;
wire            n917;
wire            n918;
wire            n919;
wire            n920;
wire            n921;
wire            n922;
wire            n923;
wire            n924;
wire            n925;
wire            n926;
wire            n927;
wire            n928;
wire            n929;
wire            n930;
wire            n931;
wire            n932;
wire            n933;
wire            n934;
wire            n935;
wire            n936;
wire            n937;
wire            n938;
wire            n939;
wire            n940;
wire            n941;
wire            n942;
wire            n943;
wire            n944;
wire            n945;
wire            n946;
wire            n947;
wire            n948;
wire            n949;
wire            n950;
wire            n951;
wire            n952;
wire            n953;
wire            n954;
wire            n955;
wire            n956;
wire            n957;
wire            n958;
wire            n959;
wire            n960;
wire            n961;
wire            n962;
wire            n963;
wire            n964;
wire            n965;
wire            n966;
wire            n967;
wire            n968;
wire            n969;
wire            n970;
wire            n971;
wire            n972;
wire            n973;
wire            n974;
wire            n975;
wire            n976;
wire            n977;
wire            n978;
wire            n979;
wire            n980;
wire            n981;
wire            n982;
wire            n983;
wire            n984;
wire            n985;
wire            n986;
wire            n987;
wire            n988;
wire            n989;
wire            n990;
wire            n991;
wire            n992;
wire            n993;
wire            n994;
wire            n995;
wire            n996;
wire            n997;
wire            n998;
wire            n999;
wire            n1000;
wire            n1001;
wire            n1002;
wire            n1003;
wire            n1004;
wire            n1005;
wire            n1006;
wire            n1007;
wire            n1008;
wire            n1009;
wire            n1010;
wire            n1011;
wire            n1012;
wire            n1013;
wire            n1014;
wire            n1015;
wire            n1016;
wire            n1017;
wire            n1018;
wire            n1019;
wire            n1020;
wire            n1021;
wire            n1022;
wire            n1023;
wire            n1024;
wire            n1025;
wire            n1026;
wire            n1027;
wire            n1028;
wire            n1029;
wire            n1030;
wire            n1031;
wire            n1032;
wire            n1033;
wire            n1034;
wire            n1035;
wire            n1036;
wire            n1037;
wire            n1038;
wire            n1039;
wire            n1040;
wire            n1041;
wire            n1042;
wire            n1043;
wire            n1044;
wire            n1045;
wire            n1046;
wire            n1047;
wire            n1048;
wire            n1049;
wire            n1050;
wire            n1051;
wire            n1052;
wire            n1053;
wire            n1054;
wire            n1055;
wire            n1056;
wire            n1057;
wire            n1058;
wire            n1059;
wire            n1060;
wire            n1061;
wire            n1062;
wire            n1063;
wire            n1064;
wire            n1065;
wire            n1066;
wire            n1067;
wire            n1068;
wire            n1069;
wire            n1070;
wire            n1071;
wire            n1072;
wire            n1073;
wire            n1074;
wire            n1075;
wire            n1076;
wire            n1077;
wire            n1078;
wire            n1079;
wire            n1080;
wire            n1081;
wire            n1082;
wire            n1083;
wire            n1084;
wire            n1085;
wire            n1086;
wire            n1087;
wire            n1088;
wire            n1089;
wire            n1090;
wire            n1091;
wire            n1092;
wire            n1093;
wire            n1094;
wire            n1095;
wire            n1096;
wire            n1097;
wire            n1098;
wire            n1099;
wire            n1100;
wire            n1101;
wire            n1102;
wire            n1103;
wire            n1104;
wire            n1105;
wire            n1106;
wire            n1107;
wire            n1108;
wire            n1109;
wire            n1110;
wire            n1111;
wire            n1112;
wire            n1113;
wire            n1114;
wire            n1115;
wire            n1116;
wire            n1117;
wire            n1118;
wire            n1119;
wire            n1120;
wire            n1121;
wire            n1122;
wire            n1123;
wire            n1124;
wire            n1125;
wire            n1126;
wire            n1127;
wire            n1128;
wire            n1129;
wire            n1130;
wire            n1131;
wire            n1132;
wire            n1133;
wire            n1134;
wire            n1135;
wire            n1136;
wire            n1137;
wire            n1138;
wire            n1139;
wire            n1140;
wire            n1141;
wire            n1142;
wire            n1143;
wire            n1144;
wire            n1145;
wire            n1146;
wire            n1147;
wire            n1148;
wire            n1149;
wire            n1150;
wire            n1151;
wire            n1152;
wire            n1153;
wire            n1154;
wire            n1155;
wire            n1156;
wire            n1157;
wire            n1158;
wire            n1159;
wire            n1160;
wire            n1161;
wire            n1162;
wire            n1163;
wire            n1164;
wire            n1165;
wire            n1166;
wire            n1167;
wire            n1168;
wire            n1169;
wire            n1170;
wire            n1171;
wire            n1172;
wire            n1173;
wire            n1174;
wire            n1175;
wire            n1176;
wire            n1177;
wire            n1178;
wire            n1179;
wire            n1180;
wire            n1181;
wire            n1182;
wire            n1183;
wire            n1184;
wire            n1185;
wire            n1186;
wire            n1187;
wire            n1188;
wire            n1189;
wire            n1190;
wire            n1191;
wire            n1192;
wire            n1193;
wire            n1194;
wire            n1195;
wire            n1196;
wire            n1197;
wire            n1198;
wire            n1199;
wire            n1200;
wire            n1201;
wire            n1202;
wire            n1203;
wire            n1204;
wire            n1205;
wire            n1206;
wire            n1207;
wire            n1208;
wire            n1209;
wire            n1210;
wire            n1211;
wire            n1212;
wire            n1213;
wire            n1214;
wire            n1215;
wire            n1216;
wire            n1217;
wire            n1218;
wire            n1219;
wire            n1220;
wire            n1221;
wire            n1222;
wire            n1223;
wire            n1224;
wire            n1225;
wire            n1226;
wire            n1227;
wire            n1228;
wire            n1229;
wire            n1230;
wire            n1231;
wire            n1232;
wire            n1233;
wire            n1234;
wire            n1235;
wire            n1236;
wire            n1237;
wire            n1238;
wire            n1239;
wire            n1240;
wire            n1241;
wire            n1242;
wire            n1243;
wire            n1244;
wire            n1245;
wire            n1246;
wire            n1247;
wire            n1248;
wire            n1249;
wire            n1250;
wire            n1251;
wire            n1252;
wire            n1253;
wire            n1254;
wire            n1255;
wire            n1256;
wire            n1257;
wire            n1258;
wire            n1259;
wire            n1260;
wire            n1261;
wire            n1262;
wire            n1263;
wire            n1264;
wire            n1265;
wire            n1266;
wire            n1267;
wire            n1268;
wire            n1269;
wire            n1270;
wire            n1271;
wire            n1272;
wire            n1273;
wire            n1274;
wire            n1275;
wire            n1276;
wire            n1277;
wire            n1278;
wire            n1279;
wire            n1280;
wire            n1281;
wire            n1282;
wire            n1283;
wire            n1284;
wire            n1285;
wire            n1286;
wire            n1287;
wire            n1288;
wire            n1289;
wire            n1290;
wire            n1291;
wire            n1292;
wire            n1293;
wire            n1294;
wire            n1295;
wire            n1296;
wire            n1297;
wire            n1298;
wire            n1299;
wire            n1300;
wire            n1301;
wire            n1302;
wire            n1303;
wire            n1304;
wire            n1305;
wire            n1306;
wire            n1307;
wire            n1308;
wire            n1309;
wire            n1310;
wire            n1311;
wire            n1312;
wire            n1313;
wire            n1314;
wire            n1315;
wire            n1316;
wire            n1317;
wire            n1318;
wire            n1319;
wire            n1320;
wire            n1321;
wire            n1322;
wire            n1323;
wire            n1324;
wire            n1325;
wire            n1326;
wire            n1327;
wire            n1328;
wire            n1329;
wire            n1330;
wire            n1331;
wire            n1332;
wire            n1333;
wire            n1334;
wire            n1335;
wire            n1336;
wire            n1337;
wire            n1338;
wire            n1339;
wire            n1340;
wire            n1341;
wire            n1342;
wire            n1343;
wire            n1344;
wire            n1345;
wire            n1346;
wire            n1347;
wire            n1348;
wire            n1349;
wire            n1350;
wire            n1351;
wire            n1352;
wire            n1353;
wire            n1354;
wire            n1355;
wire            n1356;
wire            n1357;
wire            n1358;
wire            n1359;
wire            n1360;
wire            n1361;
wire            n1362;
wire            n1363;
wire            n1364;
wire            n1365;
wire            n1366;
wire            n1367;
wire            n1368;
wire            n1369;
wire            n1370;
wire            n1371;
wire            n1372;
wire            n1373;
wire            n1374;
wire            n1375;
wire            n1376;
wire            n1377;
wire            n1378;
wire            n1379;
wire            n1380;
wire            n1381;
wire            n1382;
wire            n1383;
wire            n1384;
wire            n1385;
wire            n1386;
wire            n1387;
wire            n1388;
wire            n1389;
wire            n1390;
wire            n1391;
wire            n1392;
wire            n1393;
wire            n1394;
wire            n1395;
wire            n1396;
wire            n1397;
wire            n1398;
wire            n1399;
wire            n1400;
wire            n1401;
wire            n1402;
wire            n1403;
wire            n1404;
wire            n1405;
wire            n1406;
wire            n1407;
wire     [31:0] n1408;
wire     [31:0] n1409;
wire     [31:0] n1410;
wire     [31:0] n1411;
wire     [31:0] n1412;
wire     [31:0] n1413;
wire     [31:0] n1414;
wire     [31:0] n1415;
wire     [31:0] n1416;
wire     [31:0] n1417;
wire     [31:0] n1418;
wire     [31:0] n1419;
wire     [31:0] n1420;
wire     [31:0] n1421;
wire     [31:0] n1422;
wire     [31:0] n1423;
wire     [31:0] n1424;
wire     [31:0] n1425;
wire     [31:0] n1426;
wire     [31:0] n1427;
wire     [31:0] n1428;
wire     [31:0] n1429;
wire     [31:0] n1430;
wire     [31:0] n1431;
wire     [31:0] n1432;
wire     [31:0] n1433;
wire     [31:0] n1434;
wire     [31:0] n1435;
wire     [31:0] n1436;
wire     [31:0] n1437;
wire     [31:0] n1438;
wire     [31:0] n1439;
wire     [31:0] n1440;
wire     [31:0] n1441;
wire     [31:0] n1442;
wire     [31:0] n1443;
wire     [31:0] n1444;
wire     [31:0] n1445;
wire     [31:0] n1446;
wire     [31:0] n1447;
wire     [31:0] n1448;
wire     [31:0] n1449;
wire     [31:0] n1450;
wire     [31:0] n1451;
wire     [31:0] n1452;
wire     [31:0] n1453;
wire     [31:0] n1454;
wire     [31:0] n1455;
wire     [31:0] n1456;
wire     [31:0] n1457;
wire     [31:0] n1458;
wire     [31:0] n1459;
wire     [31:0] n1460;
wire     [31:0] n1461;
wire     [31:0] n1462;
wire     [31:0] n1463;
wire     [31:0] n1464;
wire     [31:0] n1465;
wire     [31:0] n1466;
wire     [31:0] n1467;
wire     [31:0] n1468;
wire     [31:0] n1469;
wire     [31:0] n1470;
wire     [31:0] n1471;
wire     [31:0] n1472;
wire     [31:0] n1473;
wire     [31:0] n1474;
wire     [31:0] n1475;
wire     [31:0] n1476;
wire     [31:0] n1477;
wire     [31:0] n1478;
wire     [31:0] n1479;
wire     [31:0] n1480;
wire     [31:0] n1481;
wire     [31:0] n1482;
wire     [31:0] n1483;
wire     [31:0] n1484;
wire     [31:0] n1485;
wire     [31:0] n1486;
wire     [31:0] n1487;
wire     [31:0] n1488;
wire     [31:0] n1489;
wire     [31:0] n1490;
wire     [31:0] n1491;
wire     [31:0] n1492;
wire     [31:0] n1493;
wire     [31:0] n1494;
wire     [31:0] n1495;
wire     [31:0] n1496;
wire     [31:0] n1497;
wire     [31:0] n1498;
wire     [31:0] n1499;
wire     [31:0] n1500;
wire     [31:0] n1501;
wire     [31:0] n1502;
wire     [31:0] n1503;
wire     [31:0] n1504;
wire     [31:0] n1505;
wire     [31:0] n1506;
wire     [31:0] n1507;
wire     [31:0] n1508;
wire     [31:0] n1509;
wire     [31:0] n1510;
wire     [31:0] n1511;
wire     [31:0] n1512;
wire     [31:0] n1513;
wire     [31:0] n1514;
wire     [31:0] n1515;
wire     [31:0] n1516;
wire     [31:0] n1517;
wire     [31:0] n1518;
wire     [31:0] n1519;
wire     [31:0] n1520;
wire     [31:0] n1521;
wire     [31:0] n1522;
wire     [31:0] n1523;
wire     [31:0] n1524;
wire     [31:0] n1525;
wire     [31:0] n1526;
wire     [31:0] n1527;
wire     [31:0] n1528;
wire     [31:0] n1529;
wire     [31:0] n1530;
wire     [31:0] n1531;
wire     [31:0] n1532;
wire     [31:0] n1533;
wire     [31:0] n1534;
wire     [31:0] n1535;
wire     [31:0] n1536;
wire     [31:0] n1537;
wire     [31:0] n1538;
wire     [31:0] n1539;
wire     [31:0] n1540;
wire     [31:0] n1541;
wire     [31:0] n1542;
wire     [31:0] n1543;
wire     [31:0] n1544;
wire     [31:0] n1545;
wire     [31:0] n1546;
wire     [31:0] n1547;
wire     [31:0] n1548;
wire     [31:0] n1549;
wire     [31:0] n1550;
wire     [31:0] n1551;
wire     [31:0] n1552;
wire     [31:0] n1553;
wire     [31:0] n1554;
wire     [31:0] n1555;
wire     [31:0] n1556;
wire     [31:0] n1557;
wire     [31:0] n1558;
wire     [31:0] n1559;
wire     [31:0] n1560;
wire     [31:0] n1561;
wire     [31:0] n1562;
wire     [31:0] n1563;
wire     [31:0] n1564;
wire     [31:0] n1565;
wire     [31:0] n1566;
wire     [31:0] n1567;
wire     [31:0] n1568;
wire     [31:0] n1569;
wire     [31:0] n1570;
wire     [31:0] n1571;
wire     [31:0] n1572;
wire     [31:0] n1573;
wire     [31:0] n1574;
wire     [31:0] n1575;
wire     [31:0] n1576;
wire     [31:0] n1577;
wire     [31:0] n1578;
wire     [31:0] n1579;
wire     [31:0] n1580;
wire     [31:0] n1581;
wire     [31:0] n1582;
wire     [31:0] n1583;
wire     [31:0] n1584;
wire     [31:0] n1585;
wire     [31:0] n1586;
wire     [31:0] n1587;
wire     [31:0] n1588;
wire     [31:0] n1589;
wire     [31:0] n1590;
wire     [31:0] n1591;
wire     [31:0] n1592;
wire     [31:0] n1593;
wire     [31:0] n1594;
wire     [31:0] n1595;
wire     [31:0] n1596;
wire     [31:0] n1597;
wire     [31:0] n1598;
wire     [31:0] n1599;
wire     [31:0] n1600;
wire     [31:0] n1601;
wire     [31:0] n1602;
wire     [31:0] n1603;
wire     [31:0] n1604;
wire     [31:0] n1605;
wire     [31:0] n1606;
wire     [31:0] n1607;
wire     [31:0] n1608;
wire     [31:0] n1609;
wire     [31:0] n1610;
wire     [31:0] n1611;
wire     [31:0] n1612;
wire     [31:0] n1613;
wire     [31:0] n1614;
wire     [31:0] n1615;
wire     [31:0] n1616;
wire     [31:0] n1617;
wire     [31:0] n1618;
wire     [31:0] n1619;
wire     [31:0] n1620;
wire     [31:0] n1621;
wire     [31:0] n1622;
wire     [31:0] n1623;
wire     [31:0] n1624;
wire     [31:0] n1625;
wire     [31:0] n1626;
wire     [31:0] n1627;
wire     [31:0] n1628;
wire     [31:0] n1629;
wire     [31:0] n1630;
wire     [31:0] n1631;
wire     [31:0] n1632;
wire     [31:0] n1633;
wire     [31:0] n1634;
wire     [31:0] n1635;
wire     [31:0] n1636;
wire     [31:0] n1637;
wire     [31:0] n1638;
wire     [31:0] n1639;
wire     [31:0] n1640;
wire     [31:0] n1641;
wire     [31:0] n1642;
wire     [31:0] n1643;
wire     [31:0] n1644;
wire     [31:0] n1645;
wire     [31:0] n1646;
wire     [31:0] n1647;
wire     [31:0] n1648;
wire     [31:0] n1649;
wire     [31:0] n1650;
wire     [31:0] n1651;
wire     [31:0] n1652;
wire     [31:0] n1653;
wire     [31:0] n1654;
wire     [31:0] n1655;
wire     [31:0] n1656;
wire     [31:0] n1657;
wire     [31:0] n1658;
wire     [31:0] n1659;
wire     [31:0] n1660;
wire     [31:0] n1661;
wire     [31:0] n1662;
wire     [31:0] n1663;
wire     [31:0] n1664;
wire     [31:0] n1665;
wire     [31:0] n1666;
wire     [31:0] n1667;
wire     [31:0] n1668;
wire     [31:0] n1669;
wire     [31:0] n1670;
wire     [31:0] n1671;
wire     [31:0] n1672;
wire     [31:0] n1673;
wire     [31:0] n1674;
wire     [31:0] n1675;
wire     [31:0] n1676;
wire     [31:0] n1677;
wire     [31:0] n1678;
wire     [31:0] n1679;
wire     [31:0] n1680;
wire     [31:0] n1681;
wire     [31:0] n1682;
wire     [31:0] n1683;
wire     [31:0] n1684;
wire     [31:0] n1685;
wire     [31:0] n1686;
wire     [31:0] n1687;
wire     [31:0] n1688;
wire     [31:0] n1689;
wire     [31:0] n1690;
wire     [31:0] n1691;
wire     [31:0] n1692;
wire     [31:0] n1693;
wire     [31:0] n1694;
wire     [31:0] n1695;
wire     [31:0] n1696;
wire     [31:0] n1697;
wire     [31:0] n1698;
wire     [31:0] n1699;
wire     [31:0] n1700;
wire     [31:0] n1701;
wire     [31:0] n1702;
wire     [31:0] n1703;
wire     [31:0] n1704;
wire     [31:0] n1705;
wire     [31:0] n1706;
wire     [31:0] n1707;
wire     [31:0] n1708;
wire     [31:0] n1709;
wire     [31:0] n1710;
wire     [31:0] n1711;
wire     [31:0] n1712;
wire     [31:0] n1713;
wire     [31:0] n1714;
wire     [31:0] n1715;
wire     [31:0] n1716;
wire     [31:0] n1717;
wire     [31:0] n1718;
wire     [31:0] n1719;
wire     [31:0] n1720;
wire     [31:0] n1721;
wire     [31:0] n1722;
wire     [31:0] n1723;
wire     [31:0] n1724;
wire     [31:0] n1725;
wire     [31:0] n1726;
wire     [31:0] n1727;
wire     [31:0] n1728;
wire     [31:0] n1729;
wire     [31:0] n1730;
wire     [31:0] n1731;
wire     [31:0] n1732;
wire     [31:0] n1733;
wire     [31:0] n1734;
wire     [31:0] n1735;
wire     [31:0] n1736;
wire     [31:0] n1737;
wire     [31:0] n1738;
wire     [31:0] n1739;
wire     [31:0] n1740;
wire     [31:0] n1741;
wire     [31:0] n1742;
wire     [31:0] n1743;
wire     [31:0] n1744;
wire     [31:0] n1745;
wire     [31:0] n1746;
wire     [31:0] n1747;
wire     [31:0] n1748;
wire     [31:0] n1749;
wire     [31:0] n1750;
wire     [31:0] n1751;
wire     [31:0] n1752;
wire     [31:0] n1753;
wire     [31:0] n1754;
wire     [31:0] n1755;
wire     [31:0] n1756;
wire     [31:0] n1757;
wire     [31:0] n1758;
wire     [31:0] n1759;
wire     [31:0] n1760;
wire     [31:0] n1761;
wire     [31:0] n1762;
wire     [31:0] n1763;
wire     [31:0] n1764;
wire     [31:0] n1765;
wire     [31:0] n1766;
wire     [31:0] n1767;
wire     [31:0] n1768;
wire     [31:0] n1769;
wire     [31:0] n1770;
wire     [31:0] n1771;
wire     [31:0] n1772;
wire     [31:0] n1773;
wire     [31:0] n1774;
wire     [31:0] n1775;
wire     [31:0] n1776;
wire     [31:0] n1777;
wire     [31:0] n1778;
wire     [31:0] n1779;
wire     [31:0] n1780;
wire     [31:0] n1781;
wire     [31:0] n1782;
wire     [31:0] n1783;
wire     [31:0] n1784;
wire     [31:0] n1785;
wire     [31:0] n1786;
wire     [31:0] n1787;
wire     [31:0] n1788;
wire     [31:0] n1789;
wire     [31:0] n1790;
wire     [31:0] n1791;
wire     [31:0] n1792;
wire     [31:0] n1793;
wire     [31:0] n1794;
wire     [31:0] n1795;
wire     [31:0] n1796;
wire     [31:0] n1797;
wire     [31:0] n1798;
wire     [31:0] n1799;
wire     [31:0] n1800;
wire     [31:0] n1801;
wire     [31:0] n1802;
wire     [31:0] n1803;
wire     [31:0] n1804;
wire     [31:0] n1805;
wire     [31:0] n1806;
wire     [31:0] n1807;
wire     [31:0] n1808;
wire     [31:0] n1809;
wire     [31:0] n1810;
wire     [31:0] n1811;
wire     [31:0] n1812;
wire     [31:0] n1813;
wire     [31:0] n1814;
wire     [31:0] n1815;
wire     [31:0] n1816;
wire     [31:0] n1817;
wire     [31:0] n1818;
wire     [31:0] n1819;
wire     [31:0] n1820;
wire     [31:0] n1821;
wire     [31:0] n1822;
wire     [31:0] n1823;
wire     [31:0] n1824;
wire     [31:0] n1825;
wire     [31:0] n1826;
wire     [31:0] n1827;
wire     [31:0] n1828;
wire     [31:0] n1829;
wire     [31:0] n1830;
wire     [31:0] n1831;
wire     [31:0] n1832;
wire     [31:0] n1833;
wire     [31:0] n1834;
wire     [31:0] n1835;
wire     [31:0] n1836;
wire     [31:0] n1837;
wire     [31:0] n1838;
wire     [31:0] n1839;
wire     [31:0] n1840;
wire     [31:0] n1841;
wire     [31:0] n1842;
wire     [31:0] n1843;
wire     [31:0] n1844;
wire     [31:0] n1845;
wire     [31:0] n1846;
wire     [31:0] n1847;
wire     [31:0] n1848;
wire     [31:0] n1849;
wire     [31:0] n1850;
wire     [31:0] n1851;
wire     [31:0] n1852;
wire     [31:0] n1853;
wire     [31:0] n1854;
wire     [31:0] n1855;
wire     [31:0] n1856;
wire     [31:0] n1857;
wire     [31:0] n1858;
wire     [31:0] n1859;
wire     [31:0] n1860;
wire     [31:0] n1861;
wire     [31:0] n1862;
wire     [31:0] n1863;
wire     [31:0] n1864;
wire     [31:0] n1865;
wire     [31:0] n1866;
wire     [31:0] n1867;
wire     [31:0] n1868;
wire     [31:0] n1869;
wire     [31:0] n1870;
wire     [31:0] n1871;
wire     [31:0] n1872;
wire     [31:0] n1873;
wire     [31:0] n1874;
wire     [31:0] n1875;
wire     [31:0] n1876;
wire     [31:0] n1877;
wire     [31:0] n1878;
wire     [31:0] n1879;
wire     [31:0] n1880;
wire     [31:0] n1881;
wire     [31:0] n1882;
wire     [31:0] n1883;
wire     [31:0] n1884;
wire     [31:0] n1885;
wire     [31:0] n1886;
wire     [31:0] n1887;
wire     [31:0] n1888;
wire     [31:0] n1889;
wire     [31:0] n1890;
wire     [31:0] n1891;
wire     [31:0] n1892;
wire     [31:0] n1893;
wire     [31:0] n1894;
wire     [31:0] n1895;
wire     [31:0] n1896;
wire     [31:0] n1897;
wire     [31:0] n1898;
wire     [31:0] n1899;
wire     [31:0] n1900;
wire     [31:0] n1901;
wire     [31:0] n1902;
wire     [31:0] n1903;
wire     [31:0] n1904;
wire     [31:0] n1905;
wire     [31:0] n1906;
wire     [31:0] n1907;
wire     [31:0] n1908;
wire     [31:0] n1909;
wire     [31:0] n1910;
wire     [31:0] n1911;
wire     [31:0] n1912;
wire     [31:0] n1913;
wire     [31:0] n1914;
wire     [31:0] n1915;
wire     [31:0] n1916;
wire     [31:0] n1917;
wire     [31:0] n1918;
wire     [31:0] n1919;
wire     [31:0] n1920;
wire     [31:0] n1921;
wire     [31:0] n1922;
wire     [31:0] n1923;
wire     [31:0] n1924;
wire     [31:0] n1925;
wire     [31:0] n1926;
wire     [31:0] n1927;
wire     [31:0] n1928;
wire     [31:0] n1929;
wire            n1930;
wire            n1931;
wire            n1932;
wire            n1933;
wire            n1934;
wire            n1935;
wire            n1936;
wire            n1937;
wire            n1938;
wire            n1939;
wire            n1940;
wire            n1941;
wire            n1942;
wire            n1943;
wire            n1944;
wire            n1945;
wire            n1946;
wire            n1947;
wire            n1948;
wire            n1949;
wire            n1950;
wire            n1951;
wire            n1952;
wire            n1953;
wire            n1954;
wire            n1955;
wire            n1956;
wire            n1957;
wire            n1958;
wire            n1959;
wire            n1960;
wire            n1961;
wire            n1962;
wire            n1963;
wire            n1964;
wire            n1965;
wire            n1966;
wire            n1967;
wire            n1968;
wire            n1969;
wire            n1970;
wire            n1971;
wire            n1972;
wire            n1973;
wire            n1974;
wire            n1975;
wire            n1976;
wire            n1977;
wire            n1978;
wire            n1979;
wire            n1980;
wire            n1981;
wire            n1982;
wire            n1983;
wire            n1984;
wire            n1985;
wire            n1986;
wire            n1987;
wire            n1988;
wire            n1989;
wire            n1990;
wire            n1991;
wire            n1992;
wire            n1993;
wire            n1994;
wire            n1995;
wire            n1996;
wire            n1997;
wire            n1998;
wire            n1999;
wire            n2000;
wire            n2001;
wire            n2002;
wire            n2003;
wire            n2004;
wire            n2005;
wire            n2006;
wire            n2007;
wire            n2008;
wire            n2009;
wire            n2010;
wire            n2011;
wire            n2012;
wire            n2013;
wire            n2014;
wire            n2015;
wire            n2016;
wire            n2017;
wire            n2018;
wire            n2019;
wire            n2020;
wire            n2021;
wire            n2022;
wire            n2023;
wire            n2024;
wire            n2025;
wire            n2026;
wire            n2027;
wire            n2028;
wire            n2029;
wire            n2030;
wire            n2031;
wire            n2032;
wire            n2033;
wire            n2034;
wire            n2035;
wire            n2036;
wire            n2037;
wire            n2038;
wire            n2039;
wire            n2040;
wire            n2041;
wire            n2042;
wire            n2043;
wire            n2044;
wire            n2045;
wire            n2046;
wire            n2047;
wire            n2048;
wire            n2049;
wire            n2050;
wire            n2051;
wire            n2052;
wire            n2053;
wire            n2054;
wire            n2055;
wire            n2056;
wire            n2057;
wire            n2058;
wire            n2059;
wire            n2060;
wire            n2061;
wire            n2062;
wire            n2063;
wire            n2064;
wire            n2065;
wire            n2066;
wire            n2067;
wire            n2068;
wire            n2069;
wire            n2070;
wire            n2071;
wire            n2072;
wire            n2073;
wire            n2074;
wire            n2075;
wire            n2076;
wire            n2077;
wire            n2078;
wire            n2079;
wire            n2080;
wire            n2081;
wire            n2082;
wire            n2083;
wire            n2084;
wire            n2085;
wire            n2086;
wire            n2087;
wire            n2088;
wire            n2089;
wire            n2090;
wire            n2091;
wire            n2092;
wire            n2093;
wire            n2094;
wire            n2095;
wire            n2096;
wire            n2097;
wire            n2098;
wire            n2099;
wire            n2100;
wire            n2101;
wire            n2102;
wire            n2103;
wire            n2104;
wire            n2105;
wire            n2106;
wire            n2107;
wire            n2108;
wire            n2109;
wire            n2110;
wire            n2111;
wire            n2112;
wire            n2113;
wire            n2114;
wire            n2115;
wire            n2116;
wire            n2117;
wire            n2118;
wire            n2119;
wire            n2120;
wire            n2121;
wire            n2122;
wire            n2123;
wire            n2124;
wire            n2125;
wire            n2126;
wire            n2127;
wire            n2128;
wire            n2129;
wire            n2130;
wire            n2131;
wire            n2132;
wire            n2133;
wire            n2134;
wire            n2135;
wire            n2136;
wire            n2137;
wire            n2138;
wire            n2139;
wire            n2140;
wire            n2141;
wire            n2142;
wire            n2143;
wire            n2144;
wire            n2145;
wire            n2146;
wire            n2147;
wire            n2148;
wire            n2149;
wire            n2150;
wire            n2151;
wire            n2152;
wire            n2153;
wire            n2154;
wire            n2155;
wire            n2156;
wire            n2157;
wire            n2158;
wire            n2159;
wire            n2160;
wire            n2161;
wire            n2162;
wire            n2163;
wire            n2164;
wire            n2165;
wire            n2166;
wire            n2167;
wire            n2168;
wire            n2169;
wire            n2170;
wire            n2171;
wire            n2172;
wire            n2173;
wire            n2174;
wire            n2175;
wire            n2176;
wire            n2177;
wire            n2178;
wire            n2179;
wire            n2180;
wire            n2181;
wire            n2182;
wire            n2183;
wire            n2184;
wire            n2185;
wire            n2186;
wire            n2187;
wire            n2188;
wire            n2189;
wire            n2190;
wire            n2191;
wire            n2192;
wire            n2193;
wire            n2194;
wire            n2195;
wire            n2196;
wire            n2197;
wire            n2198;
wire            n2199;
wire            n2200;
wire            n2201;
wire            n2202;
wire            n2203;
wire            n2204;
wire            n2205;
wire            n2206;
wire            n2207;
wire            n2208;
wire            n2209;
wire            n2210;
wire            n2211;
wire            n2212;
wire            n2213;
wire            n2214;
wire            n2215;
wire            n2216;
wire            n2217;
wire            n2218;
wire            n2219;
wire            n2220;
wire            n2221;
wire            n2222;
wire            n2223;
wire            n2224;
wire            n2225;
wire            n2226;
wire            n2227;
wire            n2228;
wire            n2229;
wire            n2230;
wire            n2231;
wire            n2232;
wire            n2233;
wire            n2234;
wire            n2235;
wire            n2236;
wire            n2237;
wire            n2238;
wire            n2239;
wire            n2240;
wire            n2241;
wire            n2242;
wire            n2243;
wire            n2244;
wire            n2245;
wire            n2246;
wire            n2247;
wire            n2248;
wire            n2249;
wire            n2250;
wire            n2251;
wire            n2252;
wire            n2253;
wire            n2254;
wire            n2255;
wire            n2256;
wire            n2257;
wire            n2258;
wire            n2259;
wire            n2260;
wire            n2261;
wire            n2262;
wire            n2263;
wire            n2264;
wire            n2265;
wire            n2266;
wire            n2267;
wire            n2268;
wire            n2269;
wire            n2270;
wire            n2271;
wire            n2272;
wire            n2273;
wire            n2274;
wire            n2275;
wire            n2276;
wire            n2277;
wire            n2278;
wire            n2279;
wire            n2280;
wire            n2281;
wire            n2282;
wire            n2283;
wire            n2284;
wire            n2285;
wire            n2286;
wire            n2287;
wire            n2288;
wire            n2289;
wire            n2290;
wire            n2291;
wire            n2292;
wire            n2293;
wire            n2294;
wire            n2295;
wire            n2296;
wire            n2297;
wire            n2298;
wire            n2299;
wire            n2300;
wire            n2301;
wire            n2302;
wire            n2303;
wire            n2304;
wire            n2305;
wire            n2306;
wire            n2307;
wire            n2308;
wire            n2309;
wire            n2310;
wire            n2311;
wire            n2312;
wire            n2313;
wire            n2314;
wire            n2315;
wire            n2316;
wire            n2317;
wire            n2318;
wire            n2319;
wire            n2320;
wire            n2321;
wire            n2322;
wire            n2323;
wire            n2324;
wire            n2325;
wire            n2326;
wire            n2327;
wire            n2328;
wire            n2329;
wire            n2330;
wire            n2331;
wire            n2332;
wire            n2333;
wire            n2334;
wire            n2335;
wire            n2336;
wire            n2337;
wire            n2338;
wire            n2339;
wire            n2340;
wire            n2341;
wire            n2342;
wire            n2343;
wire            n2344;
wire            n2345;
wire            n2346;
wire            n2347;
wire            n2348;
wire            n2349;
wire            n2350;
wire            n2351;
wire            n2352;
wire            n2353;
wire            n2354;
wire            n2355;
wire            n2356;
wire            n2357;
wire            n2358;
wire            n2359;
wire            n2360;
wire            n2361;
wire            n2362;
wire            n2363;
wire            n2364;
wire            n2365;
wire            n2366;
wire            n2367;
wire            n2368;
wire            n2369;
wire            n2370;
wire            n2371;
wire            n2372;
wire            n2373;
wire            n2374;
wire            n2375;
wire            n2376;
wire            n2377;
wire            n2378;
wire            n2379;
wire            n2380;
wire            n2381;
wire            n2382;
wire            n2383;
wire            n2384;
wire            n2385;
wire            n2386;
wire            n2387;
wire            n2388;
wire            n2389;
wire            n2390;
wire            n2391;
wire            n2392;
wire            n2393;
wire            n2394;
wire            n2395;
wire            n2396;
wire            n2397;
wire            n2398;
wire            n2399;
wire            n2400;
wire            n2401;
wire            n2402;
wire            n2403;
wire            n2404;
wire            n2405;
wire            n2406;
wire            n2407;
wire            n2408;
wire            n2409;
wire            n2410;
wire            n2411;
wire            n2412;
wire            n2413;
wire            n2414;
wire            n2415;
wire            n2416;
wire            n2417;
wire            n2418;
wire            n2419;
wire            n2420;
wire            n2421;
wire            n2422;
wire            n2423;
wire            n2424;
wire            n2425;
wire            n2426;
wire            n2427;
wire            n2428;
wire            n2429;
wire            n2430;
wire            n2431;
wire            n2432;
wire            n2433;
wire            n2434;
wire            n2435;
wire            n2436;
wire            n2437;
wire            n2438;
wire            n2439;
wire            n2440;
wire            n2441;
wire            n2442;
wire     [31:0] n2443;
wire     [31:0] n2444;
wire     [31:0] n2445;
wire     [31:0] n2446;
wire     [31:0] n2447;
wire     [31:0] n2448;
wire     [31:0] n2449;
wire     [31:0] n2450;
wire     [31:0] n2451;
wire     [31:0] n2452;
wire     [31:0] n2453;
wire     [31:0] n2454;
wire     [31:0] n2455;
wire     [31:0] n2456;
wire     [31:0] n2457;
wire     [31:0] n2458;
wire     [31:0] n2459;
wire     [31:0] n2460;
wire     [31:0] n2461;
wire     [31:0] n2462;
wire     [31:0] n2463;
wire     [31:0] n2464;
wire     [31:0] n2465;
wire     [31:0] n2466;
wire     [31:0] n2467;
wire     [31:0] n2468;
wire     [31:0] n2469;
wire     [31:0] n2470;
wire     [31:0] n2471;
wire     [31:0] n2472;
wire     [31:0] n2473;
wire     [31:0] n2474;
wire     [31:0] n2475;
wire     [31:0] n2476;
wire     [31:0] n2477;
wire     [31:0] n2478;
wire     [31:0] n2479;
wire     [31:0] n2480;
wire     [31:0] n2481;
wire     [31:0] n2482;
wire     [31:0] n2483;
wire     [31:0] n2484;
wire     [31:0] n2485;
wire     [31:0] n2486;
wire     [31:0] n2487;
wire     [31:0] n2488;
wire     [31:0] n2489;
wire     [31:0] n2490;
wire     [31:0] n2491;
wire     [31:0] n2492;
wire     [31:0] n2493;
wire     [31:0] n2494;
wire     [31:0] n2495;
wire     [31:0] n2496;
wire     [31:0] n2497;
wire     [31:0] n2498;
wire     [31:0] n2499;
wire     [31:0] n2500;
wire     [31:0] n2501;
wire     [31:0] n2502;
wire     [31:0] n2503;
wire     [31:0] n2504;
wire     [31:0] n2505;
wire     [31:0] n2506;
wire     [31:0] n2507;
wire     [31:0] n2508;
wire     [31:0] n2509;
wire     [31:0] n2510;
wire     [31:0] n2511;
wire     [31:0] n2512;
wire     [31:0] n2513;
wire     [31:0] n2514;
wire     [31:0] n2515;
wire     [31:0] n2516;
wire     [31:0] n2517;
wire     [31:0] n2518;
wire     [31:0] n2519;
wire     [31:0] n2520;
wire     [31:0] n2521;
wire     [31:0] n2522;
wire     [31:0] n2523;
wire     [31:0] n2524;
wire     [31:0] n2525;
wire     [31:0] n2526;
wire     [31:0] n2527;
wire     [31:0] n2528;
wire     [31:0] n2529;
wire     [31:0] n2530;
wire     [31:0] n2531;
wire     [31:0] n2532;
wire     [31:0] n2533;
wire     [31:0] n2534;
wire     [31:0] n2535;
wire     [31:0] n2536;
wire     [31:0] n2537;
wire     [31:0] n2538;
wire     [31:0] n2539;
wire     [31:0] n2540;
wire     [31:0] n2541;
wire     [31:0] n2542;
wire     [31:0] n2543;
wire     [31:0] n2544;
wire     [31:0] n2545;
wire     [31:0] n2546;
wire     [31:0] n2547;
wire     [31:0] n2548;
wire     [31:0] n2549;
wire     [31:0] n2550;
wire     [31:0] n2551;
wire     [31:0] n2552;
wire     [31:0] n2553;
wire     [31:0] n2554;
wire     [31:0] n2555;
wire     [31:0] n2556;
wire     [31:0] n2557;
wire     [31:0] n2558;
wire     [31:0] n2559;
wire     [31:0] n2560;
wire     [31:0] n2561;
wire     [31:0] n2562;
wire     [31:0] n2563;
wire     [31:0] n2564;
wire     [31:0] n2565;
wire     [31:0] n2566;
wire     [31:0] n2567;
wire     [31:0] n2568;
wire     [31:0] n2569;
wire     [31:0] n2570;
wire     [31:0] n2571;
wire     [31:0] n2572;
wire     [31:0] n2573;
wire     [31:0] n2574;
wire     [31:0] n2575;
wire     [31:0] n2576;
wire     [31:0] n2577;
wire     [31:0] n2578;
wire     [31:0] n2579;
wire     [31:0] n2580;
wire     [31:0] n2581;
wire     [31:0] n2582;
wire     [31:0] n2583;
wire     [31:0] n2584;
wire     [31:0] n2585;
wire     [31:0] n2586;
wire     [31:0] n2587;
wire     [31:0] n2588;
wire     [31:0] n2589;
wire     [31:0] n2590;
wire     [31:0] n2591;
wire     [31:0] n2592;
wire     [31:0] n2593;
wire     [31:0] n2594;
wire     [31:0] n2595;
wire     [31:0] n2596;
wire     [31:0] n2597;
wire     [31:0] n2598;
wire     [31:0] n2599;
wire     [31:0] n2600;
wire     [31:0] n2601;
wire     [31:0] n2602;
wire     [31:0] n2603;
wire     [31:0] n2604;
wire     [31:0] n2605;
wire     [31:0] n2606;
wire     [31:0] n2607;
wire     [31:0] n2608;
wire     [31:0] n2609;
wire     [31:0] n2610;
wire     [31:0] n2611;
wire     [31:0] n2612;
wire     [31:0] n2613;
wire     [31:0] n2614;
wire     [31:0] n2615;
wire     [31:0] n2616;
wire     [31:0] n2617;
wire     [31:0] n2618;
wire     [31:0] n2619;
wire     [31:0] n2620;
wire     [31:0] n2621;
wire     [31:0] n2622;
wire     [31:0] n2623;
wire     [31:0] n2624;
wire     [31:0] n2625;
wire     [31:0] n2626;
wire     [31:0] n2627;
wire     [31:0] n2628;
wire     [31:0] n2629;
wire     [31:0] n2630;
wire     [31:0] n2631;
wire     [31:0] n2632;
wire     [31:0] n2633;
wire     [31:0] n2634;
wire     [31:0] n2635;
wire     [31:0] n2636;
wire     [31:0] n2637;
wire     [31:0] n2638;
wire     [31:0] n2639;
wire     [31:0] n2640;
wire     [31:0] n2641;
wire     [31:0] n2642;
wire     [31:0] n2643;
wire     [31:0] n2644;
wire     [31:0] n2645;
wire     [31:0] n2646;
wire     [31:0] n2647;
wire     [31:0] n2648;
wire     [31:0] n2649;
wire     [31:0] n2650;
wire     [31:0] n2651;
wire     [31:0] n2652;
wire     [31:0] n2653;
wire     [31:0] n2654;
wire     [31:0] n2655;
wire     [31:0] n2656;
wire     [31:0] n2657;
wire     [31:0] n2658;
wire     [31:0] n2659;
wire     [31:0] n2660;
wire     [31:0] n2661;
wire     [31:0] n2662;
wire     [31:0] n2663;
wire     [31:0] n2664;
wire     [31:0] n2665;
wire     [31:0] n2666;
wire     [31:0] n2667;
wire     [31:0] n2668;
wire     [31:0] n2669;
wire     [31:0] n2670;
wire     [31:0] n2671;
wire     [31:0] n2672;
wire     [31:0] n2673;
wire     [31:0] n2674;
wire     [31:0] n2675;
wire     [31:0] n2676;
wire     [31:0] n2677;
wire     [31:0] n2678;
wire     [31:0] n2679;
wire     [31:0] n2680;
wire     [31:0] n2681;
wire     [31:0] n2682;
wire     [31:0] n2683;
wire     [31:0] n2684;
wire     [31:0] n2685;
wire     [31:0] n2686;
wire     [31:0] n2687;
wire     [31:0] n2688;
wire     [31:0] n2689;
wire     [31:0] n2690;
wire     [31:0] n2691;
wire     [31:0] n2692;
wire     [31:0] n2693;
wire     [31:0] n2694;
wire     [31:0] n2695;
wire     [31:0] n2696;
wire     [31:0] n2697;
wire     [31:0] n2698;
wire     [31:0] n2699;
wire     [31:0] n2700;
wire     [31:0] n2701;
wire     [31:0] n2702;
wire     [31:0] n2703;
wire     [31:0] n2704;
wire     [31:0] n2705;
wire     [31:0] n2706;
wire     [31:0] n2707;
wire     [31:0] n2708;
wire     [31:0] n2709;
wire     [31:0] n2710;
wire     [31:0] n2711;
wire     [31:0] n2712;
wire     [31:0] n2713;
wire     [31:0] n2714;
wire     [31:0] n2715;
wire     [31:0] n2716;
wire     [31:0] n2717;
wire     [31:0] n2718;
wire     [31:0] n2719;
wire     [31:0] n2720;
wire     [31:0] n2721;
wire     [31:0] n2722;
wire     [31:0] n2723;
wire     [31:0] n2724;
wire     [31:0] n2725;
wire     [31:0] n2726;
wire     [31:0] n2727;
wire     [31:0] n2728;
wire     [31:0] n2729;
wire     [31:0] n2730;
wire     [31:0] n2731;
wire     [31:0] n2732;
wire     [31:0] n2733;
wire     [31:0] n2734;
wire     [31:0] n2735;
wire     [31:0] n2736;
wire     [31:0] n2737;
wire     [31:0] n2738;
wire     [31:0] n2739;
wire     [31:0] n2740;
wire     [31:0] n2741;
wire     [31:0] n2742;
wire     [31:0] n2743;
wire     [31:0] n2744;
wire     [31:0] n2745;
wire     [31:0] n2746;
wire     [31:0] n2747;
wire     [31:0] n2748;
wire     [31:0] n2749;
wire     [31:0] n2750;
wire     [31:0] n2751;
wire     [31:0] n2752;
wire     [31:0] n2753;
wire     [31:0] n2754;
wire     [31:0] n2755;
wire     [31:0] n2756;
wire     [31:0] n2757;
wire     [31:0] n2758;
wire     [31:0] n2759;
wire     [31:0] n2760;
wire     [31:0] n2761;
wire     [31:0] n2762;
wire     [31:0] n2763;
wire     [31:0] n2764;
wire     [31:0] n2765;
wire     [31:0] n2766;
wire     [31:0] n2767;
wire     [31:0] n2768;
wire     [31:0] n2769;
wire     [31:0] n2770;
wire     [31:0] n2771;
wire     [31:0] n2772;
wire     [31:0] n2773;
wire     [31:0] n2774;
wire     [31:0] n2775;
wire     [31:0] n2776;
wire     [31:0] n2777;
wire     [31:0] n2778;
wire     [31:0] n2779;
wire     [31:0] n2780;
wire     [31:0] n2781;
wire     [31:0] n2782;
wire     [31:0] n2783;
wire     [31:0] n2784;
wire     [31:0] n2785;
wire     [31:0] n2786;
wire     [31:0] n2787;
wire     [31:0] n2788;
wire     [31:0] n2789;
wire     [31:0] n2790;
wire     [31:0] n2791;
wire     [31:0] n2792;
wire     [31:0] n2793;
wire     [31:0] n2794;
wire     [31:0] n2795;
wire     [31:0] n2796;
wire     [31:0] n2797;
wire     [31:0] n2798;
wire     [31:0] n2799;
wire     [31:0] n2800;
wire     [31:0] n2801;
wire     [31:0] n2802;
wire     [31:0] n2803;
wire     [31:0] n2804;
wire     [31:0] n2805;
wire     [31:0] n2806;
wire     [31:0] n2807;
wire     [31:0] n2808;
wire     [31:0] n2809;
wire     [31:0] n2810;
wire     [31:0] n2811;
wire     [31:0] n2812;
wire     [31:0] n2813;
wire     [31:0] n2814;
wire     [31:0] n2815;
wire     [31:0] n2816;
wire     [31:0] n2817;
wire     [31:0] n2818;
wire     [31:0] n2819;
wire     [31:0] n2820;
wire     [31:0] n2821;
wire     [31:0] n2822;
wire     [31:0] n2823;
wire     [31:0] n2824;
wire     [31:0] n2825;
wire     [31:0] n2826;
wire     [31:0] n2827;
wire     [31:0] n2828;
wire     [31:0] n2829;
wire     [31:0] n2830;
wire     [31:0] n2831;
wire     [31:0] n2832;
wire     [31:0] n2833;
wire     [31:0] n2834;
wire     [31:0] n2835;
wire     [31:0] n2836;
wire     [31:0] n2837;
wire     [31:0] n2838;
wire     [31:0] n2839;
wire     [31:0] n2840;
wire     [31:0] n2841;
wire     [31:0] n2842;
wire     [31:0] n2843;
wire     [31:0] n2844;
wire     [31:0] n2845;
wire     [31:0] n2846;
wire     [31:0] n2847;
wire     [31:0] n2848;
wire     [31:0] n2849;
wire     [31:0] n2850;
wire     [31:0] n2851;
wire     [31:0] n2852;
wire     [31:0] n2853;
wire     [31:0] n2854;
wire     [31:0] n2855;
wire     [31:0] n2856;
wire     [31:0] n2857;
wire     [31:0] n2858;
wire     [31:0] n2859;
wire     [31:0] n2860;
wire     [31:0] n2861;
wire     [31:0] n2862;
wire     [31:0] n2863;
wire     [31:0] n2864;
wire     [31:0] n2865;
wire     [31:0] n2866;
wire     [31:0] n2867;
wire     [31:0] n2868;
wire     [31:0] n2869;
wire     [31:0] n2870;
wire     [31:0] n2871;
wire     [31:0] n2872;
wire     [31:0] n2873;
wire     [31:0] n2874;
wire     [31:0] n2875;
wire     [31:0] n2876;
wire     [31:0] n2877;
wire     [31:0] n2878;
wire     [31:0] n2879;
wire     [31:0] n2880;
wire     [31:0] n2881;
wire     [31:0] n2882;
wire     [31:0] n2883;
wire     [31:0] n2884;
wire     [31:0] n2885;
wire     [31:0] n2886;
wire     [31:0] n2887;
wire     [31:0] n2888;
wire     [31:0] n2889;
wire     [31:0] n2890;
wire     [31:0] n2891;
wire     [31:0] n2892;
wire     [31:0] n2893;
wire     [31:0] n2894;
wire     [31:0] n2895;
wire     [31:0] n2896;
wire     [31:0] n2897;
wire     [31:0] n2898;
wire     [31:0] n2899;
wire     [31:0] n2900;
wire     [31:0] n2901;
wire     [31:0] n2902;
wire     [31:0] n2903;
wire     [31:0] n2904;
wire     [31:0] n2905;
wire     [31:0] n2906;
wire     [31:0] n2907;
wire     [31:0] n2908;
wire     [31:0] n2909;
wire     [31:0] n2910;
wire     [31:0] n2911;
wire     [31:0] n2912;
wire     [31:0] n2913;
wire     [31:0] n2914;
wire     [31:0] n2915;
wire     [31:0] n2916;
wire     [31:0] n2917;
wire     [31:0] n2918;
wire     [31:0] n2919;
wire     [31:0] n2920;
wire     [31:0] n2921;
wire     [31:0] n2922;
wire     [31:0] n2923;
wire     [31:0] n2924;
wire     [31:0] n2925;
wire     [31:0] n2926;
wire     [31:0] n2927;
wire     [31:0] n2928;
wire     [31:0] n2929;
wire     [31:0] n2930;
wire     [31:0] n2931;
wire     [31:0] n2932;
wire     [31:0] n2933;
wire     [31:0] n2934;
wire     [31:0] n2935;
wire     [31:0] n2936;
wire     [31:0] n2937;
wire     [31:0] n2938;
wire     [31:0] n2939;
wire     [31:0] n2940;
wire     [31:0] n2941;
wire     [31:0] n2942;
wire     [31:0] n2943;
wire     [31:0] n2944;
wire     [31:0] n2945;
wire     [31:0] n2946;
wire     [31:0] n2947;
wire     [31:0] n2948;
wire     [31:0] n2949;
wire     [31:0] n2950;
wire     [31:0] n2951;
wire     [31:0] n2952;
wire     [31:0] n2953;
wire     [31:0] n2954;
wire     [31:0] n2955;
wire     [31:0] n2956;
wire     [31:0] n2957;
wire     [31:0] n2958;
wire     [31:0] n2959;
wire     [31:0] n2960;
wire     [31:0] n2961;
wire     [31:0] n2962;
wire     [31:0] n2963;
wire     [31:0] n2964;
wire            n2965;
wire      [4:0] n2966;
wire            n2967;
wire            n2968;
wire            n2969;
wire            n2970;
wire            n2971;
wire            n2972;
wire            n2973;
wire            n2974;
wire            n2975;
wire            n2976;
wire            n2977;
wire            n2978;
wire            n2979;
wire            n2980;
wire            n2981;
wire            n2982;
wire            n2983;
wire            n2984;
wire            n2985;
wire            n2986;
wire            n2987;
wire            n2988;
wire            n2989;
wire            n2990;
wire            n2991;
wire            n2992;
wire            n2993;
wire            n2994;
wire            n2995;
wire            n2996;
wire            n2997;
wire            n2998;
wire     [31:0] n2999;
wire     [31:0] n3000;
wire     [31:0] n3001;
wire     [31:0] n3002;
wire     [31:0] n3003;
wire     [31:0] n3004;
wire     [31:0] n3005;
wire     [31:0] n3006;
wire     [31:0] n3007;
wire     [31:0] n3008;
wire     [31:0] n3009;
wire     [31:0] n3010;
wire     [31:0] n3011;
wire     [31:0] n3012;
wire     [31:0] n3013;
wire     [31:0] n3014;
wire     [31:0] n3015;
wire     [31:0] n3016;
wire     [31:0] n3017;
wire     [31:0] n3018;
wire     [31:0] n3019;
wire     [31:0] n3020;
wire     [31:0] n3021;
wire     [31:0] n3022;
wire     [31:0] n3023;
wire     [31:0] n3024;
wire     [31:0] n3025;
wire     [31:0] n3026;
wire     [31:0] n3027;
wire     [31:0] n3028;
wire     [31:0] n3029;
wire     [31:0] n3030;
wire            n3031;
wire            n3032;
wire     [31:0] n3033;
wire            n3034;
wire     [31:0] n3035;
wire     [31:0] n3036;
wire     [31:0] n3037;
wire     [31:0] n3038;
wire     [31:0] n3039;
wire            n3040;
wire     [31:0] n3041;
wire     [31:0] n3042;
wire     [31:0] n3043;
wire     [31:0] n3044;
wire     [31:0] n3045;
wire     [31:0] n3046;
wire     [31:0] n3047;
wire     [31:0] n3048;
wire     [31:0] n3049;
wire     [31:0] n3050;
wire            n3051;
wire     [31:0] n3052;
wire     [31:0] n3053;
wire     [31:0] n3054;
wire     [31:0] n3055;
wire     [31:0] n3056;
wire     [31:0] n3057;
wire     [31:0] n3058;
wire     [31:0] n3059;
wire     [31:0] n3060;
wire     [31:0] n3061;
wire     [31:0] n3062;
wire     [31:0] n3063;
wire     [31:0] n3064;
wire     [31:0] n3065;
wire     [31:0] n3066;
wire     [31:0] n3067;
wire     [31:0] n3068;
wire            n3069;
wire            n3070;
wire            n3071;
wire            n3072;
wire            n3073;
wire            n3074;
wire            n3075;
wire            n3076;
wire            n3077;
wire            n3078;
wire            n3079;
wire            n3080;
wire            n3081;
wire            n3082;
wire            n3083;
wire            n3084;
wire            n3085;
wire            n3086;
wire            n3087;
wire            n3088;
wire            n3089;
wire            n3090;
wire            n3091;
wire            n3092;
wire            n3093;
wire            n3094;
wire            n3095;
wire            n3096;
wire            n3097;
wire            n3098;
wire            n3099;
wire            n3100;
wire            n3101;
wire            n3102;
wire            n3103;
wire            n3104;
wire            n3105;
wire            n3106;
wire            n3107;
wire            n3108;
wire            n3109;
wire            n3110;
wire            n3111;
wire            n3112;
wire            n3113;
wire            n3114;
wire            n3115;
wire            n3116;
wire            n3117;
wire            n3118;
wire            n3119;
wire            n3120;
wire            n3121;
wire            n3122;
wire            n3123;
wire            n3124;
wire            n3125;
wire            n3126;
wire            n3127;
wire            n3128;
wire            n3129;
wire            n3130;
wire            n3131;
wire            n3132;
wire            n3133;
wire            n3134;
wire            n3135;
wire            n3136;
wire            n3137;
wire            n3138;
wire            n3139;
wire            n3140;
wire            n3141;
wire            n3142;
wire            n3143;
wire            n3144;
wire            n3145;
wire            n3146;
wire            n3147;
wire            n3148;
wire            n3149;
wire            n3150;
wire            n3151;
wire            n3152;
wire            n3153;
wire            n3154;
wire            n3155;
wire            n3156;
wire            n3157;
wire            n3158;
wire            n3159;
wire            n3160;
wire            n3161;
wire            n3162;
wire            n3163;
wire            n3164;
wire            n3165;
wire            n3166;
wire            n3167;
wire            n3168;
wire            n3169;
wire            n3170;
wire            n3171;
wire            n3172;
wire            n3173;
wire            n3174;
wire            n3175;
wire            n3176;
wire            n3177;
wire            n3178;
wire            n3179;
wire            n3180;
wire            n3181;
wire            n3182;
wire            n3183;
wire            n3184;
wire            n3185;
wire            n3186;
wire            n3187;
wire            n3188;
wire            n3189;
wire            n3190;
wire            n3191;
wire            n3192;
wire            n3193;
wire            n3194;
wire            n3195;
wire            n3196;
wire            n3197;
wire            n3198;
wire            n3199;
wire            n3200;
wire            n3201;
wire            n3202;
wire            n3203;
wire            n3204;
wire            n3205;
wire            n3206;
wire            n3207;
wire            n3208;
wire            n3209;
wire            n3210;
wire            n3211;
wire            n3212;
wire            n3213;
wire            n3214;
wire            n3215;
wire            n3216;
wire            n3217;
wire            n3218;
wire            n3219;
wire            n3220;
wire            n3221;
wire            n3222;
wire            n3223;
wire            n3224;
wire            n3225;
wire            n3226;
wire            n3227;
wire            n3228;
wire            n3229;
wire            n3230;
wire            n3231;
wire            n3232;
wire            n3233;
wire            n3234;
wire            n3235;
wire            n3236;
wire            n3237;
wire            n3238;
wire            n3239;
wire            n3240;
wire            n3241;
wire            n3242;
wire            n3243;
wire            n3244;
wire            n3245;
wire            n3246;
wire            n3247;
wire            n3248;
wire            n3249;
wire            n3250;
wire            n3251;
wire            n3252;
wire            n3253;
wire            n3254;
wire            n3255;
wire            n3256;
wire            n3257;
wire            n3258;
wire            n3259;
wire            n3260;
wire            n3261;
wire            n3262;
wire            n3263;
wire            n3264;
wire            n3265;
wire            n3266;
wire            n3267;
wire            n3268;
wire            n3269;
wire            n3270;
wire            n3271;
wire            n3272;
wire            n3273;
wire            n3274;
wire            n3275;
wire            n3276;
wire            n3277;
wire            n3278;
wire            n3279;
wire            n3280;
wire            n3281;
wire            n3282;
wire            n3283;
wire            n3284;
wire            n3285;
wire            n3286;
wire            n3287;
wire            n3288;
wire            n3289;
wire            n3290;
wire            n3291;
wire            n3292;
wire            n3293;
wire            n3294;
wire            n3295;
wire            n3296;
wire            n3297;
wire            n3298;
wire            n3299;
wire            n3300;
wire            n3301;
wire            n3302;
wire            n3303;
wire            n3304;
wire            n3305;
wire            n3306;
wire            n3307;
wire            n3308;
wire            n3309;
wire            n3310;
wire            n3311;
wire            n3312;
wire            n3313;
wire            n3314;
wire            n3315;
wire            n3316;
wire            n3317;
wire            n3318;
wire            n3319;
wire            n3320;
wire            n3321;
wire            n3322;
wire            n3323;
wire            n3324;
wire            n3325;
wire            n3326;
wire            n3327;
wire            n3328;
wire            n3329;
wire            n3330;
wire            n3331;
wire            n3332;
wire            n3333;
wire            n3334;
wire            n3335;
wire            n3336;
wire            n3337;
wire            n3338;
wire            n3339;
wire            n3340;
wire            n3341;
wire            n3342;
wire            n3343;
wire            n3344;
wire            n3345;
wire            n3346;
wire            n3347;
wire            n3348;
wire            n3349;
wire            n3350;
wire            n3351;
wire            n3352;
wire            n3353;
wire            n3354;
wire            n3355;
wire            n3356;
wire            n3357;
wire            n3358;
wire            n3359;
wire            n3360;
wire            n3361;
wire            n3362;
wire            n3363;
wire            n3364;
wire            n3365;
wire            n3366;
wire            n3367;
wire            n3368;
wire            n3369;
wire            n3370;
wire            n3371;
wire            n3372;
wire            n3373;
wire            n3374;
wire            n3375;
wire            n3376;
wire            n3377;
wire            n3378;
wire            n3379;
wire            n3380;
wire            n3381;
wire            n3382;
wire            n3383;
wire            n3384;
wire            n3385;
wire            n3386;
wire            n3387;
wire            n3388;
wire            n3389;
wire            n3390;
wire            n3391;
wire            n3392;
wire            n3393;
wire            n3394;
wire            n3395;
wire            n3396;
wire            n3397;
wire            n3398;
wire            n3399;
wire            n3400;
wire            n3401;
wire            n3402;
wire            n3403;
wire            n3404;
wire            n3405;
wire            n3406;
wire            n3407;
wire            n3408;
wire            n3409;
wire            n3410;
wire            n3411;
wire            n3412;
wire            n3413;
wire            n3414;
wire            n3415;
wire            n3416;
wire            n3417;
wire            n3418;
wire            n3419;
wire            n3420;
wire            n3421;
wire            n3422;
wire            n3423;
wire            n3424;
wire            n3425;
wire            n3426;
wire            n3427;
wire            n3428;
wire            n3429;
wire            n3430;
wire            n3431;
wire            n3432;
wire            n3433;
wire            n3434;
wire            n3435;
wire            n3436;
wire            n3437;
wire            n3438;
wire            n3439;
wire            n3440;
wire            n3441;
wire            n3442;
wire            n3443;
wire            n3444;
wire            n3445;
wire            n3446;
wire            n3447;
wire            n3448;
wire            n3449;
wire            n3450;
wire            n3451;
wire            n3452;
wire            n3453;
wire            n3454;
wire            n3455;
wire            n3456;
wire            n3457;
wire            n3458;
wire            n3459;
wire            n3460;
wire            n3461;
wire            n3462;
wire            n3463;
wire            n3464;
wire            n3465;
wire            n3466;
wire            n3467;
wire            n3468;
wire            n3469;
wire            n3470;
wire            n3471;
wire            n3472;
wire            n3473;
wire            n3474;
wire            n3475;
wire            n3476;
wire            n3477;
wire            n3478;
wire            n3479;
wire            n3480;
wire            n3481;
wire            n3482;
wire            n3483;
wire            n3484;
wire            n3485;
wire            n3486;
wire            n3487;
wire            n3488;
wire            n3489;
wire            n3490;
wire            n3491;
wire            n3492;
wire            n3493;
wire            n3494;
wire            n3495;
wire            n3496;
wire            n3497;
wire            n3498;
wire            n3499;
wire            n3500;
wire            n3501;
wire            n3502;
wire            n3503;
wire            n3504;
wire            n3505;
wire            n3506;
wire            n3507;
wire            n3508;
wire            n3509;
wire            n3510;
wire            n3511;
wire            n3512;
wire            n3513;
wire            n3514;
wire            n3515;
wire            n3516;
wire            n3517;
wire            n3518;
wire            n3519;
wire            n3520;
wire            n3521;
wire            n3522;
wire            n3523;
wire            n3524;
wire            n3525;
wire            n3526;
wire            n3527;
wire            n3528;
wire            n3529;
wire            n3530;
wire            n3531;
wire            n3532;
wire            n3533;
wire            n3534;
wire            n3535;
wire            n3536;
wire            n3537;
wire            n3538;
wire            n3539;
wire            n3540;
wire            n3541;
wire            n3542;
wire            n3543;
wire            n3544;
wire            n3545;
wire            n3546;
wire            n3547;
wire            n3548;
wire            n3549;
wire            n3550;
wire            n3551;
wire            n3552;
wire            n3553;
wire            n3554;
wire            n3555;
wire            n3556;
wire            n3557;
wire            n3558;
wire            n3559;
wire            n3560;
wire            n3561;
wire            n3562;
wire            n3563;
wire            n3564;
wire            n3565;
wire            n3566;
wire            n3567;
wire            n3568;
wire            n3569;
wire            n3570;
wire            n3571;
wire            n3572;
wire            n3573;
wire            n3574;
wire            n3575;
wire            n3576;
wire            n3577;
wire            n3578;
wire            n3579;
wire            n3580;
wire            n3581;
wire            n3582;
wire            n3583;
wire            n3584;
wire            n3585;
wire            n3586;
wire            n3587;
wire            n3588;
wire            n3589;
wire            n3590;
wire            n3591;
wire            n3592;
wire            n3593;
wire            n3594;
wire            n3595;
wire            n3596;
wire     [31:0] n3597;
wire     [31:0] n3598;
wire     [31:0] n3599;
wire     [31:0] n3600;
wire     [31:0] n3601;
wire     [31:0] n3602;
wire     [31:0] n3603;
wire     [31:0] n3604;
wire     [31:0] n3605;
wire     [31:0] n3606;
wire     [31:0] n3607;
wire     [31:0] n3608;
wire     [31:0] n3609;
wire     [31:0] n3610;
wire     [31:0] n3611;
wire     [31:0] n3612;
wire     [31:0] n3613;
wire     [31:0] n3614;
wire     [31:0] n3615;
wire     [31:0] n3616;
wire     [31:0] n3617;
wire     [31:0] n3618;
wire     [31:0] n3619;
wire     [31:0] n3620;
wire     [31:0] n3621;
wire     [31:0] n3622;
wire     [31:0] n3623;
wire     [31:0] n3624;
wire     [31:0] n3625;
wire     [31:0] n3626;
wire     [31:0] n3627;
wire     [31:0] n3628;
wire     [31:0] n3629;
wire     [31:0] n3630;
wire     [31:0] n3631;
wire     [31:0] n3632;
wire     [31:0] n3633;
wire     [31:0] n3634;
wire     [31:0] n3635;
wire     [31:0] n3636;
wire     [31:0] n3637;
wire     [31:0] n3638;
wire     [31:0] n3639;
wire     [31:0] n3640;
wire     [31:0] n3641;
wire     [31:0] n3642;
wire     [31:0] n3643;
wire     [31:0] n3644;
wire     [31:0] n3645;
wire     [31:0] n3646;
wire     [31:0] n3647;
wire     [31:0] n3648;
wire     [31:0] n3649;
wire     [31:0] n3650;
wire     [31:0] n3651;
wire     [31:0] n3652;
wire     [31:0] n3653;
wire     [31:0] n3654;
wire     [31:0] n3655;
wire     [31:0] n3656;
wire     [31:0] n3657;
wire     [31:0] n3658;
wire     [31:0] n3659;
wire     [31:0] n3660;
wire     [31:0] n3661;
wire     [31:0] n3662;
wire     [31:0] n3663;
wire     [31:0] n3664;
wire     [31:0] n3665;
wire     [31:0] n3666;
wire     [31:0] n3667;
wire     [31:0] n3668;
wire     [31:0] n3669;
wire     [31:0] n3670;
wire     [31:0] n3671;
wire     [31:0] n3672;
wire     [31:0] n3673;
wire     [31:0] n3674;
wire     [31:0] n3675;
wire     [31:0] n3676;
wire     [31:0] n3677;
wire     [31:0] n3678;
wire     [31:0] n3679;
wire     [31:0] n3680;
wire     [31:0] n3681;
wire     [31:0] n3682;
wire     [31:0] n3683;
wire     [31:0] n3684;
wire     [31:0] n3685;
wire     [31:0] n3686;
wire     [31:0] n3687;
wire     [31:0] n3688;
wire     [31:0] n3689;
wire     [31:0] n3690;
wire     [31:0] n3691;
wire     [31:0] n3692;
wire     [31:0] n3693;
wire     [31:0] n3694;
wire     [31:0] n3695;
wire     [31:0] n3696;
wire     [31:0] n3697;
wire     [31:0] n3698;
wire     [31:0] n3699;
wire     [31:0] n3700;
wire     [31:0] n3701;
wire     [31:0] n3702;
wire     [31:0] n3703;
wire     [31:0] n3704;
wire     [31:0] n3705;
wire     [31:0] n3706;
wire     [31:0] n3707;
wire     [31:0] n3708;
wire     [31:0] n3709;
wire     [31:0] n3710;
wire     [31:0] n3711;
wire     [31:0] n3712;
wire     [31:0] n3713;
wire     [31:0] n3714;
wire     [31:0] n3715;
wire     [31:0] n3716;
wire     [31:0] n3717;
wire     [31:0] n3718;
wire     [31:0] n3719;
wire     [31:0] n3720;
wire     [31:0] n3721;
wire     [31:0] n3722;
wire     [31:0] n3723;
wire     [31:0] n3724;
wire     [31:0] n3725;
wire     [31:0] n3726;
wire     [31:0] n3727;
wire     [31:0] n3728;
wire     [31:0] n3729;
wire     [31:0] n3730;
wire     [31:0] n3731;
wire     [31:0] n3732;
wire     [31:0] n3733;
wire     [31:0] n3734;
wire     [31:0] n3735;
wire     [31:0] n3736;
wire     [31:0] n3737;
wire     [31:0] n3738;
wire     [31:0] n3739;
wire     [31:0] n3740;
wire     [31:0] n3741;
wire     [31:0] n3742;
wire     [31:0] n3743;
wire     [31:0] n3744;
wire     [31:0] n3745;
wire     [31:0] n3746;
wire     [31:0] n3747;
wire     [31:0] n3748;
wire     [31:0] n3749;
wire     [31:0] n3750;
wire     [31:0] n3751;
wire     [31:0] n3752;
wire     [31:0] n3753;
wire     [31:0] n3754;
wire     [31:0] n3755;
wire     [31:0] n3756;
wire     [31:0] n3757;
wire     [31:0] n3758;
wire     [31:0] n3759;
wire     [31:0] n3760;
wire     [31:0] n3761;
wire     [31:0] n3762;
wire     [31:0] n3763;
wire     [31:0] n3764;
wire     [31:0] n3765;
wire     [31:0] n3766;
wire     [31:0] n3767;
wire     [31:0] n3768;
wire     [31:0] n3769;
wire     [31:0] n3770;
wire     [31:0] n3771;
wire     [31:0] n3772;
wire     [31:0] n3773;
wire     [31:0] n3774;
wire     [31:0] n3775;
wire     [31:0] n3776;
wire     [31:0] n3777;
wire     [31:0] n3778;
wire     [31:0] n3779;
wire     [31:0] n3780;
wire     [31:0] n3781;
wire     [31:0] n3782;
wire     [31:0] n3783;
wire     [31:0] n3784;
wire     [31:0] n3785;
wire     [31:0] n3786;
wire     [31:0] n3787;
wire     [31:0] n3788;
wire     [31:0] n3789;
wire     [31:0] n3790;
wire     [31:0] n3791;
wire     [31:0] n3792;
wire     [31:0] n3793;
wire     [31:0] n3794;
wire     [31:0] n3795;
wire     [31:0] n3796;
wire     [31:0] n3797;
wire     [31:0] n3798;
wire     [31:0] n3799;
wire     [31:0] n3800;
wire     [31:0] n3801;
wire     [31:0] n3802;
wire     [31:0] n3803;
wire     [31:0] n3804;
wire     [31:0] n3805;
wire     [31:0] n3806;
wire     [31:0] n3807;
wire     [31:0] n3808;
wire     [31:0] n3809;
wire     [31:0] n3810;
wire     [31:0] n3811;
wire     [31:0] n3812;
wire     [31:0] n3813;
wire     [31:0] n3814;
wire     [31:0] n3815;
wire     [31:0] n3816;
wire     [31:0] n3817;
wire     [31:0] n3818;
wire     [31:0] n3819;
wire     [31:0] n3820;
wire     [31:0] n3821;
wire     [31:0] n3822;
wire     [31:0] n3823;
wire     [31:0] n3824;
wire     [31:0] n3825;
wire     [31:0] n3826;
wire     [31:0] n3827;
wire     [31:0] n3828;
wire     [31:0] n3829;
wire     [31:0] n3830;
wire     [31:0] n3831;
wire     [31:0] n3832;
wire     [31:0] n3833;
wire     [31:0] n3834;
wire     [31:0] n3835;
wire     [31:0] n3836;
wire     [31:0] n3837;
wire     [31:0] n3838;
wire     [31:0] n3839;
wire     [31:0] n3840;
wire     [31:0] n3841;
wire     [31:0] n3842;
wire     [31:0] n3843;
wire     [31:0] n3844;
wire     [31:0] n3845;
wire     [31:0] n3846;
wire     [31:0] n3847;
wire     [31:0] n3848;
wire     [31:0] n3849;
wire     [31:0] n3850;
wire     [31:0] n3851;
wire     [31:0] n3852;
wire     [31:0] n3853;
wire     [31:0] n3854;
wire     [31:0] n3855;
wire     [31:0] n3856;
wire     [31:0] n3857;
wire     [31:0] n3858;
wire     [31:0] n3859;
wire     [31:0] n3860;
wire     [31:0] n3861;
wire     [31:0] n3862;
wire     [31:0] n3863;
wire     [31:0] n3864;
wire     [31:0] n3865;
wire     [31:0] n3866;
wire     [31:0] n3867;
wire     [31:0] n3868;
wire     [31:0] n3869;
wire     [31:0] n3870;
wire     [31:0] n3871;
wire     [31:0] n3872;
wire     [31:0] n3873;
wire     [31:0] n3874;
wire     [31:0] n3875;
wire     [31:0] n3876;
wire     [31:0] n3877;
wire     [31:0] n3878;
wire     [31:0] n3879;
wire     [31:0] n3880;
wire     [31:0] n3881;
wire     [31:0] n3882;
wire     [31:0] n3883;
wire     [31:0] n3884;
wire     [31:0] n3885;
wire     [31:0] n3886;
wire     [31:0] n3887;
wire     [31:0] n3888;
wire     [31:0] n3889;
wire     [31:0] n3890;
wire     [31:0] n3891;
wire     [31:0] n3892;
wire     [31:0] n3893;
wire     [31:0] n3894;
wire     [31:0] n3895;
wire     [31:0] n3896;
wire     [31:0] n3897;
wire     [31:0] n3898;
wire     [31:0] n3899;
wire     [31:0] n3900;
wire     [31:0] n3901;
wire     [31:0] n3902;
wire     [31:0] n3903;
wire     [31:0] n3904;
wire     [31:0] n3905;
wire     [31:0] n3906;
wire     [31:0] n3907;
wire     [31:0] n3908;
wire     [31:0] n3909;
wire     [31:0] n3910;
wire     [31:0] n3911;
wire     [31:0] n3912;
wire     [31:0] n3913;
wire     [31:0] n3914;
wire     [31:0] n3915;
wire     [31:0] n3916;
wire     [31:0] n3917;
wire     [31:0] n3918;
wire     [31:0] n3919;
wire     [31:0] n3920;
wire     [31:0] n3921;
wire     [31:0] n3922;
wire     [31:0] n3923;
wire     [31:0] n3924;
wire     [31:0] n3925;
wire     [31:0] n3926;
wire     [31:0] n3927;
wire     [31:0] n3928;
wire     [31:0] n3929;
wire     [31:0] n3930;
wire     [31:0] n3931;
wire     [31:0] n3932;
wire     [31:0] n3933;
wire     [31:0] n3934;
wire     [31:0] n3935;
wire     [31:0] n3936;
wire     [31:0] n3937;
wire     [31:0] n3938;
wire     [31:0] n3939;
wire     [31:0] n3940;
wire     [31:0] n3941;
wire     [31:0] n3942;
wire     [31:0] n3943;
wire     [31:0] n3944;
wire     [31:0] n3945;
wire     [31:0] n3946;
wire     [31:0] n3947;
wire     [31:0] n3948;
wire     [31:0] n3949;
wire     [31:0] n3950;
wire     [31:0] n3951;
wire     [31:0] n3952;
wire     [31:0] n3953;
wire     [31:0] n3954;
wire     [31:0] n3955;
wire     [31:0] n3956;
wire     [31:0] n3957;
wire     [31:0] n3958;
wire     [31:0] n3959;
wire     [31:0] n3960;
wire     [31:0] n3961;
wire     [31:0] n3962;
wire     [31:0] n3963;
wire     [31:0] n3964;
wire     [31:0] n3965;
wire     [31:0] n3966;
wire     [31:0] n3967;
wire     [31:0] n3968;
wire     [31:0] n3969;
wire     [31:0] n3970;
wire     [31:0] n3971;
wire     [31:0] n3972;
wire     [31:0] n3973;
wire     [31:0] n3974;
wire     [31:0] n3975;
wire     [31:0] n3976;
wire     [31:0] n3977;
wire     [31:0] n3978;
wire     [31:0] n3979;
wire     [31:0] n3980;
wire     [31:0] n3981;
wire     [31:0] n3982;
wire     [31:0] n3983;
wire     [31:0] n3984;
wire     [31:0] n3985;
wire     [31:0] n3986;
wire     [31:0] n3987;
wire     [31:0] n3988;
wire     [31:0] n3989;
wire     [31:0] n3990;
wire     [31:0] n3991;
wire     [31:0] n3992;
wire     [31:0] n3993;
wire     [31:0] n3994;
wire     [31:0] n3995;
wire     [31:0] n3996;
wire     [31:0] n3997;
wire     [31:0] n3998;
wire     [31:0] n3999;
wire     [31:0] n4000;
wire     [31:0] n4001;
wire     [31:0] n4002;
wire     [31:0] n4003;
wire     [31:0] n4004;
wire     [31:0] n4005;
wire     [31:0] n4006;
wire     [31:0] n4007;
wire     [31:0] n4008;
wire     [31:0] n4009;
wire     [31:0] n4010;
wire     [31:0] n4011;
wire     [31:0] n4012;
wire     [31:0] n4013;
wire     [31:0] n4014;
wire     [31:0] n4015;
wire     [31:0] n4016;
wire     [31:0] n4017;
wire     [31:0] n4018;
wire     [31:0] n4019;
wire     [31:0] n4020;
wire     [31:0] n4021;
wire     [31:0] n4022;
wire     [31:0] n4023;
wire     [31:0] n4024;
wire     [31:0] n4025;
wire     [31:0] n4026;
wire     [31:0] n4027;
wire     [31:0] n4028;
wire     [31:0] n4029;
wire     [31:0] n4030;
wire     [31:0] n4031;
wire     [31:0] n4032;
wire     [31:0] n4033;
wire     [31:0] n4034;
wire     [31:0] n4035;
wire     [31:0] n4036;
wire     [31:0] n4037;
wire     [31:0] n4038;
wire     [31:0] n4039;
wire     [31:0] n4040;
wire     [31:0] n4041;
wire     [31:0] n4042;
wire     [31:0] n4043;
wire     [31:0] n4044;
wire     [31:0] n4045;
wire     [31:0] n4046;
wire     [31:0] n4047;
wire     [31:0] n4048;
wire     [31:0] n4049;
wire     [31:0] n4050;
wire     [31:0] n4051;
wire     [31:0] n4052;
wire     [31:0] n4053;
wire     [31:0] n4054;
wire     [31:0] n4055;
wire     [31:0] n4056;
wire     [31:0] n4057;
wire     [31:0] n4058;
wire     [31:0] n4059;
wire     [31:0] n4060;
wire     [31:0] n4061;
wire     [31:0] n4062;
wire     [31:0] n4063;
wire     [31:0] n4064;
wire     [31:0] n4065;
wire     [31:0] n4066;
wire     [31:0] n4067;
wire     [31:0] n4068;
wire     [31:0] n4069;
wire     [31:0] n4070;
wire     [31:0] n4071;
wire     [31:0] n4072;
wire     [31:0] n4073;
wire     [31:0] n4074;
wire     [31:0] n4075;
wire     [31:0] n4076;
wire     [31:0] n4077;
wire     [31:0] n4078;
wire     [31:0] n4079;
wire     [31:0] n4080;
wire     [31:0] n4081;
wire     [31:0] n4082;
wire     [31:0] n4083;
wire     [31:0] n4084;
wire     [31:0] n4085;
wire     [31:0] n4086;
wire     [31:0] n4087;
wire     [31:0] n4088;
wire     [31:0] n4089;
wire     [31:0] n4090;
wire     [31:0] n4091;
wire     [31:0] n4092;
wire     [31:0] n4093;
wire     [31:0] n4094;
wire     [31:0] n4095;
wire     [31:0] n4096;
wire     [31:0] n4097;
wire     [31:0] n4098;
wire     [31:0] n4099;
wire     [31:0] n4100;
wire     [31:0] n4101;
wire     [31:0] n4102;
wire     [31:0] n4103;
wire     [31:0] n4104;
wire     [31:0] n4105;
wire     [31:0] n4106;
wire     [31:0] n4107;
wire     [31:0] n4108;
wire     [31:0] n4109;
wire     [31:0] n4110;
wire     [31:0] n4111;
wire     [31:0] n4112;
wire     [31:0] n4113;
wire     [31:0] n4114;
wire     [31:0] n4115;
wire     [31:0] n4116;
wire     [31:0] n4117;
wire     [31:0] n4118;
wire            n4119;
wire            n4120;
wire            n4121;
wire            n4122;
wire            n4123;
wire            n4124;
wire            n4125;
wire            n4126;
wire            n4127;
wire            n4128;
wire            n4129;
wire            n4130;
wire            n4131;
wire            n4132;
wire            n4133;
wire            n4134;
wire            n4135;
wire            n4136;
wire            n4137;
wire            n4138;
wire            n4139;
wire            n4140;
wire            n4141;
wire            n4142;
wire            n4143;
wire            n4144;
wire            n4145;
wire            n4146;
wire            n4147;
wire            n4148;
wire            n4149;
wire            n4150;
wire            n4151;
wire            n4152;
wire            n4153;
wire            n4154;
wire            n4155;
wire            n4156;
wire            n4157;
wire            n4158;
wire            n4159;
wire            n4160;
wire            n4161;
wire            n4162;
wire            n4163;
wire            n4164;
wire            n4165;
wire            n4166;
wire            n4167;
wire            n4168;
wire            n4169;
wire            n4170;
wire            n4171;
wire            n4172;
wire            n4173;
wire            n4174;
wire            n4175;
wire            n4176;
wire            n4177;
wire            n4178;
wire            n4179;
wire            n4180;
wire            n4181;
wire            n4182;
wire            n4183;
wire            n4184;
wire            n4185;
wire            n4186;
wire            n4187;
wire            n4188;
wire            n4189;
wire            n4190;
wire            n4191;
wire            n4192;
wire            n4193;
wire            n4194;
wire            n4195;
wire            n4196;
wire            n4197;
wire            n4198;
wire            n4199;
wire            n4200;
wire            n4201;
wire            n4202;
wire            n4203;
wire            n4204;
wire            n4205;
wire            n4206;
wire            n4207;
wire            n4208;
wire            n4209;
wire            n4210;
wire            n4211;
wire            n4212;
wire            n4213;
wire            n4214;
wire            n4215;
wire            n4216;
wire            n4217;
wire            n4218;
wire            n4219;
wire            n4220;
wire            n4221;
wire            n4222;
wire            n4223;
wire            n4224;
wire            n4225;
wire            n4226;
wire            n4227;
wire            n4228;
wire            n4229;
wire            n4230;
wire            n4231;
wire            n4232;
wire            n4233;
wire            n4234;
wire            n4235;
wire            n4236;
wire            n4237;
wire            n4238;
wire            n4239;
wire            n4240;
wire            n4241;
wire            n4242;
wire            n4243;
wire            n4244;
wire            n4245;
wire            n4246;
wire            n4247;
wire            n4248;
wire            n4249;
wire            n4250;
wire            n4251;
wire            n4252;
wire            n4253;
wire            n4254;
wire            n4255;
wire            n4256;
wire            n4257;
wire            n4258;
wire            n4259;
wire            n4260;
wire            n4261;
wire            n4262;
wire            n4263;
wire            n4264;
wire            n4265;
wire            n4266;
wire            n4267;
wire            n4268;
wire            n4269;
wire            n4270;
wire            n4271;
wire            n4272;
wire            n4273;
wire            n4274;
wire            n4275;
wire            n4276;
wire            n4277;
wire            n4278;
wire            n4279;
wire            n4280;
wire            n4281;
wire            n4282;
wire            n4283;
wire            n4284;
wire            n4285;
wire            n4286;
wire            n4287;
wire            n4288;
wire            n4289;
wire            n4290;
wire            n4291;
wire            n4292;
wire            n4293;
wire            n4294;
wire            n4295;
wire            n4296;
wire            n4297;
wire            n4298;
wire            n4299;
wire            n4300;
wire            n4301;
wire            n4302;
wire            n4303;
wire            n4304;
wire            n4305;
wire            n4306;
wire            n4307;
wire            n4308;
wire            n4309;
wire            n4310;
wire            n4311;
wire            n4312;
wire            n4313;
wire            n4314;
wire            n4315;
wire            n4316;
wire            n4317;
wire            n4318;
wire            n4319;
wire            n4320;
wire            n4321;
wire            n4322;
wire            n4323;
wire            n4324;
wire            n4325;
wire            n4326;
wire            n4327;
wire            n4328;
wire            n4329;
wire            n4330;
wire            n4331;
wire            n4332;
wire            n4333;
wire            n4334;
wire            n4335;
wire            n4336;
wire            n4337;
wire            n4338;
wire            n4339;
wire            n4340;
wire            n4341;
wire            n4342;
wire            n4343;
wire            n4344;
wire            n4345;
wire            n4346;
wire            n4347;
wire            n4348;
wire            n4349;
wire            n4350;
wire            n4351;
wire            n4352;
wire            n4353;
wire            n4354;
wire            n4355;
wire            n4356;
wire            n4357;
wire            n4358;
wire            n4359;
wire            n4360;
wire            n4361;
wire            n4362;
wire            n4363;
wire            n4364;
wire            n4365;
wire            n4366;
wire            n4367;
wire            n4368;
wire            n4369;
wire            n4370;
wire            n4371;
wire            n4372;
wire            n4373;
wire            n4374;
wire            n4375;
wire            n4376;
wire            n4377;
wire            n4378;
wire            n4379;
wire            n4380;
wire            n4381;
wire            n4382;
wire            n4383;
wire            n4384;
wire            n4385;
wire            n4386;
wire            n4387;
wire            n4388;
wire            n4389;
wire            n4390;
wire            n4391;
wire            n4392;
wire            n4393;
wire            n4394;
wire            n4395;
wire            n4396;
wire            n4397;
wire            n4398;
wire            n4399;
wire            n4400;
wire            n4401;
wire            n4402;
wire            n4403;
wire            n4404;
wire            n4405;
wire            n4406;
wire            n4407;
wire            n4408;
wire            n4409;
wire            n4410;
wire            n4411;
wire            n4412;
wire            n4413;
wire            n4414;
wire            n4415;
wire            n4416;
wire            n4417;
wire            n4418;
wire            n4419;
wire            n4420;
wire            n4421;
wire            n4422;
wire            n4423;
wire            n4424;
wire            n4425;
wire            n4426;
wire            n4427;
wire            n4428;
wire            n4429;
wire            n4430;
wire            n4431;
wire            n4432;
wire            n4433;
wire            n4434;
wire            n4435;
wire            n4436;
wire            n4437;
wire            n4438;
wire            n4439;
wire            n4440;
wire            n4441;
wire            n4442;
wire            n4443;
wire            n4444;
wire            n4445;
wire            n4446;
wire            n4447;
wire            n4448;
wire            n4449;
wire            n4450;
wire            n4451;
wire            n4452;
wire            n4453;
wire            n4454;
wire            n4455;
wire            n4456;
wire            n4457;
wire            n4458;
wire            n4459;
wire            n4460;
wire            n4461;
wire            n4462;
wire            n4463;
wire            n4464;
wire            n4465;
wire            n4466;
wire            n4467;
wire            n4468;
wire            n4469;
wire            n4470;
wire            n4471;
wire            n4472;
wire            n4473;
wire            n4474;
wire            n4475;
wire            n4476;
wire            n4477;
wire            n4478;
wire            n4479;
wire            n4480;
wire            n4481;
wire            n4482;
wire            n4483;
wire            n4484;
wire            n4485;
wire            n4486;
wire            n4487;
wire            n4488;
wire            n4489;
wire            n4490;
wire            n4491;
wire            n4492;
wire            n4493;
wire            n4494;
wire            n4495;
wire            n4496;
wire            n4497;
wire            n4498;
wire            n4499;
wire            n4500;
wire            n4501;
wire            n4502;
wire            n4503;
wire            n4504;
wire            n4505;
wire            n4506;
wire            n4507;
wire            n4508;
wire            n4509;
wire            n4510;
wire            n4511;
wire            n4512;
wire            n4513;
wire            n4514;
wire            n4515;
wire            n4516;
wire            n4517;
wire            n4518;
wire            n4519;
wire            n4520;
wire            n4521;
wire            n4522;
wire            n4523;
wire            n4524;
wire            n4525;
wire            n4526;
wire            n4527;
wire            n4528;
wire            n4529;
wire            n4530;
wire            n4531;
wire            n4532;
wire            n4533;
wire            n4534;
wire            n4535;
wire            n4536;
wire            n4537;
wire            n4538;
wire            n4539;
wire            n4540;
wire            n4541;
wire            n4542;
wire            n4543;
wire            n4544;
wire            n4545;
wire            n4546;
wire            n4547;
wire            n4548;
wire            n4549;
wire            n4550;
wire            n4551;
wire            n4552;
wire            n4553;
wire            n4554;
wire            n4555;
wire            n4556;
wire            n4557;
wire            n4558;
wire            n4559;
wire            n4560;
wire            n4561;
wire            n4562;
wire            n4563;
wire            n4564;
wire            n4565;
wire            n4566;
wire            n4567;
wire            n4568;
wire            n4569;
wire            n4570;
wire            n4571;
wire            n4572;
wire            n4573;
wire            n4574;
wire            n4575;
wire            n4576;
wire            n4577;
wire            n4578;
wire            n4579;
wire            n4580;
wire            n4581;
wire            n4582;
wire            n4583;
wire            n4584;
wire            n4585;
wire            n4586;
wire            n4587;
wire            n4588;
wire            n4589;
wire            n4590;
wire            n4591;
wire            n4592;
wire            n4593;
wire            n4594;
wire            n4595;
wire            n4596;
wire            n4597;
wire            n4598;
wire            n4599;
wire            n4600;
wire            n4601;
wire            n4602;
wire            n4603;
wire            n4604;
wire            n4605;
wire            n4606;
wire            n4607;
wire            n4608;
wire            n4609;
wire            n4610;
wire            n4611;
wire            n4612;
wire            n4613;
wire            n4614;
wire            n4615;
wire            n4616;
wire            n4617;
wire            n4618;
wire            n4619;
wire            n4620;
wire            n4621;
wire            n4622;
wire            n4623;
wire            n4624;
wire            n4625;
wire            n4626;
wire            n4627;
wire            n4628;
wire            n4629;
wire            n4630;
wire     [31:0] n4631;
wire     [31:0] n4632;
wire     [31:0] n4633;
wire     [31:0] n4634;
wire     [31:0] n4635;
wire     [31:0] n4636;
wire     [31:0] n4637;
wire     [31:0] n4638;
wire     [31:0] n4639;
wire     [31:0] n4640;
wire     [31:0] n4641;
wire     [31:0] n4642;
wire     [31:0] n4643;
wire     [31:0] n4644;
wire     [31:0] n4645;
wire     [31:0] n4646;
wire     [31:0] n4647;
wire     [31:0] n4648;
wire     [31:0] n4649;
wire     [31:0] n4650;
wire     [31:0] n4651;
wire     [31:0] n4652;
wire     [31:0] n4653;
wire     [31:0] n4654;
wire     [31:0] n4655;
wire     [31:0] n4656;
wire     [31:0] n4657;
wire     [31:0] n4658;
wire     [31:0] n4659;
wire     [31:0] n4660;
wire     [31:0] n4661;
wire     [31:0] n4662;
wire     [31:0] n4663;
wire     [31:0] n4664;
wire     [31:0] n4665;
wire     [31:0] n4666;
wire     [31:0] n4667;
wire     [31:0] n4668;
wire     [31:0] n4669;
wire     [31:0] n4670;
wire     [31:0] n4671;
wire     [31:0] n4672;
wire     [31:0] n4673;
wire     [31:0] n4674;
wire     [31:0] n4675;
wire     [31:0] n4676;
wire     [31:0] n4677;
wire     [31:0] n4678;
wire     [31:0] n4679;
wire     [31:0] n4680;
wire     [31:0] n4681;
wire     [31:0] n4682;
wire     [31:0] n4683;
wire     [31:0] n4684;
wire     [31:0] n4685;
wire     [31:0] n4686;
wire     [31:0] n4687;
wire     [31:0] n4688;
wire     [31:0] n4689;
wire     [31:0] n4690;
wire     [31:0] n4691;
wire     [31:0] n4692;
wire     [31:0] n4693;
wire     [31:0] n4694;
wire     [31:0] n4695;
wire     [31:0] n4696;
wire     [31:0] n4697;
wire     [31:0] n4698;
wire     [31:0] n4699;
wire     [31:0] n4700;
wire     [31:0] n4701;
wire     [31:0] n4702;
wire     [31:0] n4703;
wire     [31:0] n4704;
wire     [31:0] n4705;
wire     [31:0] n4706;
wire     [31:0] n4707;
wire     [31:0] n4708;
wire     [31:0] n4709;
wire     [31:0] n4710;
wire     [31:0] n4711;
wire     [31:0] n4712;
wire     [31:0] n4713;
wire     [31:0] n4714;
wire     [31:0] n4715;
wire     [31:0] n4716;
wire     [31:0] n4717;
wire     [31:0] n4718;
wire     [31:0] n4719;
wire     [31:0] n4720;
wire     [31:0] n4721;
wire     [31:0] n4722;
wire     [31:0] n4723;
wire     [31:0] n4724;
wire     [31:0] n4725;
wire     [31:0] n4726;
wire     [31:0] n4727;
wire     [31:0] n4728;
wire     [31:0] n4729;
wire     [31:0] n4730;
wire     [31:0] n4731;
wire     [31:0] n4732;
wire     [31:0] n4733;
wire     [31:0] n4734;
wire     [31:0] n4735;
wire     [31:0] n4736;
wire     [31:0] n4737;
wire     [31:0] n4738;
wire     [31:0] n4739;
wire     [31:0] n4740;
wire     [31:0] n4741;
wire     [31:0] n4742;
wire     [31:0] n4743;
wire     [31:0] n4744;
wire     [31:0] n4745;
wire     [31:0] n4746;
wire     [31:0] n4747;
wire     [31:0] n4748;
wire     [31:0] n4749;
wire     [31:0] n4750;
wire     [31:0] n4751;
wire     [31:0] n4752;
wire     [31:0] n4753;
wire     [31:0] n4754;
wire     [31:0] n4755;
wire     [31:0] n4756;
wire     [31:0] n4757;
wire     [31:0] n4758;
wire     [31:0] n4759;
wire     [31:0] n4760;
wire     [31:0] n4761;
wire     [31:0] n4762;
wire     [31:0] n4763;
wire     [31:0] n4764;
wire     [31:0] n4765;
wire     [31:0] n4766;
wire     [31:0] n4767;
wire     [31:0] n4768;
wire     [31:0] n4769;
wire     [31:0] n4770;
wire     [31:0] n4771;
wire     [31:0] n4772;
wire     [31:0] n4773;
wire     [31:0] n4774;
wire     [31:0] n4775;
wire     [31:0] n4776;
wire     [31:0] n4777;
wire     [31:0] n4778;
wire     [31:0] n4779;
wire     [31:0] n4780;
wire     [31:0] n4781;
wire     [31:0] n4782;
wire     [31:0] n4783;
wire     [31:0] n4784;
wire     [31:0] n4785;
wire     [31:0] n4786;
wire     [31:0] n4787;
wire     [31:0] n4788;
wire     [31:0] n4789;
wire     [31:0] n4790;
wire     [31:0] n4791;
wire     [31:0] n4792;
wire     [31:0] n4793;
wire     [31:0] n4794;
wire     [31:0] n4795;
wire     [31:0] n4796;
wire     [31:0] n4797;
wire     [31:0] n4798;
wire     [31:0] n4799;
wire     [31:0] n4800;
wire     [31:0] n4801;
wire     [31:0] n4802;
wire     [31:0] n4803;
wire     [31:0] n4804;
wire     [31:0] n4805;
wire     [31:0] n4806;
wire     [31:0] n4807;
wire     [31:0] n4808;
wire     [31:0] n4809;
wire     [31:0] n4810;
wire     [31:0] n4811;
wire     [31:0] n4812;
wire     [31:0] n4813;
wire     [31:0] n4814;
wire     [31:0] n4815;
wire     [31:0] n4816;
wire     [31:0] n4817;
wire     [31:0] n4818;
wire     [31:0] n4819;
wire     [31:0] n4820;
wire     [31:0] n4821;
wire     [31:0] n4822;
wire     [31:0] n4823;
wire     [31:0] n4824;
wire     [31:0] n4825;
wire     [31:0] n4826;
wire     [31:0] n4827;
wire     [31:0] n4828;
wire     [31:0] n4829;
wire     [31:0] n4830;
wire     [31:0] n4831;
wire     [31:0] n4832;
wire     [31:0] n4833;
wire     [31:0] n4834;
wire     [31:0] n4835;
wire     [31:0] n4836;
wire     [31:0] n4837;
wire     [31:0] n4838;
wire     [31:0] n4839;
wire     [31:0] n4840;
wire     [31:0] n4841;
wire     [31:0] n4842;
wire     [31:0] n4843;
wire     [31:0] n4844;
wire     [31:0] n4845;
wire     [31:0] n4846;
wire     [31:0] n4847;
wire     [31:0] n4848;
wire     [31:0] n4849;
wire     [31:0] n4850;
wire     [31:0] n4851;
wire     [31:0] n4852;
wire     [31:0] n4853;
wire     [31:0] n4854;
wire     [31:0] n4855;
wire     [31:0] n4856;
wire     [31:0] n4857;
wire     [31:0] n4858;
wire     [31:0] n4859;
wire     [31:0] n4860;
wire     [31:0] n4861;
wire     [31:0] n4862;
wire     [31:0] n4863;
wire     [31:0] n4864;
wire     [31:0] n4865;
wire     [31:0] n4866;
wire     [31:0] n4867;
wire     [31:0] n4868;
wire     [31:0] n4869;
wire     [31:0] n4870;
wire     [31:0] n4871;
wire     [31:0] n4872;
wire     [31:0] n4873;
wire     [31:0] n4874;
wire     [31:0] n4875;
wire     [31:0] n4876;
wire     [31:0] n4877;
wire     [31:0] n4878;
wire     [31:0] n4879;
wire     [31:0] n4880;
wire     [31:0] n4881;
wire     [31:0] n4882;
wire     [31:0] n4883;
wire     [31:0] n4884;
wire     [31:0] n4885;
wire     [31:0] n4886;
wire     [31:0] n4887;
wire     [31:0] n4888;
wire     [31:0] n4889;
wire     [31:0] n4890;
wire     [31:0] n4891;
wire     [31:0] n4892;
wire     [31:0] n4893;
wire     [31:0] n4894;
wire     [31:0] n4895;
wire     [31:0] n4896;
wire     [31:0] n4897;
wire     [31:0] n4898;
wire     [31:0] n4899;
wire     [31:0] n4900;
wire     [31:0] n4901;
wire     [31:0] n4902;
wire     [31:0] n4903;
wire     [31:0] n4904;
wire     [31:0] n4905;
wire     [31:0] n4906;
wire     [31:0] n4907;
wire     [31:0] n4908;
wire     [31:0] n4909;
wire     [31:0] n4910;
wire     [31:0] n4911;
wire     [31:0] n4912;
wire     [31:0] n4913;
wire     [31:0] n4914;
wire     [31:0] n4915;
wire     [31:0] n4916;
wire     [31:0] n4917;
wire     [31:0] n4918;
wire     [31:0] n4919;
wire     [31:0] n4920;
wire     [31:0] n4921;
wire     [31:0] n4922;
wire     [31:0] n4923;
wire     [31:0] n4924;
wire     [31:0] n4925;
wire     [31:0] n4926;
wire     [31:0] n4927;
wire     [31:0] n4928;
wire     [31:0] n4929;
wire     [31:0] n4930;
wire     [31:0] n4931;
wire     [31:0] n4932;
wire     [31:0] n4933;
wire     [31:0] n4934;
wire     [31:0] n4935;
wire     [31:0] n4936;
wire     [31:0] n4937;
wire     [31:0] n4938;
wire     [31:0] n4939;
wire     [31:0] n4940;
wire     [31:0] n4941;
wire     [31:0] n4942;
wire     [31:0] n4943;
wire     [31:0] n4944;
wire     [31:0] n4945;
wire     [31:0] n4946;
wire     [31:0] n4947;
wire     [31:0] n4948;
wire     [31:0] n4949;
wire     [31:0] n4950;
wire     [31:0] n4951;
wire     [31:0] n4952;
wire     [31:0] n4953;
wire     [31:0] n4954;
wire     [31:0] n4955;
wire     [31:0] n4956;
wire     [31:0] n4957;
wire     [31:0] n4958;
wire     [31:0] n4959;
wire     [31:0] n4960;
wire     [31:0] n4961;
wire     [31:0] n4962;
wire     [31:0] n4963;
wire     [31:0] n4964;
wire     [31:0] n4965;
wire     [31:0] n4966;
wire     [31:0] n4967;
wire     [31:0] n4968;
wire     [31:0] n4969;
wire     [31:0] n4970;
wire     [31:0] n4971;
wire     [31:0] n4972;
wire     [31:0] n4973;
wire     [31:0] n4974;
wire     [31:0] n4975;
wire     [31:0] n4976;
wire     [31:0] n4977;
wire     [31:0] n4978;
wire     [31:0] n4979;
wire     [31:0] n4980;
wire     [31:0] n4981;
wire     [31:0] n4982;
wire     [31:0] n4983;
wire     [31:0] n4984;
wire     [31:0] n4985;
wire     [31:0] n4986;
wire     [31:0] n4987;
wire     [31:0] n4988;
wire     [31:0] n4989;
wire     [31:0] n4990;
wire     [31:0] n4991;
wire     [31:0] n4992;
wire     [31:0] n4993;
wire     [31:0] n4994;
wire     [31:0] n4995;
wire     [31:0] n4996;
wire     [31:0] n4997;
wire     [31:0] n4998;
wire     [31:0] n4999;
wire     [31:0] n5000;
wire     [31:0] n5001;
wire     [31:0] n5002;
wire     [31:0] n5003;
wire     [31:0] n5004;
wire     [31:0] n5005;
wire     [31:0] n5006;
wire     [31:0] n5007;
wire     [31:0] n5008;
wire     [31:0] n5009;
wire     [31:0] n5010;
wire     [31:0] n5011;
wire     [31:0] n5012;
wire     [31:0] n5013;
wire     [31:0] n5014;
wire     [31:0] n5015;
wire     [31:0] n5016;
wire     [31:0] n5017;
wire     [31:0] n5018;
wire     [31:0] n5019;
wire     [31:0] n5020;
wire     [31:0] n5021;
wire     [31:0] n5022;
wire     [31:0] n5023;
wire     [31:0] n5024;
wire     [31:0] n5025;
wire     [31:0] n5026;
wire     [31:0] n5027;
wire     [31:0] n5028;
wire     [31:0] n5029;
wire     [31:0] n5030;
wire     [31:0] n5031;
wire     [31:0] n5032;
wire     [31:0] n5033;
wire     [31:0] n5034;
wire     [31:0] n5035;
wire     [31:0] n5036;
wire     [31:0] n5037;
wire     [31:0] n5038;
wire     [31:0] n5039;
wire     [31:0] n5040;
wire     [31:0] n5041;
wire     [31:0] n5042;
wire     [31:0] n5043;
wire     [31:0] n5044;
wire     [31:0] n5045;
wire     [31:0] n5046;
wire     [31:0] n5047;
wire     [31:0] n5048;
wire     [31:0] n5049;
wire     [31:0] n5050;
wire     [31:0] n5051;
wire     [31:0] n5052;
wire     [31:0] n5053;
wire     [31:0] n5054;
wire     [31:0] n5055;
wire     [31:0] n5056;
wire     [31:0] n5057;
wire     [31:0] n5058;
wire     [31:0] n5059;
wire     [31:0] n5060;
wire     [31:0] n5061;
wire     [31:0] n5062;
wire     [31:0] n5063;
wire     [31:0] n5064;
wire     [31:0] n5065;
wire     [31:0] n5066;
wire     [31:0] n5067;
wire     [31:0] n5068;
wire     [31:0] n5069;
wire     [31:0] n5070;
wire     [31:0] n5071;
wire     [31:0] n5072;
wire     [31:0] n5073;
wire     [31:0] n5074;
wire     [31:0] n5075;
wire     [31:0] n5076;
wire     [31:0] n5077;
wire     [31:0] n5078;
wire     [31:0] n5079;
wire     [31:0] n5080;
wire     [31:0] n5081;
wire     [31:0] n5082;
wire     [31:0] n5083;
wire     [31:0] n5084;
wire     [31:0] n5085;
wire     [31:0] n5086;
wire     [31:0] n5087;
wire     [31:0] n5088;
wire     [31:0] n5089;
wire     [31:0] n5090;
wire     [31:0] n5091;
wire     [31:0] n5092;
wire     [31:0] n5093;
wire     [31:0] n5094;
wire     [31:0] n5095;
wire     [31:0] n5096;
wire     [31:0] n5097;
wire     [31:0] n5098;
wire     [31:0] n5099;
wire     [31:0] n5100;
wire     [31:0] n5101;
wire     [31:0] n5102;
wire     [31:0] n5103;
wire     [31:0] n5104;
wire     [31:0] n5105;
wire     [31:0] n5106;
wire     [31:0] n5107;
wire     [31:0] n5108;
wire     [31:0] n5109;
wire     [31:0] n5110;
wire     [31:0] n5111;
wire     [31:0] n5112;
wire     [31:0] n5113;
wire     [31:0] n5114;
wire     [31:0] n5115;
wire     [31:0] n5116;
wire     [31:0] n5117;
wire     [31:0] n5118;
wire     [31:0] n5119;
wire     [31:0] n5120;
wire     [31:0] n5121;
wire     [31:0] n5122;
wire     [31:0] n5123;
wire     [31:0] n5124;
wire     [31:0] n5125;
wire     [31:0] n5126;
wire     [31:0] n5127;
wire     [31:0] n5128;
wire     [31:0] n5129;
wire     [31:0] n5130;
wire     [31:0] n5131;
wire     [31:0] n5132;
wire     [31:0] n5133;
wire     [31:0] n5134;
wire     [31:0] n5135;
wire     [31:0] n5136;
wire     [31:0] n5137;
wire     [31:0] n5138;
wire     [31:0] n5139;
wire     [31:0] n5140;
wire     [31:0] n5141;
wire     [31:0] n5142;
wire     [31:0] n5143;
wire     [31:0] n5144;
wire     [31:0] n5145;
wire     [31:0] n5146;
wire     [31:0] n5147;
wire     [31:0] n5148;
wire     [31:0] n5149;
wire     [31:0] n5150;
wire     [31:0] n5151;
wire     [31:0] n5152;
wire            n5153;
wire            n5154;
wire     [31:0] n5155;
wire     [31:0] n5156;
wire     [31:0] n5157;
wire     [31:0] n5158;
wire     [31:0] n5159;
wire     [31:0] n5160;
wire     [31:0] n5161;
wire     [31:0] n5162;
wire     [31:0] n5163;
wire     [31:0] n5164;
wire     [31:0] n5165;
wire     [31:0] n5166;
wire     [31:0] n5167;
wire     [31:0] n5168;
wire     [31:0] n5169;
wire     [31:0] n5170;
wire     [31:0] n5171;
wire     [31:0] n5172;
wire     [31:0] n5173;
wire     [31:0] n5174;
wire     [31:0] n5175;
wire     [31:0] n5176;
wire     [31:0] n5177;
wire     [31:0] n5178;
wire     [31:0] n5179;
wire     [31:0] n5180;
wire     [31:0] n5181;
wire     [31:0] n5182;
wire     [31:0] n5183;
wire     [31:0] n5184;
wire     [31:0] n5185;
wire     [31:0] n5186;
wire     [31:0] n5187;
wire            n5188;
wire            n5189;
wire            n5190;
wire            n5191;
wire            n5192;
wire            n5193;
wire            n5194;
wire            n5195;
wire            n5196;
wire            n5197;
wire            n5198;
wire            n5199;
wire            n5200;
wire            n5201;
wire            n5202;
wire            n5203;
wire            n5204;
wire            n5205;
wire            n5206;
wire            n5207;
wire            n5208;
wire            n5209;
wire            n5210;
wire            n5211;
wire            n5212;
wire            n5213;
wire            n5214;
wire            n5215;
wire            n5216;
wire            n5217;
wire            n5218;
wire            n5219;
wire            n5220;
wire            n5221;
wire            n5222;
wire            n5223;
wire            n5224;
wire            n5225;
wire            n5226;
wire            n5227;
wire            n5228;
wire            n5229;
wire            n5230;
wire            n5231;
wire            n5232;
wire            n5233;
wire            n5234;
wire            n5235;
wire            n5236;
wire            n5237;
wire            n5238;
wire            n5239;
wire            n5240;
wire            n5241;
wire            n5242;
wire            n5243;
wire            n5244;
wire            n5245;
wire            n5246;
wire            n5247;
wire            n5248;
wire            n5249;
wire            n5250;
wire            n5251;
wire            n5252;
wire            n5253;
wire            n5254;
wire            n5255;
wire            n5256;
wire            n5257;
wire            n5258;
wire            n5259;
wire            n5260;
wire            n5261;
wire            n5262;
wire            n5263;
wire            n5264;
wire            n5265;
wire            n5266;
wire            n5267;
wire            n5268;
wire            n5269;
wire            n5270;
wire            n5271;
wire            n5272;
wire            n5273;
wire            n5274;
wire            n5275;
wire            n5276;
wire            n5277;
wire            n5278;
wire            n5279;
wire            n5280;
wire            n5281;
wire            n5282;
wire            n5283;
wire            n5284;
wire            n5285;
wire            n5286;
wire            n5287;
wire            n5288;
wire            n5289;
wire            n5290;
wire            n5291;
wire            n5292;
wire            n5293;
wire            n5294;
wire            n5295;
wire            n5296;
wire            n5297;
wire            n5298;
wire            n5299;
wire            n5300;
wire            n5301;
wire            n5302;
wire            n5303;
wire            n5304;
wire            n5305;
wire            n5306;
wire            n5307;
wire            n5308;
wire            n5309;
wire            n5310;
wire            n5311;
wire            n5312;
wire            n5313;
wire            n5314;
wire            n5315;
wire            n5316;
wire            n5317;
wire            n5318;
wire            n5319;
wire            n5320;
wire            n5321;
wire            n5322;
wire            n5323;
wire            n5324;
wire            n5325;
wire            n5326;
wire            n5327;
wire            n5328;
wire            n5329;
wire            n5330;
wire            n5331;
wire            n5332;
wire            n5333;
wire            n5334;
wire            n5335;
wire            n5336;
wire            n5337;
wire            n5338;
wire            n5339;
wire            n5340;
wire            n5341;
wire            n5342;
wire            n5343;
wire            n5344;
wire            n5345;
wire            n5346;
wire            n5347;
wire            n5348;
wire            n5349;
wire            n5350;
wire            n5351;
wire            n5352;
wire            n5353;
wire            n5354;
wire            n5355;
wire            n5356;
wire            n5357;
wire            n5358;
wire            n5359;
wire            n5360;
wire            n5361;
wire            n5362;
wire            n5363;
wire            n5364;
wire            n5365;
wire            n5366;
wire            n5367;
wire            n5368;
wire            n5369;
wire            n5370;
wire            n5371;
wire            n5372;
wire            n5373;
wire            n5374;
wire            n5375;
wire            n5376;
wire            n5377;
wire            n5378;
wire            n5379;
wire            n5380;
wire            n5381;
wire            n5382;
wire            n5383;
wire            n5384;
wire            n5385;
wire            n5386;
wire            n5387;
wire            n5388;
wire            n5389;
wire            n5390;
wire            n5391;
wire            n5392;
wire            n5393;
wire            n5394;
wire            n5395;
wire            n5396;
wire            n5397;
wire            n5398;
wire            n5399;
wire            n5400;
wire            n5401;
wire            n5402;
wire            n5403;
wire            n5404;
wire            n5405;
wire            n5406;
wire            n5407;
wire            n5408;
wire            n5409;
wire            n5410;
wire            n5411;
wire            n5412;
wire            n5413;
wire            n5414;
wire            n5415;
wire            n5416;
wire            n5417;
wire            n5418;
wire            n5419;
wire            n5420;
wire            n5421;
wire            n5422;
wire            n5423;
wire            n5424;
wire            n5425;
wire            n5426;
wire            n5427;
wire            n5428;
wire            n5429;
wire            n5430;
wire            n5431;
wire            n5432;
wire            n5433;
wire            n5434;
wire            n5435;
wire            n5436;
wire            n5437;
wire            n5438;
wire            n5439;
wire            n5440;
wire            n5441;
wire            n5442;
wire            n5443;
wire            n5444;
wire            n5445;
wire            n5446;
wire            n5447;
wire            n5448;
wire            n5449;
wire            n5450;
wire            n5451;
wire            n5452;
wire            n5453;
wire            n5454;
wire            n5455;
wire            n5456;
wire            n5457;
wire            n5458;
wire            n5459;
wire            n5460;
wire            n5461;
wire            n5462;
wire            n5463;
wire            n5464;
wire            n5465;
wire            n5466;
wire            n5467;
wire            n5468;
wire            n5469;
wire            n5470;
wire            n5471;
wire            n5472;
wire            n5473;
wire            n5474;
wire            n5475;
wire            n5476;
wire            n5477;
wire            n5478;
wire            n5479;
wire            n5480;
wire            n5481;
wire            n5482;
wire            n5483;
wire            n5484;
wire            n5485;
wire            n5486;
wire            n5487;
wire            n5488;
wire            n5489;
wire            n5490;
wire            n5491;
wire            n5492;
wire            n5493;
wire            n5494;
wire            n5495;
wire            n5496;
wire            n5497;
wire            n5498;
wire            n5499;
wire            n5500;
wire            n5501;
wire            n5502;
wire            n5503;
wire            n5504;
wire            n5505;
wire            n5506;
wire            n5507;
wire            n5508;
wire            n5509;
wire            n5510;
wire            n5511;
wire            n5512;
wire            n5513;
wire            n5514;
wire            n5515;
wire            n5516;
wire            n5517;
wire            n5518;
wire            n5519;
wire            n5520;
wire            n5521;
wire            n5522;
wire            n5523;
wire            n5524;
wire            n5525;
wire            n5526;
wire            n5527;
wire            n5528;
wire            n5529;
wire            n5530;
wire            n5531;
wire            n5532;
wire            n5533;
wire            n5534;
wire            n5535;
wire            n5536;
wire            n5537;
wire            n5538;
wire            n5539;
wire            n5540;
wire            n5541;
wire            n5542;
wire            n5543;
wire            n5544;
wire            n5545;
wire            n5546;
wire            n5547;
wire            n5548;
wire            n5549;
wire            n5550;
wire            n5551;
wire            n5552;
wire            n5553;
wire            n5554;
wire            n5555;
wire            n5556;
wire            n5557;
wire            n5558;
wire            n5559;
wire            n5560;
wire            n5561;
wire            n5562;
wire            n5563;
wire            n5564;
wire            n5565;
wire            n5566;
wire            n5567;
wire            n5568;
wire            n5569;
wire            n5570;
wire            n5571;
wire            n5572;
wire            n5573;
wire            n5574;
wire            n5575;
wire            n5576;
wire            n5577;
wire            n5578;
wire            n5579;
wire            n5580;
wire            n5581;
wire            n5582;
wire            n5583;
wire            n5584;
wire            n5585;
wire            n5586;
wire            n5587;
wire            n5588;
wire            n5589;
wire            n5590;
wire            n5591;
wire            n5592;
wire            n5593;
wire            n5594;
wire            n5595;
wire            n5596;
wire            n5597;
wire            n5598;
wire            n5599;
wire            n5600;
wire            n5601;
wire            n5602;
wire            n5603;
wire            n5604;
wire            n5605;
wire            n5606;
wire            n5607;
wire            n5608;
wire            n5609;
wire            n5610;
wire            n5611;
wire            n5612;
wire            n5613;
wire            n5614;
wire            n5615;
wire            n5616;
wire            n5617;
wire            n5618;
wire            n5619;
wire            n5620;
wire            n5621;
wire            n5622;
wire            n5623;
wire            n5624;
wire            n5625;
wire            n5626;
wire            n5627;
wire            n5628;
wire            n5629;
wire            n5630;
wire            n5631;
wire            n5632;
wire            n5633;
wire            n5634;
wire            n5635;
wire            n5636;
wire            n5637;
wire            n5638;
wire            n5639;
wire            n5640;
wire            n5641;
wire            n5642;
wire            n5643;
wire            n5644;
wire            n5645;
wire            n5646;
wire            n5647;
wire            n5648;
wire            n5649;
wire            n5650;
wire            n5651;
wire            n5652;
wire            n5653;
wire            n5654;
wire            n5655;
wire            n5656;
wire            n5657;
wire            n5658;
wire            n5659;
wire            n5660;
wire            n5661;
wire            n5662;
wire            n5663;
wire            n5664;
wire            n5665;
wire            n5666;
wire            n5667;
wire            n5668;
wire            n5669;
wire            n5670;
wire            n5671;
wire            n5672;
wire            n5673;
wire            n5674;
wire            n5675;
wire            n5676;
wire            n5677;
wire            n5678;
wire            n5679;
wire            n5680;
wire            n5681;
wire            n5682;
wire            n5683;
wire            n5684;
wire            n5685;
wire            n5686;
wire            n5687;
wire            n5688;
wire            n5689;
wire            n5690;
wire            n5691;
wire            n5692;
wire            n5693;
wire            n5694;
wire            n5695;
wire            n5696;
wire            n5697;
wire            n5698;
wire            n5699;
wire            n5700;
wire            n5701;
wire            n5702;
wire            n5703;
wire            n5704;
wire            n5705;
wire            n5706;
wire            n5707;
wire            n5708;
wire            n5709;
wire            n5710;
wire            n5711;
wire            n5712;
wire            n5713;
wire            n5714;
wire            n5715;
wire     [31:0] n5716;
wire     [31:0] n5717;
wire     [31:0] n5718;
wire     [31:0] n5719;
wire     [31:0] n5720;
wire     [31:0] n5721;
wire     [31:0] n5722;
wire     [31:0] n5723;
wire     [31:0] n5724;
wire     [31:0] n5725;
wire     [31:0] n5726;
wire     [31:0] n5727;
wire     [31:0] n5728;
wire     [31:0] n5729;
wire     [31:0] n5730;
wire     [31:0] n5731;
wire     [31:0] n5732;
wire     [31:0] n5733;
wire     [31:0] n5734;
wire     [31:0] n5735;
wire     [31:0] n5736;
wire     [31:0] n5737;
wire     [31:0] n5738;
wire     [31:0] n5739;
wire     [31:0] n5740;
wire     [31:0] n5741;
wire     [31:0] n5742;
wire     [31:0] n5743;
wire     [31:0] n5744;
wire     [31:0] n5745;
wire     [31:0] n5746;
wire     [31:0] n5747;
wire     [31:0] n5748;
wire     [31:0] n5749;
wire     [31:0] n5750;
wire     [31:0] n5751;
wire     [31:0] n5752;
wire     [31:0] n5753;
wire     [31:0] n5754;
wire     [31:0] n5755;
wire     [31:0] n5756;
wire     [31:0] n5757;
wire     [31:0] n5758;
wire     [31:0] n5759;
wire     [31:0] n5760;
wire     [31:0] n5761;
wire     [31:0] n5762;
wire     [31:0] n5763;
wire     [31:0] n5764;
wire     [31:0] n5765;
wire     [31:0] n5766;
wire     [31:0] n5767;
wire     [31:0] n5768;
wire     [31:0] n5769;
wire     [31:0] n5770;
wire     [31:0] n5771;
wire     [31:0] n5772;
wire     [31:0] n5773;
wire     [31:0] n5774;
wire     [31:0] n5775;
wire     [31:0] n5776;
wire     [31:0] n5777;
wire     [31:0] n5778;
wire     [31:0] n5779;
wire     [31:0] n5780;
wire     [31:0] n5781;
wire     [31:0] n5782;
wire     [31:0] n5783;
wire     [31:0] n5784;
wire     [31:0] n5785;
wire     [31:0] n5786;
wire     [31:0] n5787;
wire     [31:0] n5788;
wire     [31:0] n5789;
wire     [31:0] n5790;
wire     [31:0] n5791;
wire     [31:0] n5792;
wire     [31:0] n5793;
wire     [31:0] n5794;
wire     [31:0] n5795;
wire     [31:0] n5796;
wire     [31:0] n5797;
wire     [31:0] n5798;
wire     [31:0] n5799;
wire     [31:0] n5800;
wire     [31:0] n5801;
wire     [31:0] n5802;
wire     [31:0] n5803;
wire     [31:0] n5804;
wire     [31:0] n5805;
wire     [31:0] n5806;
wire     [31:0] n5807;
wire     [31:0] n5808;
wire     [31:0] n5809;
wire     [31:0] n5810;
wire     [31:0] n5811;
wire     [31:0] n5812;
wire     [31:0] n5813;
wire     [31:0] n5814;
wire     [31:0] n5815;
wire     [31:0] n5816;
wire     [31:0] n5817;
wire     [31:0] n5818;
wire     [31:0] n5819;
wire     [31:0] n5820;
wire     [31:0] n5821;
wire     [31:0] n5822;
wire     [31:0] n5823;
wire     [31:0] n5824;
wire     [31:0] n5825;
wire     [31:0] n5826;
wire     [31:0] n5827;
wire     [31:0] n5828;
wire     [31:0] n5829;
wire     [31:0] n5830;
wire     [31:0] n5831;
wire     [31:0] n5832;
wire     [31:0] n5833;
wire     [31:0] n5834;
wire     [31:0] n5835;
wire     [31:0] n5836;
wire     [31:0] n5837;
wire     [31:0] n5838;
wire     [31:0] n5839;
wire     [31:0] n5840;
wire     [31:0] n5841;
wire     [31:0] n5842;
wire     [31:0] n5843;
wire     [31:0] n5844;
wire     [31:0] n5845;
wire     [31:0] n5846;
wire     [31:0] n5847;
wire     [31:0] n5848;
wire     [31:0] n5849;
wire     [31:0] n5850;
wire     [31:0] n5851;
wire     [31:0] n5852;
wire     [31:0] n5853;
wire     [31:0] n5854;
wire     [31:0] n5855;
wire     [31:0] n5856;
wire     [31:0] n5857;
wire     [31:0] n5858;
wire     [31:0] n5859;
wire     [31:0] n5860;
wire     [31:0] n5861;
wire     [31:0] n5862;
wire     [31:0] n5863;
wire     [31:0] n5864;
wire     [31:0] n5865;
wire     [31:0] n5866;
wire     [31:0] n5867;
wire     [31:0] n5868;
wire     [31:0] n5869;
wire     [31:0] n5870;
wire     [31:0] n5871;
wire     [31:0] n5872;
wire     [31:0] n5873;
wire     [31:0] n5874;
wire     [31:0] n5875;
wire     [31:0] n5876;
wire     [31:0] n5877;
wire     [31:0] n5878;
wire     [31:0] n5879;
wire     [31:0] n5880;
wire     [31:0] n5881;
wire     [31:0] n5882;
wire     [31:0] n5883;
wire     [31:0] n5884;
wire     [31:0] n5885;
wire     [31:0] n5886;
wire     [31:0] n5887;
wire     [31:0] n5888;
wire     [31:0] n5889;
wire     [31:0] n5890;
wire     [31:0] n5891;
wire     [31:0] n5892;
wire     [31:0] n5893;
wire     [31:0] n5894;
wire     [31:0] n5895;
wire     [31:0] n5896;
wire     [31:0] n5897;
wire     [31:0] n5898;
wire     [31:0] n5899;
wire     [31:0] n5900;
wire     [31:0] n5901;
wire     [31:0] n5902;
wire     [31:0] n5903;
wire     [31:0] n5904;
wire     [31:0] n5905;
wire     [31:0] n5906;
wire     [31:0] n5907;
wire     [31:0] n5908;
wire     [31:0] n5909;
wire     [31:0] n5910;
wire     [31:0] n5911;
wire     [31:0] n5912;
wire     [31:0] n5913;
wire     [31:0] n5914;
wire     [31:0] n5915;
wire     [31:0] n5916;
wire     [31:0] n5917;
wire     [31:0] n5918;
wire     [31:0] n5919;
wire     [31:0] n5920;
wire     [31:0] n5921;
wire     [31:0] n5922;
wire     [31:0] n5923;
wire     [31:0] n5924;
wire     [31:0] n5925;
wire     [31:0] n5926;
wire     [31:0] n5927;
wire     [31:0] n5928;
wire     [31:0] n5929;
wire     [31:0] n5930;
wire     [31:0] n5931;
wire     [31:0] n5932;
wire     [31:0] n5933;
wire     [31:0] n5934;
wire     [31:0] n5935;
wire     [31:0] n5936;
wire     [31:0] n5937;
wire     [31:0] n5938;
wire     [31:0] n5939;
wire     [31:0] n5940;
wire     [31:0] n5941;
wire     [31:0] n5942;
wire     [31:0] n5943;
wire     [31:0] n5944;
wire     [31:0] n5945;
wire     [31:0] n5946;
wire     [31:0] n5947;
wire     [31:0] n5948;
wire     [31:0] n5949;
wire     [31:0] n5950;
wire     [31:0] n5951;
wire     [31:0] n5952;
wire     [31:0] n5953;
wire     [31:0] n5954;
wire     [31:0] n5955;
wire     [31:0] n5956;
wire     [31:0] n5957;
wire     [31:0] n5958;
wire     [31:0] n5959;
wire     [31:0] n5960;
wire     [31:0] n5961;
wire     [31:0] n5962;
wire     [31:0] n5963;
wire     [31:0] n5964;
wire     [31:0] n5965;
wire     [31:0] n5966;
wire     [31:0] n5967;
wire     [31:0] n5968;
wire     [31:0] n5969;
wire     [31:0] n5970;
wire     [31:0] n5971;
wire     [31:0] n5972;
wire     [31:0] n5973;
wire     [31:0] n5974;
wire     [31:0] n5975;
wire     [31:0] n5976;
wire     [31:0] n5977;
wire     [31:0] n5978;
wire     [31:0] n5979;
wire     [31:0] n5980;
wire     [31:0] n5981;
wire     [31:0] n5982;
wire     [31:0] n5983;
wire     [31:0] n5984;
wire     [31:0] n5985;
wire     [31:0] n5986;
wire     [31:0] n5987;
wire     [31:0] n5988;
wire     [31:0] n5989;
wire     [31:0] n5990;
wire     [31:0] n5991;
wire     [31:0] n5992;
wire     [31:0] n5993;
wire     [31:0] n5994;
wire     [31:0] n5995;
wire     [31:0] n5996;
wire     [31:0] n5997;
wire     [31:0] n5998;
wire     [31:0] n5999;
wire     [31:0] n6000;
wire     [31:0] n6001;
wire     [31:0] n6002;
wire     [31:0] n6003;
wire     [31:0] n6004;
wire     [31:0] n6005;
wire     [31:0] n6006;
wire     [31:0] n6007;
wire     [31:0] n6008;
wire     [31:0] n6009;
wire     [31:0] n6010;
wire     [31:0] n6011;
wire     [31:0] n6012;
wire     [31:0] n6013;
wire     [31:0] n6014;
wire     [31:0] n6015;
wire     [31:0] n6016;
wire     [31:0] n6017;
wire     [31:0] n6018;
wire     [31:0] n6019;
wire     [31:0] n6020;
wire     [31:0] n6021;
wire     [31:0] n6022;
wire     [31:0] n6023;
wire     [31:0] n6024;
wire     [31:0] n6025;
wire     [31:0] n6026;
wire     [31:0] n6027;
wire     [31:0] n6028;
wire     [31:0] n6029;
wire     [31:0] n6030;
wire     [31:0] n6031;
wire     [31:0] n6032;
wire     [31:0] n6033;
wire     [31:0] n6034;
wire     [31:0] n6035;
wire     [31:0] n6036;
wire     [31:0] n6037;
wire     [31:0] n6038;
wire     [31:0] n6039;
wire     [31:0] n6040;
wire     [31:0] n6041;
wire     [31:0] n6042;
wire     [31:0] n6043;
wire     [31:0] n6044;
wire     [31:0] n6045;
wire     [31:0] n6046;
wire     [31:0] n6047;
wire     [31:0] n6048;
wire     [31:0] n6049;
wire     [31:0] n6050;
wire     [31:0] n6051;
wire     [31:0] n6052;
wire     [31:0] n6053;
wire     [31:0] n6054;
wire     [31:0] n6055;
wire     [31:0] n6056;
wire     [31:0] n6057;
wire     [31:0] n6058;
wire     [31:0] n6059;
wire     [31:0] n6060;
wire     [31:0] n6061;
wire     [31:0] n6062;
wire     [31:0] n6063;
wire     [31:0] n6064;
wire     [31:0] n6065;
wire     [31:0] n6066;
wire     [31:0] n6067;
wire     [31:0] n6068;
wire     [31:0] n6069;
wire     [31:0] n6070;
wire     [31:0] n6071;
wire     [31:0] n6072;
wire     [31:0] n6073;
wire     [31:0] n6074;
wire     [31:0] n6075;
wire     [31:0] n6076;
wire     [31:0] n6077;
wire     [31:0] n6078;
wire     [31:0] n6079;
wire     [31:0] n6080;
wire     [31:0] n6081;
wire     [31:0] n6082;
wire     [31:0] n6083;
wire     [31:0] n6084;
wire     [31:0] n6085;
wire     [31:0] n6086;
wire     [31:0] n6087;
wire     [31:0] n6088;
wire     [31:0] n6089;
wire     [31:0] n6090;
wire     [31:0] n6091;
wire     [31:0] n6092;
wire     [31:0] n6093;
wire     [31:0] n6094;
wire     [31:0] n6095;
wire     [31:0] n6096;
wire     [31:0] n6097;
wire     [31:0] n6098;
wire     [31:0] n6099;
wire     [31:0] n6100;
wire     [31:0] n6101;
wire     [31:0] n6102;
wire     [31:0] n6103;
wire     [31:0] n6104;
wire     [31:0] n6105;
wire     [31:0] n6106;
wire     [31:0] n6107;
wire     [31:0] n6108;
wire     [31:0] n6109;
wire     [31:0] n6110;
wire     [31:0] n6111;
wire     [31:0] n6112;
wire     [31:0] n6113;
wire     [31:0] n6114;
wire     [31:0] n6115;
wire     [31:0] n6116;
wire     [31:0] n6117;
wire     [31:0] n6118;
wire     [31:0] n6119;
wire     [31:0] n6120;
wire     [31:0] n6121;
wire     [31:0] n6122;
wire     [31:0] n6123;
wire     [31:0] n6124;
wire     [31:0] n6125;
wire     [31:0] n6126;
wire     [31:0] n6127;
wire     [31:0] n6128;
wire     [31:0] n6129;
wire     [31:0] n6130;
wire     [31:0] n6131;
wire     [31:0] n6132;
wire     [31:0] n6133;
wire     [31:0] n6134;
wire     [31:0] n6135;
wire     [31:0] n6136;
wire     [31:0] n6137;
wire     [31:0] n6138;
wire     [31:0] n6139;
wire     [31:0] n6140;
wire     [31:0] n6141;
wire     [31:0] n6142;
wire     [31:0] n6143;
wire     [31:0] n6144;
wire     [31:0] n6145;
wire     [31:0] n6146;
wire     [31:0] n6147;
wire     [31:0] n6148;
wire     [31:0] n6149;
wire     [31:0] n6150;
wire     [31:0] n6151;
wire     [31:0] n6152;
wire     [31:0] n6153;
wire     [31:0] n6154;
wire     [31:0] n6155;
wire     [31:0] n6156;
wire     [31:0] n6157;
wire     [31:0] n6158;
wire     [31:0] n6159;
wire     [31:0] n6160;
wire     [31:0] n6161;
wire     [31:0] n6162;
wire     [31:0] n6163;
wire     [31:0] n6164;
wire     [31:0] n6165;
wire     [31:0] n6166;
wire     [31:0] n6167;
wire     [31:0] n6168;
wire     [31:0] n6169;
wire     [31:0] n6170;
wire     [31:0] n6171;
wire     [31:0] n6172;
wire     [31:0] n6173;
wire     [31:0] n6174;
wire     [31:0] n6175;
wire     [31:0] n6176;
wire     [31:0] n6177;
wire     [31:0] n6178;
wire     [31:0] n6179;
wire     [31:0] n6180;
wire     [31:0] n6181;
wire     [31:0] n6182;
wire     [31:0] n6183;
wire     [31:0] n6184;
wire     [31:0] n6185;
wire     [31:0] n6186;
wire     [31:0] n6187;
wire     [31:0] n6188;
wire     [31:0] n6189;
wire     [31:0] n6190;
wire     [31:0] n6191;
wire     [31:0] n6192;
wire     [31:0] n6193;
wire     [31:0] n6194;
wire     [31:0] n6195;
wire     [31:0] n6196;
wire     [31:0] n6197;
wire     [31:0] n6198;
wire     [31:0] n6199;
wire     [31:0] n6200;
wire     [31:0] n6201;
wire     [31:0] n6202;
wire     [31:0] n6203;
wire     [31:0] n6204;
wire     [31:0] n6205;
wire     [31:0] n6206;
wire     [31:0] n6207;
wire     [31:0] n6208;
wire     [31:0] n6209;
wire     [31:0] n6210;
wire     [31:0] n6211;
wire     [31:0] n6212;
wire     [31:0] n6213;
wire     [31:0] n6214;
wire     [31:0] n6215;
wire     [31:0] n6216;
wire     [31:0] n6217;
wire     [31:0] n6218;
wire     [31:0] n6219;
wire     [31:0] n6220;
wire     [31:0] n6221;
wire     [31:0] n6222;
wire     [31:0] n6223;
wire     [31:0] n6224;
wire     [31:0] n6225;
wire     [31:0] n6226;
wire     [31:0] n6227;
wire     [31:0] n6228;
wire     [31:0] n6229;
wire     [31:0] n6230;
wire     [31:0] n6231;
wire     [31:0] n6232;
wire     [31:0] n6233;
wire     [31:0] n6234;
wire     [31:0] n6235;
wire     [31:0] n6236;
wire     [31:0] n6237;
wire            n6238;
wire            n6239;
wire            n6240;
wire            n6241;
wire            n6242;
wire            n6243;
wire            n6244;
wire            n6245;
wire            n6246;
wire            n6247;
wire            n6248;
wire            n6249;
wire            n6250;
wire            n6251;
wire            n6252;
wire            n6253;
wire            n6254;
wire            n6255;
wire            n6256;
wire            n6257;
wire            n6258;
wire            n6259;
wire            n6260;
wire            n6261;
wire            n6262;
wire            n6263;
wire            n6264;
wire            n6265;
wire            n6266;
wire            n6267;
wire            n6268;
wire            n6269;
wire            n6270;
wire            n6271;
wire            n6272;
wire            n6273;
wire            n6274;
wire            n6275;
wire            n6276;
wire            n6277;
wire            n6278;
wire            n6279;
wire            n6280;
wire            n6281;
wire            n6282;
wire            n6283;
wire            n6284;
wire            n6285;
wire            n6286;
wire            n6287;
wire            n6288;
wire            n6289;
wire            n6290;
wire            n6291;
wire            n6292;
wire            n6293;
wire            n6294;
wire            n6295;
wire            n6296;
wire            n6297;
wire            n6298;
wire            n6299;
wire            n6300;
wire            n6301;
wire            n6302;
wire            n6303;
wire            n6304;
wire            n6305;
wire            n6306;
wire            n6307;
wire            n6308;
wire            n6309;
wire            n6310;
wire            n6311;
wire            n6312;
wire            n6313;
wire            n6314;
wire            n6315;
wire            n6316;
wire            n6317;
wire            n6318;
wire            n6319;
wire            n6320;
wire            n6321;
wire            n6322;
wire            n6323;
wire            n6324;
wire            n6325;
wire            n6326;
wire            n6327;
wire            n6328;
wire            n6329;
wire            n6330;
wire            n6331;
wire            n6332;
wire            n6333;
wire            n6334;
wire            n6335;
wire            n6336;
wire            n6337;
wire            n6338;
wire            n6339;
wire            n6340;
wire            n6341;
wire            n6342;
wire            n6343;
wire            n6344;
wire            n6345;
wire            n6346;
wire            n6347;
wire            n6348;
wire            n6349;
wire            n6350;
wire            n6351;
wire            n6352;
wire            n6353;
wire            n6354;
wire            n6355;
wire            n6356;
wire            n6357;
wire            n6358;
wire            n6359;
wire            n6360;
wire            n6361;
wire            n6362;
wire            n6363;
wire            n6364;
wire            n6365;
wire            n6366;
wire            n6367;
wire            n6368;
wire            n6369;
wire            n6370;
wire            n6371;
wire            n6372;
wire            n6373;
wire            n6374;
wire            n6375;
wire            n6376;
wire            n6377;
wire            n6378;
wire            n6379;
wire            n6380;
wire            n6381;
wire            n6382;
wire            n6383;
wire            n6384;
wire            n6385;
wire            n6386;
wire            n6387;
wire            n6388;
wire            n6389;
wire            n6390;
wire            n6391;
wire            n6392;
wire            n6393;
wire            n6394;
wire            n6395;
wire            n6396;
wire            n6397;
wire            n6398;
wire            n6399;
wire            n6400;
wire            n6401;
wire            n6402;
wire            n6403;
wire            n6404;
wire            n6405;
wire            n6406;
wire            n6407;
wire            n6408;
wire            n6409;
wire            n6410;
wire            n6411;
wire            n6412;
wire            n6413;
wire            n6414;
wire            n6415;
wire            n6416;
wire            n6417;
wire            n6418;
wire            n6419;
wire            n6420;
wire            n6421;
wire            n6422;
wire            n6423;
wire            n6424;
wire            n6425;
wire            n6426;
wire            n6427;
wire            n6428;
wire            n6429;
wire            n6430;
wire            n6431;
wire            n6432;
wire            n6433;
wire            n6434;
wire            n6435;
wire            n6436;
wire            n6437;
wire            n6438;
wire            n6439;
wire            n6440;
wire            n6441;
wire            n6442;
wire            n6443;
wire            n6444;
wire            n6445;
wire            n6446;
wire            n6447;
wire            n6448;
wire            n6449;
wire            n6450;
wire            n6451;
wire            n6452;
wire            n6453;
wire            n6454;
wire            n6455;
wire            n6456;
wire            n6457;
wire            n6458;
wire            n6459;
wire            n6460;
wire            n6461;
wire            n6462;
wire            n6463;
wire            n6464;
wire            n6465;
wire            n6466;
wire            n6467;
wire            n6468;
wire            n6469;
wire            n6470;
wire            n6471;
wire            n6472;
wire            n6473;
wire            n6474;
wire            n6475;
wire            n6476;
wire            n6477;
wire            n6478;
wire            n6479;
wire            n6480;
wire            n6481;
wire            n6482;
wire            n6483;
wire            n6484;
wire            n6485;
wire            n6486;
wire            n6487;
wire            n6488;
wire            n6489;
wire            n6490;
wire            n6491;
wire            n6492;
wire            n6493;
wire            n6494;
wire            n6495;
wire            n6496;
wire            n6497;
wire            n6498;
wire            n6499;
wire            n6500;
wire            n6501;
wire            n6502;
wire            n6503;
wire            n6504;
wire            n6505;
wire            n6506;
wire            n6507;
wire            n6508;
wire            n6509;
wire            n6510;
wire            n6511;
wire            n6512;
wire            n6513;
wire            n6514;
wire            n6515;
wire            n6516;
wire            n6517;
wire            n6518;
wire            n6519;
wire            n6520;
wire            n6521;
wire            n6522;
wire            n6523;
wire            n6524;
wire            n6525;
wire            n6526;
wire            n6527;
wire            n6528;
wire            n6529;
wire            n6530;
wire            n6531;
wire            n6532;
wire            n6533;
wire            n6534;
wire            n6535;
wire            n6536;
wire            n6537;
wire            n6538;
wire            n6539;
wire            n6540;
wire            n6541;
wire            n6542;
wire            n6543;
wire            n6544;
wire            n6545;
wire            n6546;
wire            n6547;
wire            n6548;
wire            n6549;
wire            n6550;
wire            n6551;
wire            n6552;
wire            n6553;
wire            n6554;
wire            n6555;
wire            n6556;
wire            n6557;
wire            n6558;
wire            n6559;
wire            n6560;
wire            n6561;
wire            n6562;
wire            n6563;
wire            n6564;
wire            n6565;
wire            n6566;
wire            n6567;
wire            n6568;
wire            n6569;
wire            n6570;
wire            n6571;
wire            n6572;
wire            n6573;
wire            n6574;
wire            n6575;
wire            n6576;
wire            n6577;
wire            n6578;
wire            n6579;
wire            n6580;
wire            n6581;
wire            n6582;
wire            n6583;
wire            n6584;
wire            n6585;
wire            n6586;
wire            n6587;
wire            n6588;
wire            n6589;
wire            n6590;
wire            n6591;
wire            n6592;
wire            n6593;
wire            n6594;
wire            n6595;
wire            n6596;
wire            n6597;
wire            n6598;
wire            n6599;
wire            n6600;
wire            n6601;
wire            n6602;
wire            n6603;
wire            n6604;
wire            n6605;
wire            n6606;
wire            n6607;
wire            n6608;
wire            n6609;
wire            n6610;
wire            n6611;
wire            n6612;
wire            n6613;
wire            n6614;
wire            n6615;
wire            n6616;
wire            n6617;
wire            n6618;
wire            n6619;
wire            n6620;
wire            n6621;
wire            n6622;
wire            n6623;
wire            n6624;
wire            n6625;
wire            n6626;
wire            n6627;
wire            n6628;
wire            n6629;
wire            n6630;
wire            n6631;
wire            n6632;
wire            n6633;
wire            n6634;
wire            n6635;
wire            n6636;
wire            n6637;
wire            n6638;
wire            n6639;
wire            n6640;
wire            n6641;
wire            n6642;
wire            n6643;
wire            n6644;
wire            n6645;
wire            n6646;
wire            n6647;
wire            n6648;
wire            n6649;
wire            n6650;
wire            n6651;
wire            n6652;
wire            n6653;
wire            n6654;
wire            n6655;
wire            n6656;
wire            n6657;
wire            n6658;
wire            n6659;
wire            n6660;
wire            n6661;
wire            n6662;
wire            n6663;
wire            n6664;
wire            n6665;
wire            n6666;
wire            n6667;
wire            n6668;
wire            n6669;
wire            n6670;
wire            n6671;
wire            n6672;
wire            n6673;
wire            n6674;
wire            n6675;
wire            n6676;
wire            n6677;
wire            n6678;
wire            n6679;
wire            n6680;
wire            n6681;
wire            n6682;
wire            n6683;
wire            n6684;
wire            n6685;
wire            n6686;
wire            n6687;
wire            n6688;
wire            n6689;
wire            n6690;
wire            n6691;
wire            n6692;
wire            n6693;
wire            n6694;
wire            n6695;
wire            n6696;
wire            n6697;
wire            n6698;
wire            n6699;
wire            n6700;
wire            n6701;
wire            n6702;
wire            n6703;
wire            n6704;
wire            n6705;
wire            n6706;
wire            n6707;
wire            n6708;
wire            n6709;
wire            n6710;
wire            n6711;
wire            n6712;
wire            n6713;
wire            n6714;
wire            n6715;
wire            n6716;
wire            n6717;
wire            n6718;
wire            n6719;
wire            n6720;
wire            n6721;
wire            n6722;
wire            n6723;
wire            n6724;
wire            n6725;
wire            n6726;
wire            n6727;
wire            n6728;
wire            n6729;
wire            n6730;
wire            n6731;
wire            n6732;
wire            n6733;
wire            n6734;
wire            n6735;
wire            n6736;
wire            n6737;
wire            n6738;
wire            n6739;
wire            n6740;
wire            n6741;
wire            n6742;
wire            n6743;
wire            n6744;
wire            n6745;
wire            n6746;
wire            n6747;
wire            n6748;
wire            n6749;
wire     [31:0] n6750;
wire     [31:0] n6751;
wire     [31:0] n6752;
wire     [31:0] n6753;
wire     [31:0] n6754;
wire     [31:0] n6755;
wire     [31:0] n6756;
wire     [31:0] n6757;
wire     [31:0] n6758;
wire     [31:0] n6759;
wire     [31:0] n6760;
wire     [31:0] n6761;
wire     [31:0] n6762;
wire     [31:0] n6763;
wire     [31:0] n6764;
wire     [31:0] n6765;
wire     [31:0] n6766;
wire     [31:0] n6767;
wire     [31:0] n6768;
wire     [31:0] n6769;
wire     [31:0] n6770;
wire     [31:0] n6771;
wire     [31:0] n6772;
wire     [31:0] n6773;
wire     [31:0] n6774;
wire     [31:0] n6775;
wire     [31:0] n6776;
wire     [31:0] n6777;
wire     [31:0] n6778;
wire     [31:0] n6779;
wire     [31:0] n6780;
wire     [31:0] n6781;
wire     [31:0] n6782;
wire     [31:0] n6783;
wire     [31:0] n6784;
wire     [31:0] n6785;
wire     [31:0] n6786;
wire     [31:0] n6787;
wire     [31:0] n6788;
wire     [31:0] n6789;
wire     [31:0] n6790;
wire     [31:0] n6791;
wire     [31:0] n6792;
wire     [31:0] n6793;
wire     [31:0] n6794;
wire     [31:0] n6795;
wire     [31:0] n6796;
wire     [31:0] n6797;
wire     [31:0] n6798;
wire     [31:0] n6799;
wire     [31:0] n6800;
wire     [31:0] n6801;
wire     [31:0] n6802;
wire     [31:0] n6803;
wire     [31:0] n6804;
wire     [31:0] n6805;
wire     [31:0] n6806;
wire     [31:0] n6807;
wire     [31:0] n6808;
wire     [31:0] n6809;
wire     [31:0] n6810;
wire     [31:0] n6811;
wire     [31:0] n6812;
wire     [31:0] n6813;
wire     [31:0] n6814;
wire     [31:0] n6815;
wire     [31:0] n6816;
wire     [31:0] n6817;
wire     [31:0] n6818;
wire     [31:0] n6819;
wire     [31:0] n6820;
wire     [31:0] n6821;
wire     [31:0] n6822;
wire     [31:0] n6823;
wire     [31:0] n6824;
wire     [31:0] n6825;
wire     [31:0] n6826;
wire     [31:0] n6827;
wire     [31:0] n6828;
wire     [31:0] n6829;
wire     [31:0] n6830;
wire     [31:0] n6831;
wire     [31:0] n6832;
wire     [31:0] n6833;
wire     [31:0] n6834;
wire     [31:0] n6835;
wire     [31:0] n6836;
wire     [31:0] n6837;
wire     [31:0] n6838;
wire     [31:0] n6839;
wire     [31:0] n6840;
wire     [31:0] n6841;
wire     [31:0] n6842;
wire     [31:0] n6843;
wire     [31:0] n6844;
wire     [31:0] n6845;
wire     [31:0] n6846;
wire     [31:0] n6847;
wire     [31:0] n6848;
wire     [31:0] n6849;
wire     [31:0] n6850;
wire     [31:0] n6851;
wire     [31:0] n6852;
wire     [31:0] n6853;
wire     [31:0] n6854;
wire     [31:0] n6855;
wire     [31:0] n6856;
wire     [31:0] n6857;
wire     [31:0] n6858;
wire     [31:0] n6859;
wire     [31:0] n6860;
wire     [31:0] n6861;
wire     [31:0] n6862;
wire     [31:0] n6863;
wire     [31:0] n6864;
wire     [31:0] n6865;
wire     [31:0] n6866;
wire     [31:0] n6867;
wire     [31:0] n6868;
wire     [31:0] n6869;
wire     [31:0] n6870;
wire     [31:0] n6871;
wire     [31:0] n6872;
wire     [31:0] n6873;
wire     [31:0] n6874;
wire     [31:0] n6875;
wire     [31:0] n6876;
wire     [31:0] n6877;
wire     [31:0] n6878;
wire     [31:0] n6879;
wire     [31:0] n6880;
wire     [31:0] n6881;
wire     [31:0] n6882;
wire     [31:0] n6883;
wire     [31:0] n6884;
wire     [31:0] n6885;
wire     [31:0] n6886;
wire     [31:0] n6887;
wire     [31:0] n6888;
wire     [31:0] n6889;
wire     [31:0] n6890;
wire     [31:0] n6891;
wire     [31:0] n6892;
wire     [31:0] n6893;
wire     [31:0] n6894;
wire     [31:0] n6895;
wire     [31:0] n6896;
wire     [31:0] n6897;
wire     [31:0] n6898;
wire     [31:0] n6899;
wire     [31:0] n6900;
wire     [31:0] n6901;
wire     [31:0] n6902;
wire     [31:0] n6903;
wire     [31:0] n6904;
wire     [31:0] n6905;
wire     [31:0] n6906;
wire     [31:0] n6907;
wire     [31:0] n6908;
wire     [31:0] n6909;
wire     [31:0] n6910;
wire     [31:0] n6911;
wire     [31:0] n6912;
wire     [31:0] n6913;
wire     [31:0] n6914;
wire     [31:0] n6915;
wire     [31:0] n6916;
wire     [31:0] n6917;
wire     [31:0] n6918;
wire     [31:0] n6919;
wire     [31:0] n6920;
wire     [31:0] n6921;
wire     [31:0] n6922;
wire     [31:0] n6923;
wire     [31:0] n6924;
wire     [31:0] n6925;
wire     [31:0] n6926;
wire     [31:0] n6927;
wire     [31:0] n6928;
wire     [31:0] n6929;
wire     [31:0] n6930;
wire     [31:0] n6931;
wire     [31:0] n6932;
wire     [31:0] n6933;
wire     [31:0] n6934;
wire     [31:0] n6935;
wire     [31:0] n6936;
wire     [31:0] n6937;
wire     [31:0] n6938;
wire     [31:0] n6939;
wire     [31:0] n6940;
wire     [31:0] n6941;
wire     [31:0] n6942;
wire     [31:0] n6943;
wire     [31:0] n6944;
wire     [31:0] n6945;
wire     [31:0] n6946;
wire     [31:0] n6947;
wire     [31:0] n6948;
wire     [31:0] n6949;
wire     [31:0] n6950;
wire     [31:0] n6951;
wire     [31:0] n6952;
wire     [31:0] n6953;
wire     [31:0] n6954;
wire     [31:0] n6955;
wire     [31:0] n6956;
wire     [31:0] n6957;
wire     [31:0] n6958;
wire     [31:0] n6959;
wire     [31:0] n6960;
wire     [31:0] n6961;
wire     [31:0] n6962;
wire     [31:0] n6963;
wire     [31:0] n6964;
wire     [31:0] n6965;
wire     [31:0] n6966;
wire     [31:0] n6967;
wire     [31:0] n6968;
wire     [31:0] n6969;
wire     [31:0] n6970;
wire     [31:0] n6971;
wire     [31:0] n6972;
wire     [31:0] n6973;
wire     [31:0] n6974;
wire     [31:0] n6975;
wire     [31:0] n6976;
wire     [31:0] n6977;
wire     [31:0] n6978;
wire     [31:0] n6979;
wire     [31:0] n6980;
wire     [31:0] n6981;
wire     [31:0] n6982;
wire     [31:0] n6983;
wire     [31:0] n6984;
wire     [31:0] n6985;
wire     [31:0] n6986;
wire     [31:0] n6987;
wire     [31:0] n6988;
wire     [31:0] n6989;
wire     [31:0] n6990;
wire     [31:0] n6991;
wire     [31:0] n6992;
wire     [31:0] n6993;
wire     [31:0] n6994;
wire     [31:0] n6995;
wire     [31:0] n6996;
wire     [31:0] n6997;
wire     [31:0] n6998;
wire     [31:0] n6999;
wire     [31:0] n7000;
wire     [31:0] n7001;
wire     [31:0] n7002;
wire     [31:0] n7003;
wire     [31:0] n7004;
wire     [31:0] n7005;
wire     [31:0] n7006;
wire     [31:0] n7007;
wire     [31:0] n7008;
wire     [31:0] n7009;
wire     [31:0] n7010;
wire     [31:0] n7011;
wire     [31:0] n7012;
wire     [31:0] n7013;
wire     [31:0] n7014;
wire     [31:0] n7015;
wire     [31:0] n7016;
wire     [31:0] n7017;
wire     [31:0] n7018;
wire     [31:0] n7019;
wire     [31:0] n7020;
wire     [31:0] n7021;
wire     [31:0] n7022;
wire     [31:0] n7023;
wire     [31:0] n7024;
wire     [31:0] n7025;
wire     [31:0] n7026;
wire     [31:0] n7027;
wire     [31:0] n7028;
wire     [31:0] n7029;
wire     [31:0] n7030;
wire     [31:0] n7031;
wire     [31:0] n7032;
wire     [31:0] n7033;
wire     [31:0] n7034;
wire     [31:0] n7035;
wire     [31:0] n7036;
wire     [31:0] n7037;
wire     [31:0] n7038;
wire     [31:0] n7039;
wire     [31:0] n7040;
wire     [31:0] n7041;
wire     [31:0] n7042;
wire     [31:0] n7043;
wire     [31:0] n7044;
wire     [31:0] n7045;
wire     [31:0] n7046;
wire     [31:0] n7047;
wire     [31:0] n7048;
wire     [31:0] n7049;
wire     [31:0] n7050;
wire     [31:0] n7051;
wire     [31:0] n7052;
wire     [31:0] n7053;
wire     [31:0] n7054;
wire     [31:0] n7055;
wire     [31:0] n7056;
wire     [31:0] n7057;
wire     [31:0] n7058;
wire     [31:0] n7059;
wire     [31:0] n7060;
wire     [31:0] n7061;
wire     [31:0] n7062;
wire     [31:0] n7063;
wire     [31:0] n7064;
wire     [31:0] n7065;
wire     [31:0] n7066;
wire     [31:0] n7067;
wire     [31:0] n7068;
wire     [31:0] n7069;
wire     [31:0] n7070;
wire     [31:0] n7071;
wire     [31:0] n7072;
wire     [31:0] n7073;
wire     [31:0] n7074;
wire     [31:0] n7075;
wire     [31:0] n7076;
wire     [31:0] n7077;
wire     [31:0] n7078;
wire     [31:0] n7079;
wire     [31:0] n7080;
wire     [31:0] n7081;
wire     [31:0] n7082;
wire     [31:0] n7083;
wire     [31:0] n7084;
wire     [31:0] n7085;
wire     [31:0] n7086;
wire     [31:0] n7087;
wire     [31:0] n7088;
wire     [31:0] n7089;
wire     [31:0] n7090;
wire     [31:0] n7091;
wire     [31:0] n7092;
wire     [31:0] n7093;
wire     [31:0] n7094;
wire     [31:0] n7095;
wire     [31:0] n7096;
wire     [31:0] n7097;
wire     [31:0] n7098;
wire     [31:0] n7099;
wire     [31:0] n7100;
wire     [31:0] n7101;
wire     [31:0] n7102;
wire     [31:0] n7103;
wire     [31:0] n7104;
wire     [31:0] n7105;
wire     [31:0] n7106;
wire     [31:0] n7107;
wire     [31:0] n7108;
wire     [31:0] n7109;
wire     [31:0] n7110;
wire     [31:0] n7111;
wire     [31:0] n7112;
wire     [31:0] n7113;
wire     [31:0] n7114;
wire     [31:0] n7115;
wire     [31:0] n7116;
wire     [31:0] n7117;
wire     [31:0] n7118;
wire     [31:0] n7119;
wire     [31:0] n7120;
wire     [31:0] n7121;
wire     [31:0] n7122;
wire     [31:0] n7123;
wire     [31:0] n7124;
wire     [31:0] n7125;
wire     [31:0] n7126;
wire     [31:0] n7127;
wire     [31:0] n7128;
wire     [31:0] n7129;
wire     [31:0] n7130;
wire     [31:0] n7131;
wire     [31:0] n7132;
wire     [31:0] n7133;
wire     [31:0] n7134;
wire     [31:0] n7135;
wire     [31:0] n7136;
wire     [31:0] n7137;
wire     [31:0] n7138;
wire     [31:0] n7139;
wire     [31:0] n7140;
wire     [31:0] n7141;
wire     [31:0] n7142;
wire     [31:0] n7143;
wire     [31:0] n7144;
wire     [31:0] n7145;
wire     [31:0] n7146;
wire     [31:0] n7147;
wire     [31:0] n7148;
wire     [31:0] n7149;
wire     [31:0] n7150;
wire     [31:0] n7151;
wire     [31:0] n7152;
wire     [31:0] n7153;
wire     [31:0] n7154;
wire     [31:0] n7155;
wire     [31:0] n7156;
wire     [31:0] n7157;
wire     [31:0] n7158;
wire     [31:0] n7159;
wire     [31:0] n7160;
wire     [31:0] n7161;
wire     [31:0] n7162;
wire     [31:0] n7163;
wire     [31:0] n7164;
wire     [31:0] n7165;
wire     [31:0] n7166;
wire     [31:0] n7167;
wire     [31:0] n7168;
wire     [31:0] n7169;
wire     [31:0] n7170;
wire     [31:0] n7171;
wire     [31:0] n7172;
wire     [31:0] n7173;
wire     [31:0] n7174;
wire     [31:0] n7175;
wire     [31:0] n7176;
wire     [31:0] n7177;
wire     [31:0] n7178;
wire     [31:0] n7179;
wire     [31:0] n7180;
wire     [31:0] n7181;
wire     [31:0] n7182;
wire     [31:0] n7183;
wire     [31:0] n7184;
wire     [31:0] n7185;
wire     [31:0] n7186;
wire     [31:0] n7187;
wire     [31:0] n7188;
wire     [31:0] n7189;
wire     [31:0] n7190;
wire     [31:0] n7191;
wire     [31:0] n7192;
wire     [31:0] n7193;
wire     [31:0] n7194;
wire     [31:0] n7195;
wire     [31:0] n7196;
wire     [31:0] n7197;
wire     [31:0] n7198;
wire     [31:0] n7199;
wire     [31:0] n7200;
wire     [31:0] n7201;
wire     [31:0] n7202;
wire     [31:0] n7203;
wire     [31:0] n7204;
wire     [31:0] n7205;
wire     [31:0] n7206;
wire     [31:0] n7207;
wire     [31:0] n7208;
wire     [31:0] n7209;
wire     [31:0] n7210;
wire     [31:0] n7211;
wire     [31:0] n7212;
wire     [31:0] n7213;
wire     [31:0] n7214;
wire     [31:0] n7215;
wire     [31:0] n7216;
wire     [31:0] n7217;
wire     [31:0] n7218;
wire     [31:0] n7219;
wire     [31:0] n7220;
wire     [31:0] n7221;
wire     [31:0] n7222;
wire     [31:0] n7223;
wire     [31:0] n7224;
wire     [31:0] n7225;
wire     [31:0] n7226;
wire     [31:0] n7227;
wire     [31:0] n7228;
wire     [31:0] n7229;
wire     [31:0] n7230;
wire     [31:0] n7231;
wire     [31:0] n7232;
wire     [31:0] n7233;
wire     [31:0] n7234;
wire     [31:0] n7235;
wire     [31:0] n7236;
wire     [31:0] n7237;
wire     [31:0] n7238;
wire     [31:0] n7239;
wire     [31:0] n7240;
wire     [31:0] n7241;
wire     [31:0] n7242;
wire     [31:0] n7243;
wire     [31:0] n7244;
wire     [31:0] n7245;
wire     [31:0] n7246;
wire     [31:0] n7247;
wire     [31:0] n7248;
wire     [31:0] n7249;
wire     [31:0] n7250;
wire     [31:0] n7251;
wire     [31:0] n7252;
wire     [31:0] n7253;
wire     [31:0] n7254;
wire     [31:0] n7255;
wire     [31:0] n7256;
wire     [31:0] n7257;
wire     [31:0] n7258;
wire     [31:0] n7259;
wire     [31:0] n7260;
wire     [31:0] n7261;
wire     [31:0] n7262;
wire     [31:0] n7263;
wire     [31:0] n7264;
wire     [31:0] n7265;
wire     [31:0] n7266;
wire     [31:0] n7267;
wire     [31:0] n7268;
wire     [31:0] n7269;
wire     [31:0] n7270;
wire     [31:0] n7271;
wire            n7272;
wire            n7273;
wire     [31:0] n7274;
wire     [31:0] n7275;
wire     [31:0] n7276;
wire     [31:0] n7277;
wire     [31:0] n7278;
wire     [31:0] n7279;
wire     [31:0] n7280;
wire     [31:0] n7281;
wire     [31:0] n7282;
wire     [31:0] n7283;
wire     [31:0] n7284;
wire     [31:0] n7285;
wire     [31:0] n7286;
wire     [31:0] n7287;
wire     [31:0] n7288;
wire     [31:0] n7289;
wire     [31:0] n7290;
wire     [31:0] n7291;
wire     [31:0] n7292;
wire     [31:0] n7293;
wire     [31:0] n7294;
wire     [31:0] n7295;
wire     [31:0] n7296;
wire     [31:0] n7297;
wire     [31:0] n7298;
wire     [31:0] n7299;
wire     [31:0] n7300;
wire     [31:0] n7301;
wire     [31:0] n7302;
wire     [31:0] n7303;
wire     [31:0] n7304;
wire     [31:0] n7305;
wire     [31:0] n7306;
wire            n7307;
wire            n7308;
wire            n7309;
wire            n7310;
wire            n7311;
wire            n7312;
wire            n7313;
wire            n7314;
wire            n7315;
wire            n7316;
wire            n7317;
wire            n7318;
wire            n7319;
wire            n7320;
wire            n7321;
wire            n7322;
wire            n7323;
wire            n7324;
wire            n7325;
wire            n7326;
wire            n7327;
wire            n7328;
wire            n7329;
wire            n7330;
wire            n7331;
wire            n7332;
wire            n7333;
wire            n7334;
wire            n7335;
wire            n7336;
wire            n7337;
wire            n7338;
wire            n7339;
wire            n7340;
wire            n7341;
wire            n7342;
wire            n7343;
wire            n7344;
wire            n7345;
wire            n7346;
wire            n7347;
wire            n7348;
wire            n7349;
wire            n7350;
wire            n7351;
wire            n7352;
wire            n7353;
wire            n7354;
wire            n7355;
wire            n7356;
wire            n7357;
wire            n7358;
wire            n7359;
wire            n7360;
wire            n7361;
wire            n7362;
wire            n7363;
wire            n7364;
wire            n7365;
wire            n7366;
wire            n7367;
wire            n7368;
wire            n7369;
wire            n7370;
wire            n7371;
wire            n7372;
wire            n7373;
wire            n7374;
wire            n7375;
wire            n7376;
wire            n7377;
wire            n7378;
wire            n7379;
wire            n7380;
wire            n7381;
wire            n7382;
wire            n7383;
wire            n7384;
wire            n7385;
wire            n7386;
wire            n7387;
wire            n7388;
wire            n7389;
wire            n7390;
wire            n7391;
wire            n7392;
wire            n7393;
wire            n7394;
wire            n7395;
wire            n7396;
wire            n7397;
wire            n7398;
wire            n7399;
wire            n7400;
wire            n7401;
wire            n7402;
wire            n7403;
wire            n7404;
wire            n7405;
wire            n7406;
wire            n7407;
wire            n7408;
wire            n7409;
wire            n7410;
wire            n7411;
wire            n7412;
wire            n7413;
wire            n7414;
wire            n7415;
wire            n7416;
wire            n7417;
wire            n7418;
wire            n7419;
wire            n7420;
wire            n7421;
wire            n7422;
wire            n7423;
wire            n7424;
wire            n7425;
wire            n7426;
wire            n7427;
wire            n7428;
wire            n7429;
wire            n7430;
wire            n7431;
wire            n7432;
wire            n7433;
wire            n7434;
wire            n7435;
wire            n7436;
wire            n7437;
wire            n7438;
wire            n7439;
wire            n7440;
wire            n7441;
wire            n7442;
wire            n7443;
wire            n7444;
wire            n7445;
wire            n7446;
wire            n7447;
wire            n7448;
wire            n7449;
wire            n7450;
wire            n7451;
wire            n7452;
wire            n7453;
wire            n7454;
wire            n7455;
wire            n7456;
wire            n7457;
wire            n7458;
wire            n7459;
wire            n7460;
wire            n7461;
wire            n7462;
wire            n7463;
wire            n7464;
wire            n7465;
wire            n7466;
wire            n7467;
wire            n7468;
wire            n7469;
wire            n7470;
wire            n7471;
wire            n7472;
wire            n7473;
wire            n7474;
wire            n7475;
wire            n7476;
wire            n7477;
wire            n7478;
wire            n7479;
wire            n7480;
wire            n7481;
wire            n7482;
wire            n7483;
wire            n7484;
wire            n7485;
wire            n7486;
wire            n7487;
wire            n7488;
wire            n7489;
wire            n7490;
wire            n7491;
wire            n7492;
wire            n7493;
wire            n7494;
wire            n7495;
wire            n7496;
wire            n7497;
wire            n7498;
wire            n7499;
wire            n7500;
wire            n7501;
wire            n7502;
wire            n7503;
wire            n7504;
wire            n7505;
wire            n7506;
wire            n7507;
wire            n7508;
wire            n7509;
wire            n7510;
wire            n7511;
wire            n7512;
wire            n7513;
wire            n7514;
wire            n7515;
wire            n7516;
wire            n7517;
wire            n7518;
wire            n7519;
wire            n7520;
wire            n7521;
wire            n7522;
wire            n7523;
wire            n7524;
wire            n7525;
wire            n7526;
wire            n7527;
wire            n7528;
wire            n7529;
wire            n7530;
wire            n7531;
wire            n7532;
wire            n7533;
wire            n7534;
wire            n7535;
wire            n7536;
wire            n7537;
wire            n7538;
wire            n7539;
wire            n7540;
wire            n7541;
wire            n7542;
wire            n7543;
wire            n7544;
wire            n7545;
wire            n7546;
wire            n7547;
wire            n7548;
wire            n7549;
wire            n7550;
wire            n7551;
wire            n7552;
wire            n7553;
wire            n7554;
wire            n7555;
wire            n7556;
wire            n7557;
wire            n7558;
wire            n7559;
wire            n7560;
wire            n7561;
wire            n7562;
wire            n7563;
wire            n7564;
wire            n7565;
wire            n7566;
wire            n7567;
wire            n7568;
wire            n7569;
wire            n7570;
wire            n7571;
wire            n7572;
wire            n7573;
wire            n7574;
wire            n7575;
wire            n7576;
wire            n7577;
wire            n7578;
wire            n7579;
wire            n7580;
wire            n7581;
wire            n7582;
wire            n7583;
wire            n7584;
wire            n7585;
wire            n7586;
wire            n7587;
wire            n7588;
wire            n7589;
wire            n7590;
wire            n7591;
wire            n7592;
wire            n7593;
wire            n7594;
wire            n7595;
wire            n7596;
wire            n7597;
wire            n7598;
wire            n7599;
wire            n7600;
wire            n7601;
wire            n7602;
wire            n7603;
wire            n7604;
wire            n7605;
wire            n7606;
wire            n7607;
wire            n7608;
wire            n7609;
wire            n7610;
wire            n7611;
wire            n7612;
wire            n7613;
wire            n7614;
wire            n7615;
wire            n7616;
wire            n7617;
wire            n7618;
wire            n7619;
wire            n7620;
wire            n7621;
wire            n7622;
wire            n7623;
wire            n7624;
wire            n7625;
wire            n7626;
wire            n7627;
wire            n7628;
wire            n7629;
wire            n7630;
wire            n7631;
wire            n7632;
wire            n7633;
wire            n7634;
wire            n7635;
wire            n7636;
wire            n7637;
wire            n7638;
wire            n7639;
wire            n7640;
wire            n7641;
wire            n7642;
wire            n7643;
wire            n7644;
wire            n7645;
wire            n7646;
wire            n7647;
wire            n7648;
wire            n7649;
wire            n7650;
wire            n7651;
wire            n7652;
wire            n7653;
wire            n7654;
wire            n7655;
wire            n7656;
wire            n7657;
wire            n7658;
wire            n7659;
wire            n7660;
wire            n7661;
wire            n7662;
wire            n7663;
wire            n7664;
wire            n7665;
wire            n7666;
wire            n7667;
wire            n7668;
wire            n7669;
wire            n7670;
wire            n7671;
wire            n7672;
wire            n7673;
wire            n7674;
wire            n7675;
wire            n7676;
wire            n7677;
wire            n7678;
wire            n7679;
wire            n7680;
wire            n7681;
wire            n7682;
wire            n7683;
wire            n7684;
wire            n7685;
wire            n7686;
wire            n7687;
wire            n7688;
wire            n7689;
wire            n7690;
wire            n7691;
wire            n7692;
wire            n7693;
wire            n7694;
wire            n7695;
wire            n7696;
wire            n7697;
wire            n7698;
wire            n7699;
wire            n7700;
wire            n7701;
wire            n7702;
wire            n7703;
wire            n7704;
wire            n7705;
wire            n7706;
wire            n7707;
wire            n7708;
wire            n7709;
wire            n7710;
wire            n7711;
wire            n7712;
wire            n7713;
wire            n7714;
wire            n7715;
wire            n7716;
wire            n7717;
wire            n7718;
wire            n7719;
wire            n7720;
wire            n7721;
wire            n7722;
wire            n7723;
wire            n7724;
wire            n7725;
wire            n7726;
wire            n7727;
wire            n7728;
wire            n7729;
wire            n7730;
wire            n7731;
wire            n7732;
wire            n7733;
wire            n7734;
wire            n7735;
wire            n7736;
wire            n7737;
wire            n7738;
wire            n7739;
wire            n7740;
wire            n7741;
wire            n7742;
wire            n7743;
wire            n7744;
wire            n7745;
wire            n7746;
wire            n7747;
wire            n7748;
wire            n7749;
wire            n7750;
wire            n7751;
wire            n7752;
wire            n7753;
wire            n7754;
wire            n7755;
wire            n7756;
wire            n7757;
wire            n7758;
wire            n7759;
wire            n7760;
wire            n7761;
wire            n7762;
wire            n7763;
wire            n7764;
wire            n7765;
wire            n7766;
wire            n7767;
wire            n7768;
wire            n7769;
wire            n7770;
wire            n7771;
wire            n7772;
wire            n7773;
wire            n7774;
wire            n7775;
wire            n7776;
wire            n7777;
wire            n7778;
wire            n7779;
wire            n7780;
wire            n7781;
wire            n7782;
wire            n7783;
wire            n7784;
wire            n7785;
wire            n7786;
wire            n7787;
wire            n7788;
wire            n7789;
wire            n7790;
wire            n7791;
wire            n7792;
wire            n7793;
wire            n7794;
wire            n7795;
wire            n7796;
wire            n7797;
wire            n7798;
wire            n7799;
wire            n7800;
wire            n7801;
wire            n7802;
wire            n7803;
wire            n7804;
wire            n7805;
wire            n7806;
wire            n7807;
wire            n7808;
wire            n7809;
wire            n7810;
wire            n7811;
wire            n7812;
wire            n7813;
wire            n7814;
wire            n7815;
wire            n7816;
wire            n7817;
wire            n7818;
wire            n7819;
wire            n7820;
wire            n7821;
wire            n7822;
wire            n7823;
wire            n7824;
wire            n7825;
wire            n7826;
wire            n7827;
wire            n7828;
wire            n7829;
wire            n7830;
wire            n7831;
wire            n7832;
wire            n7833;
wire            n7834;
wire     [31:0] n7835;
wire     [31:0] n7836;
wire     [31:0] n7837;
wire     [31:0] n7838;
wire     [31:0] n7839;
wire     [31:0] n7840;
wire     [31:0] n7841;
wire     [31:0] n7842;
wire     [31:0] n7843;
wire     [31:0] n7844;
wire     [31:0] n7845;
wire     [31:0] n7846;
wire     [31:0] n7847;
wire     [31:0] n7848;
wire     [31:0] n7849;
wire     [31:0] n7850;
wire     [31:0] n7851;
wire     [31:0] n7852;
wire     [31:0] n7853;
wire     [31:0] n7854;
wire     [31:0] n7855;
wire     [31:0] n7856;
wire     [31:0] n7857;
wire     [31:0] n7858;
wire     [31:0] n7859;
wire     [31:0] n7860;
wire     [31:0] n7861;
wire     [31:0] n7862;
wire     [31:0] n7863;
wire     [31:0] n7864;
wire     [31:0] n7865;
wire     [31:0] n7866;
wire     [31:0] n7867;
wire     [31:0] n7868;
wire     [31:0] n7869;
wire     [31:0] n7870;
wire     [31:0] n7871;
wire     [31:0] n7872;
wire     [31:0] n7873;
wire     [31:0] n7874;
wire     [31:0] n7875;
wire     [31:0] n7876;
wire     [31:0] n7877;
wire     [31:0] n7878;
wire     [31:0] n7879;
wire     [31:0] n7880;
wire     [31:0] n7881;
wire     [31:0] n7882;
wire     [31:0] n7883;
wire     [31:0] n7884;
wire     [31:0] n7885;
wire     [31:0] n7886;
wire     [31:0] n7887;
wire     [31:0] n7888;
wire     [31:0] n7889;
wire     [31:0] n7890;
wire     [31:0] n7891;
wire     [31:0] n7892;
wire     [31:0] n7893;
wire     [31:0] n7894;
wire     [31:0] n7895;
wire     [31:0] n7896;
wire     [31:0] n7897;
wire     [31:0] n7898;
wire     [31:0] n7899;
wire     [31:0] n7900;
wire     [31:0] n7901;
wire     [31:0] n7902;
wire     [31:0] n7903;
wire     [31:0] n7904;
wire     [31:0] n7905;
wire     [31:0] n7906;
wire     [31:0] n7907;
wire     [31:0] n7908;
wire     [31:0] n7909;
wire     [31:0] n7910;
wire     [31:0] n7911;
wire     [31:0] n7912;
wire     [31:0] n7913;
wire     [31:0] n7914;
wire     [31:0] n7915;
wire     [31:0] n7916;
wire     [31:0] n7917;
wire     [31:0] n7918;
wire     [31:0] n7919;
wire     [31:0] n7920;
wire     [31:0] n7921;
wire     [31:0] n7922;
wire     [31:0] n7923;
wire     [31:0] n7924;
wire     [31:0] n7925;
wire     [31:0] n7926;
wire     [31:0] n7927;
wire     [31:0] n7928;
wire     [31:0] n7929;
wire     [31:0] n7930;
wire     [31:0] n7931;
wire     [31:0] n7932;
wire     [31:0] n7933;
wire     [31:0] n7934;
wire     [31:0] n7935;
wire     [31:0] n7936;
wire     [31:0] n7937;
wire     [31:0] n7938;
wire     [31:0] n7939;
wire     [31:0] n7940;
wire     [31:0] n7941;
wire     [31:0] n7942;
wire     [31:0] n7943;
wire     [31:0] n7944;
wire     [31:0] n7945;
wire     [31:0] n7946;
wire     [31:0] n7947;
wire     [31:0] n7948;
wire     [31:0] n7949;
wire     [31:0] n7950;
wire     [31:0] n7951;
wire     [31:0] n7952;
wire     [31:0] n7953;
wire     [31:0] n7954;
wire     [31:0] n7955;
wire     [31:0] n7956;
wire     [31:0] n7957;
wire     [31:0] n7958;
wire     [31:0] n7959;
wire     [31:0] n7960;
wire     [31:0] n7961;
wire     [31:0] n7962;
wire     [31:0] n7963;
wire     [31:0] n7964;
wire     [31:0] n7965;
wire     [31:0] n7966;
wire     [31:0] n7967;
wire     [31:0] n7968;
wire     [31:0] n7969;
wire     [31:0] n7970;
wire     [31:0] n7971;
wire     [31:0] n7972;
wire     [31:0] n7973;
wire     [31:0] n7974;
wire     [31:0] n7975;
wire     [31:0] n7976;
wire     [31:0] n7977;
wire     [31:0] n7978;
wire     [31:0] n7979;
wire     [31:0] n7980;
wire     [31:0] n7981;
wire     [31:0] n7982;
wire     [31:0] n7983;
wire     [31:0] n7984;
wire     [31:0] n7985;
wire     [31:0] n7986;
wire     [31:0] n7987;
wire     [31:0] n7988;
wire     [31:0] n7989;
wire     [31:0] n7990;
wire     [31:0] n7991;
wire     [31:0] n7992;
wire     [31:0] n7993;
wire     [31:0] n7994;
wire     [31:0] n7995;
wire     [31:0] n7996;
wire     [31:0] n7997;
wire     [31:0] n7998;
wire     [31:0] n7999;
wire     [31:0] n8000;
wire     [31:0] n8001;
wire     [31:0] n8002;
wire     [31:0] n8003;
wire     [31:0] n8004;
wire     [31:0] n8005;
wire     [31:0] n8006;
wire     [31:0] n8007;
wire     [31:0] n8008;
wire     [31:0] n8009;
wire     [31:0] n8010;
wire     [31:0] n8011;
wire     [31:0] n8012;
wire     [31:0] n8013;
wire     [31:0] n8014;
wire     [31:0] n8015;
wire     [31:0] n8016;
wire     [31:0] n8017;
wire     [31:0] n8018;
wire     [31:0] n8019;
wire     [31:0] n8020;
wire     [31:0] n8021;
wire     [31:0] n8022;
wire     [31:0] n8023;
wire     [31:0] n8024;
wire     [31:0] n8025;
wire     [31:0] n8026;
wire     [31:0] n8027;
wire     [31:0] n8028;
wire     [31:0] n8029;
wire     [31:0] n8030;
wire     [31:0] n8031;
wire     [31:0] n8032;
wire     [31:0] n8033;
wire     [31:0] n8034;
wire     [31:0] n8035;
wire     [31:0] n8036;
wire     [31:0] n8037;
wire     [31:0] n8038;
wire     [31:0] n8039;
wire     [31:0] n8040;
wire     [31:0] n8041;
wire     [31:0] n8042;
wire     [31:0] n8043;
wire     [31:0] n8044;
wire     [31:0] n8045;
wire     [31:0] n8046;
wire     [31:0] n8047;
wire     [31:0] n8048;
wire     [31:0] n8049;
wire     [31:0] n8050;
wire     [31:0] n8051;
wire     [31:0] n8052;
wire     [31:0] n8053;
wire     [31:0] n8054;
wire     [31:0] n8055;
wire     [31:0] n8056;
wire     [31:0] n8057;
wire     [31:0] n8058;
wire     [31:0] n8059;
wire     [31:0] n8060;
wire     [31:0] n8061;
wire     [31:0] n8062;
wire     [31:0] n8063;
wire     [31:0] n8064;
wire     [31:0] n8065;
wire     [31:0] n8066;
wire     [31:0] n8067;
wire     [31:0] n8068;
wire     [31:0] n8069;
wire     [31:0] n8070;
wire     [31:0] n8071;
wire     [31:0] n8072;
wire     [31:0] n8073;
wire     [31:0] n8074;
wire     [31:0] n8075;
wire     [31:0] n8076;
wire     [31:0] n8077;
wire     [31:0] n8078;
wire     [31:0] n8079;
wire     [31:0] n8080;
wire     [31:0] n8081;
wire     [31:0] n8082;
wire     [31:0] n8083;
wire     [31:0] n8084;
wire     [31:0] n8085;
wire     [31:0] n8086;
wire     [31:0] n8087;
wire     [31:0] n8088;
wire     [31:0] n8089;
wire     [31:0] n8090;
wire     [31:0] n8091;
wire     [31:0] n8092;
wire     [31:0] n8093;
wire     [31:0] n8094;
wire     [31:0] n8095;
wire     [31:0] n8096;
wire     [31:0] n8097;
wire     [31:0] n8098;
wire     [31:0] n8099;
wire     [31:0] n8100;
wire     [31:0] n8101;
wire     [31:0] n8102;
wire     [31:0] n8103;
wire     [31:0] n8104;
wire     [31:0] n8105;
wire     [31:0] n8106;
wire     [31:0] n8107;
wire     [31:0] n8108;
wire     [31:0] n8109;
wire     [31:0] n8110;
wire     [31:0] n8111;
wire     [31:0] n8112;
wire     [31:0] n8113;
wire     [31:0] n8114;
wire     [31:0] n8115;
wire     [31:0] n8116;
wire     [31:0] n8117;
wire     [31:0] n8118;
wire     [31:0] n8119;
wire     [31:0] n8120;
wire     [31:0] n8121;
wire     [31:0] n8122;
wire     [31:0] n8123;
wire     [31:0] n8124;
wire     [31:0] n8125;
wire     [31:0] n8126;
wire     [31:0] n8127;
wire     [31:0] n8128;
wire     [31:0] n8129;
wire     [31:0] n8130;
wire     [31:0] n8131;
wire     [31:0] n8132;
wire     [31:0] n8133;
wire     [31:0] n8134;
wire     [31:0] n8135;
wire     [31:0] n8136;
wire     [31:0] n8137;
wire     [31:0] n8138;
wire     [31:0] n8139;
wire     [31:0] n8140;
wire     [31:0] n8141;
wire     [31:0] n8142;
wire     [31:0] n8143;
wire     [31:0] n8144;
wire     [31:0] n8145;
wire     [31:0] n8146;
wire     [31:0] n8147;
wire     [31:0] n8148;
wire     [31:0] n8149;
wire     [31:0] n8150;
wire     [31:0] n8151;
wire     [31:0] n8152;
wire     [31:0] n8153;
wire     [31:0] n8154;
wire     [31:0] n8155;
wire     [31:0] n8156;
wire     [31:0] n8157;
wire     [31:0] n8158;
wire     [31:0] n8159;
wire     [31:0] n8160;
wire     [31:0] n8161;
wire     [31:0] n8162;
wire     [31:0] n8163;
wire     [31:0] n8164;
wire     [31:0] n8165;
wire     [31:0] n8166;
wire     [31:0] n8167;
wire     [31:0] n8168;
wire     [31:0] n8169;
wire     [31:0] n8170;
wire     [31:0] n8171;
wire     [31:0] n8172;
wire     [31:0] n8173;
wire     [31:0] n8174;
wire     [31:0] n8175;
wire     [31:0] n8176;
wire     [31:0] n8177;
wire     [31:0] n8178;
wire     [31:0] n8179;
wire     [31:0] n8180;
wire     [31:0] n8181;
wire     [31:0] n8182;
wire     [31:0] n8183;
wire     [31:0] n8184;
wire     [31:0] n8185;
wire     [31:0] n8186;
wire     [31:0] n8187;
wire     [31:0] n8188;
wire     [31:0] n8189;
wire     [31:0] n8190;
wire     [31:0] n8191;
wire     [31:0] n8192;
wire     [31:0] n8193;
wire     [31:0] n8194;
wire     [31:0] n8195;
wire     [31:0] n8196;
wire     [31:0] n8197;
wire     [31:0] n8198;
wire     [31:0] n8199;
wire     [31:0] n8200;
wire     [31:0] n8201;
wire     [31:0] n8202;
wire     [31:0] n8203;
wire     [31:0] n8204;
wire     [31:0] n8205;
wire     [31:0] n8206;
wire     [31:0] n8207;
wire     [31:0] n8208;
wire     [31:0] n8209;
wire     [31:0] n8210;
wire     [31:0] n8211;
wire     [31:0] n8212;
wire     [31:0] n8213;
wire     [31:0] n8214;
wire     [31:0] n8215;
wire     [31:0] n8216;
wire     [31:0] n8217;
wire     [31:0] n8218;
wire     [31:0] n8219;
wire     [31:0] n8220;
wire     [31:0] n8221;
wire     [31:0] n8222;
wire     [31:0] n8223;
wire     [31:0] n8224;
wire     [31:0] n8225;
wire     [31:0] n8226;
wire     [31:0] n8227;
wire     [31:0] n8228;
wire     [31:0] n8229;
wire     [31:0] n8230;
wire     [31:0] n8231;
wire     [31:0] n8232;
wire     [31:0] n8233;
wire     [31:0] n8234;
wire     [31:0] n8235;
wire     [31:0] n8236;
wire     [31:0] n8237;
wire     [31:0] n8238;
wire     [31:0] n8239;
wire     [31:0] n8240;
wire     [31:0] n8241;
wire     [31:0] n8242;
wire     [31:0] n8243;
wire     [31:0] n8244;
wire     [31:0] n8245;
wire     [31:0] n8246;
wire     [31:0] n8247;
wire     [31:0] n8248;
wire     [31:0] n8249;
wire     [31:0] n8250;
wire     [31:0] n8251;
wire     [31:0] n8252;
wire     [31:0] n8253;
wire     [31:0] n8254;
wire     [31:0] n8255;
wire     [31:0] n8256;
wire     [31:0] n8257;
wire     [31:0] n8258;
wire     [31:0] n8259;
wire     [31:0] n8260;
wire     [31:0] n8261;
wire     [31:0] n8262;
wire     [31:0] n8263;
wire     [31:0] n8264;
wire     [31:0] n8265;
wire     [31:0] n8266;
wire     [31:0] n8267;
wire     [31:0] n8268;
wire     [31:0] n8269;
wire     [31:0] n8270;
wire     [31:0] n8271;
wire     [31:0] n8272;
wire     [31:0] n8273;
wire     [31:0] n8274;
wire     [31:0] n8275;
wire     [31:0] n8276;
wire     [31:0] n8277;
wire     [31:0] n8278;
wire     [31:0] n8279;
wire     [31:0] n8280;
wire     [31:0] n8281;
wire     [31:0] n8282;
wire     [31:0] n8283;
wire     [31:0] n8284;
wire     [31:0] n8285;
wire     [31:0] n8286;
wire     [31:0] n8287;
wire     [31:0] n8288;
wire     [31:0] n8289;
wire     [31:0] n8290;
wire     [31:0] n8291;
wire     [31:0] n8292;
wire     [31:0] n8293;
wire     [31:0] n8294;
wire     [31:0] n8295;
wire     [31:0] n8296;
wire     [31:0] n8297;
wire     [31:0] n8298;
wire     [31:0] n8299;
wire     [31:0] n8300;
wire     [31:0] n8301;
wire     [31:0] n8302;
wire     [31:0] n8303;
wire     [31:0] n8304;
wire     [31:0] n8305;
wire     [31:0] n8306;
wire     [31:0] n8307;
wire     [31:0] n8308;
wire     [31:0] n8309;
wire     [31:0] n8310;
wire     [31:0] n8311;
wire     [31:0] n8312;
wire     [31:0] n8313;
wire     [31:0] n8314;
wire     [31:0] n8315;
wire     [31:0] n8316;
wire     [31:0] n8317;
wire     [31:0] n8318;
wire     [31:0] n8319;
wire     [31:0] n8320;
wire     [31:0] n8321;
wire     [31:0] n8322;
wire     [31:0] n8323;
wire     [31:0] n8324;
wire     [31:0] n8325;
wire     [31:0] n8326;
wire     [31:0] n8327;
wire     [31:0] n8328;
wire     [31:0] n8329;
wire     [31:0] n8330;
wire     [31:0] n8331;
wire     [31:0] n8332;
wire     [31:0] n8333;
wire     [31:0] n8334;
wire     [31:0] n8335;
wire     [31:0] n8336;
wire     [31:0] n8337;
wire     [31:0] n8338;
wire     [31:0] n8339;
wire     [31:0] n8340;
wire     [31:0] n8341;
wire     [31:0] n8342;
wire     [31:0] n8343;
wire     [31:0] n8344;
wire     [31:0] n8345;
wire     [31:0] n8346;
wire     [31:0] n8347;
wire     [31:0] n8348;
wire     [31:0] n8349;
wire     [31:0] n8350;
wire     [31:0] n8351;
wire     [31:0] n8352;
wire     [31:0] n8353;
wire     [31:0] n8354;
wire     [31:0] n8355;
wire     [31:0] n8356;
wire            n8357;
wire            n8358;
wire            n8359;
wire            n8360;
wire            n8361;
wire            n8362;
wire            n8363;
wire            n8364;
wire            n8365;
wire            n8366;
wire            n8367;
wire            n8368;
wire            n8369;
wire            n8370;
wire            n8371;
wire            n8372;
wire            n8373;
wire            n8374;
wire            n8375;
wire            n8376;
wire            n8377;
wire            n8378;
wire            n8379;
wire            n8380;
wire            n8381;
wire            n8382;
wire            n8383;
wire            n8384;
wire            n8385;
wire            n8386;
wire            n8387;
wire            n8388;
wire            n8389;
wire            n8390;
wire            n8391;
wire            n8392;
wire            n8393;
wire            n8394;
wire            n8395;
wire            n8396;
wire            n8397;
wire            n8398;
wire            n8399;
wire            n8400;
wire            n8401;
wire            n8402;
wire            n8403;
wire            n8404;
wire            n8405;
wire            n8406;
wire            n8407;
wire            n8408;
wire            n8409;
wire            n8410;
wire            n8411;
wire            n8412;
wire            n8413;
wire            n8414;
wire            n8415;
wire            n8416;
wire            n8417;
wire            n8418;
wire            n8419;
wire            n8420;
wire            n8421;
wire            n8422;
wire            n8423;
wire            n8424;
wire            n8425;
wire            n8426;
wire            n8427;
wire            n8428;
wire            n8429;
wire            n8430;
wire            n8431;
wire            n8432;
wire            n8433;
wire            n8434;
wire            n8435;
wire            n8436;
wire            n8437;
wire            n8438;
wire            n8439;
wire            n8440;
wire            n8441;
wire            n8442;
wire            n8443;
wire            n8444;
wire            n8445;
wire            n8446;
wire            n8447;
wire            n8448;
wire            n8449;
wire            n8450;
wire            n8451;
wire            n8452;
wire            n8453;
wire            n8454;
wire            n8455;
wire            n8456;
wire            n8457;
wire            n8458;
wire            n8459;
wire            n8460;
wire            n8461;
wire            n8462;
wire            n8463;
wire            n8464;
wire            n8465;
wire            n8466;
wire            n8467;
wire            n8468;
wire            n8469;
wire            n8470;
wire            n8471;
wire            n8472;
wire            n8473;
wire            n8474;
wire            n8475;
wire            n8476;
wire            n8477;
wire            n8478;
wire            n8479;
wire            n8480;
wire            n8481;
wire            n8482;
wire            n8483;
wire            n8484;
wire            n8485;
wire            n8486;
wire            n8487;
wire            n8488;
wire            n8489;
wire            n8490;
wire            n8491;
wire            n8492;
wire            n8493;
wire            n8494;
wire            n8495;
wire            n8496;
wire            n8497;
wire            n8498;
wire            n8499;
wire            n8500;
wire            n8501;
wire            n8502;
wire            n8503;
wire            n8504;
wire            n8505;
wire            n8506;
wire            n8507;
wire            n8508;
wire            n8509;
wire            n8510;
wire            n8511;
wire            n8512;
wire            n8513;
wire            n8514;
wire            n8515;
wire            n8516;
wire            n8517;
wire            n8518;
wire            n8519;
wire            n8520;
wire            n8521;
wire            n8522;
wire            n8523;
wire            n8524;
wire            n8525;
wire            n8526;
wire            n8527;
wire            n8528;
wire            n8529;
wire            n8530;
wire            n8531;
wire            n8532;
wire            n8533;
wire            n8534;
wire            n8535;
wire            n8536;
wire            n8537;
wire            n8538;
wire            n8539;
wire            n8540;
wire            n8541;
wire            n8542;
wire            n8543;
wire            n8544;
wire            n8545;
wire            n8546;
wire            n8547;
wire            n8548;
wire            n8549;
wire            n8550;
wire            n8551;
wire            n8552;
wire            n8553;
wire            n8554;
wire            n8555;
wire            n8556;
wire            n8557;
wire            n8558;
wire            n8559;
wire            n8560;
wire            n8561;
wire            n8562;
wire            n8563;
wire            n8564;
wire            n8565;
wire            n8566;
wire            n8567;
wire            n8568;
wire            n8569;
wire            n8570;
wire            n8571;
wire            n8572;
wire            n8573;
wire            n8574;
wire            n8575;
wire            n8576;
wire            n8577;
wire            n8578;
wire            n8579;
wire            n8580;
wire            n8581;
wire            n8582;
wire            n8583;
wire            n8584;
wire            n8585;
wire            n8586;
wire            n8587;
wire            n8588;
wire            n8589;
wire            n8590;
wire            n8591;
wire            n8592;
wire            n8593;
wire            n8594;
wire            n8595;
wire            n8596;
wire            n8597;
wire            n8598;
wire            n8599;
wire            n8600;
wire            n8601;
wire            n8602;
wire            n8603;
wire            n8604;
wire            n8605;
wire            n8606;
wire            n8607;
wire            n8608;
wire            n8609;
wire            n8610;
wire            n8611;
wire            n8612;
wire            n8613;
wire            n8614;
wire            n8615;
wire            n8616;
wire            n8617;
wire            n8618;
wire            n8619;
wire            n8620;
wire            n8621;
wire            n8622;
wire            n8623;
wire            n8624;
wire            n8625;
wire            n8626;
wire            n8627;
wire            n8628;
wire            n8629;
wire            n8630;
wire            n8631;
wire            n8632;
wire            n8633;
wire            n8634;
wire            n8635;
wire            n8636;
wire            n8637;
wire            n8638;
wire            n8639;
wire            n8640;
wire            n8641;
wire            n8642;
wire            n8643;
wire            n8644;
wire            n8645;
wire            n8646;
wire            n8647;
wire            n8648;
wire            n8649;
wire            n8650;
wire            n8651;
wire            n8652;
wire            n8653;
wire            n8654;
wire            n8655;
wire            n8656;
wire            n8657;
wire            n8658;
wire            n8659;
wire            n8660;
wire            n8661;
wire            n8662;
wire            n8663;
wire            n8664;
wire            n8665;
wire            n8666;
wire            n8667;
wire            n8668;
wire            n8669;
wire            n8670;
wire            n8671;
wire            n8672;
wire            n8673;
wire            n8674;
wire            n8675;
wire            n8676;
wire            n8677;
wire            n8678;
wire            n8679;
wire            n8680;
wire            n8681;
wire            n8682;
wire            n8683;
wire            n8684;
wire            n8685;
wire            n8686;
wire            n8687;
wire            n8688;
wire            n8689;
wire            n8690;
wire            n8691;
wire            n8692;
wire            n8693;
wire            n8694;
wire            n8695;
wire            n8696;
wire            n8697;
wire            n8698;
wire            n8699;
wire            n8700;
wire            n8701;
wire            n8702;
wire            n8703;
wire            n8704;
wire            n8705;
wire            n8706;
wire            n8707;
wire            n8708;
wire            n8709;
wire            n8710;
wire            n8711;
wire            n8712;
wire            n8713;
wire            n8714;
wire            n8715;
wire            n8716;
wire            n8717;
wire            n8718;
wire            n8719;
wire            n8720;
wire            n8721;
wire            n8722;
wire            n8723;
wire            n8724;
wire            n8725;
wire            n8726;
wire            n8727;
wire            n8728;
wire            n8729;
wire            n8730;
wire            n8731;
wire            n8732;
wire            n8733;
wire            n8734;
wire            n8735;
wire            n8736;
wire            n8737;
wire            n8738;
wire            n8739;
wire            n8740;
wire            n8741;
wire            n8742;
wire            n8743;
wire            n8744;
wire            n8745;
wire            n8746;
wire            n8747;
wire            n8748;
wire            n8749;
wire            n8750;
wire            n8751;
wire            n8752;
wire            n8753;
wire            n8754;
wire            n8755;
wire            n8756;
wire            n8757;
wire            n8758;
wire            n8759;
wire            n8760;
wire            n8761;
wire            n8762;
wire            n8763;
wire            n8764;
wire            n8765;
wire            n8766;
wire            n8767;
wire            n8768;
wire            n8769;
wire            n8770;
wire            n8771;
wire            n8772;
wire            n8773;
wire            n8774;
wire            n8775;
wire            n8776;
wire            n8777;
wire            n8778;
wire            n8779;
wire            n8780;
wire            n8781;
wire            n8782;
wire            n8783;
wire            n8784;
wire            n8785;
wire            n8786;
wire            n8787;
wire            n8788;
wire            n8789;
wire            n8790;
wire            n8791;
wire            n8792;
wire            n8793;
wire            n8794;
wire            n8795;
wire            n8796;
wire            n8797;
wire            n8798;
wire            n8799;
wire            n8800;
wire            n8801;
wire            n8802;
wire            n8803;
wire            n8804;
wire            n8805;
wire            n8806;
wire            n8807;
wire            n8808;
wire            n8809;
wire            n8810;
wire            n8811;
wire            n8812;
wire            n8813;
wire            n8814;
wire            n8815;
wire            n8816;
wire            n8817;
wire            n8818;
wire            n8819;
wire            n8820;
wire            n8821;
wire            n8822;
wire            n8823;
wire            n8824;
wire            n8825;
wire            n8826;
wire            n8827;
wire            n8828;
wire            n8829;
wire            n8830;
wire            n8831;
wire            n8832;
wire            n8833;
wire            n8834;
wire            n8835;
wire            n8836;
wire            n8837;
wire            n8838;
wire            n8839;
wire            n8840;
wire            n8841;
wire            n8842;
wire            n8843;
wire            n8844;
wire            n8845;
wire            n8846;
wire            n8847;
wire            n8848;
wire            n8849;
wire            n8850;
wire            n8851;
wire            n8852;
wire            n8853;
wire            n8854;
wire            n8855;
wire            n8856;
wire            n8857;
wire            n8858;
wire            n8859;
wire            n8860;
wire            n8861;
wire            n8862;
wire            n8863;
wire            n8864;
wire            n8865;
wire            n8866;
wire            n8867;
wire            n8868;
wire     [31:0] n8869;
wire     [31:0] n8870;
wire     [31:0] n8871;
wire     [31:0] n8872;
wire     [31:0] n8873;
wire     [31:0] n8874;
wire     [31:0] n8875;
wire     [31:0] n8876;
wire     [31:0] n8877;
wire     [31:0] n8878;
wire     [31:0] n8879;
wire     [31:0] n8880;
wire     [31:0] n8881;
wire     [31:0] n8882;
wire     [31:0] n8883;
wire     [31:0] n8884;
wire     [31:0] n8885;
wire     [31:0] n8886;
wire     [31:0] n8887;
wire     [31:0] n8888;
wire     [31:0] n8889;
wire     [31:0] n8890;
wire     [31:0] n8891;
wire     [31:0] n8892;
wire     [31:0] n8893;
wire     [31:0] n8894;
wire     [31:0] n8895;
wire     [31:0] n8896;
wire     [31:0] n8897;
wire     [31:0] n8898;
wire     [31:0] n8899;
wire     [31:0] n8900;
wire     [31:0] n8901;
wire     [31:0] n8902;
wire     [31:0] n8903;
wire     [31:0] n8904;
wire     [31:0] n8905;
wire     [31:0] n8906;
wire     [31:0] n8907;
wire     [31:0] n8908;
wire     [31:0] n8909;
wire     [31:0] n8910;
wire     [31:0] n8911;
wire     [31:0] n8912;
wire     [31:0] n8913;
wire     [31:0] n8914;
wire     [31:0] n8915;
wire     [31:0] n8916;
wire     [31:0] n8917;
wire     [31:0] n8918;
wire     [31:0] n8919;
wire     [31:0] n8920;
wire     [31:0] n8921;
wire     [31:0] n8922;
wire     [31:0] n8923;
wire     [31:0] n8924;
wire     [31:0] n8925;
wire     [31:0] n8926;
wire     [31:0] n8927;
wire     [31:0] n8928;
wire     [31:0] n8929;
wire     [31:0] n8930;
wire     [31:0] n8931;
wire     [31:0] n8932;
wire     [31:0] n8933;
wire     [31:0] n8934;
wire     [31:0] n8935;
wire     [31:0] n8936;
wire     [31:0] n8937;
wire     [31:0] n8938;
wire     [31:0] n8939;
wire     [31:0] n8940;
wire     [31:0] n8941;
wire     [31:0] n8942;
wire     [31:0] n8943;
wire     [31:0] n8944;
wire     [31:0] n8945;
wire     [31:0] n8946;
wire     [31:0] n8947;
wire     [31:0] n8948;
wire     [31:0] n8949;
wire     [31:0] n8950;
wire     [31:0] n8951;
wire     [31:0] n8952;
wire     [31:0] n8953;
wire     [31:0] n8954;
wire     [31:0] n8955;
wire     [31:0] n8956;
wire     [31:0] n8957;
wire     [31:0] n8958;
wire     [31:0] n8959;
wire     [31:0] n8960;
wire     [31:0] n8961;
wire     [31:0] n8962;
wire     [31:0] n8963;
wire     [31:0] n8964;
wire     [31:0] n8965;
wire     [31:0] n8966;
wire     [31:0] n8967;
wire     [31:0] n8968;
wire     [31:0] n8969;
wire     [31:0] n8970;
wire     [31:0] n8971;
wire     [31:0] n8972;
wire     [31:0] n8973;
wire     [31:0] n8974;
wire     [31:0] n8975;
wire     [31:0] n8976;
wire     [31:0] n8977;
wire     [31:0] n8978;
wire     [31:0] n8979;
wire     [31:0] n8980;
wire     [31:0] n8981;
wire     [31:0] n8982;
wire     [31:0] n8983;
wire     [31:0] n8984;
wire     [31:0] n8985;
wire     [31:0] n8986;
wire     [31:0] n8987;
wire     [31:0] n8988;
wire     [31:0] n8989;
wire     [31:0] n8990;
wire     [31:0] n8991;
wire     [31:0] n8992;
wire     [31:0] n8993;
wire     [31:0] n8994;
wire     [31:0] n8995;
wire     [31:0] n8996;
wire     [31:0] n8997;
wire     [31:0] n8998;
wire     [31:0] n8999;
wire     [31:0] n9000;
wire     [31:0] n9001;
wire     [31:0] n9002;
wire     [31:0] n9003;
wire     [31:0] n9004;
wire     [31:0] n9005;
wire     [31:0] n9006;
wire     [31:0] n9007;
wire     [31:0] n9008;
wire     [31:0] n9009;
wire     [31:0] n9010;
wire     [31:0] n9011;
wire     [31:0] n9012;
wire     [31:0] n9013;
wire     [31:0] n9014;
wire     [31:0] n9015;
wire     [31:0] n9016;
wire     [31:0] n9017;
wire     [31:0] n9018;
wire     [31:0] n9019;
wire     [31:0] n9020;
wire     [31:0] n9021;
wire     [31:0] n9022;
wire     [31:0] n9023;
wire     [31:0] n9024;
wire     [31:0] n9025;
wire     [31:0] n9026;
wire     [31:0] n9027;
wire     [31:0] n9028;
wire     [31:0] n9029;
wire     [31:0] n9030;
wire     [31:0] n9031;
wire     [31:0] n9032;
wire     [31:0] n9033;
wire     [31:0] n9034;
wire     [31:0] n9035;
wire     [31:0] n9036;
wire     [31:0] n9037;
wire     [31:0] n9038;
wire     [31:0] n9039;
wire     [31:0] n9040;
wire     [31:0] n9041;
wire     [31:0] n9042;
wire     [31:0] n9043;
wire     [31:0] n9044;
wire     [31:0] n9045;
wire     [31:0] n9046;
wire     [31:0] n9047;
wire     [31:0] n9048;
wire     [31:0] n9049;
wire     [31:0] n9050;
wire     [31:0] n9051;
wire     [31:0] n9052;
wire     [31:0] n9053;
wire     [31:0] n9054;
wire     [31:0] n9055;
wire     [31:0] n9056;
wire     [31:0] n9057;
wire     [31:0] n9058;
wire     [31:0] n9059;
wire     [31:0] n9060;
wire     [31:0] n9061;
wire     [31:0] n9062;
wire     [31:0] n9063;
wire     [31:0] n9064;
wire     [31:0] n9065;
wire     [31:0] n9066;
wire     [31:0] n9067;
wire     [31:0] n9068;
wire     [31:0] n9069;
wire     [31:0] n9070;
wire     [31:0] n9071;
wire     [31:0] n9072;
wire     [31:0] n9073;
wire     [31:0] n9074;
wire     [31:0] n9075;
wire     [31:0] n9076;
wire     [31:0] n9077;
wire     [31:0] n9078;
wire     [31:0] n9079;
wire     [31:0] n9080;
wire     [31:0] n9081;
wire     [31:0] n9082;
wire     [31:0] n9083;
wire     [31:0] n9084;
wire     [31:0] n9085;
wire     [31:0] n9086;
wire     [31:0] n9087;
wire     [31:0] n9088;
wire     [31:0] n9089;
wire     [31:0] n9090;
wire     [31:0] n9091;
wire     [31:0] n9092;
wire     [31:0] n9093;
wire     [31:0] n9094;
wire     [31:0] n9095;
wire     [31:0] n9096;
wire     [31:0] n9097;
wire     [31:0] n9098;
wire     [31:0] n9099;
wire     [31:0] n9100;
wire     [31:0] n9101;
wire     [31:0] n9102;
wire     [31:0] n9103;
wire     [31:0] n9104;
wire     [31:0] n9105;
wire     [31:0] n9106;
wire     [31:0] n9107;
wire     [31:0] n9108;
wire     [31:0] n9109;
wire     [31:0] n9110;
wire     [31:0] n9111;
wire     [31:0] n9112;
wire     [31:0] n9113;
wire     [31:0] n9114;
wire     [31:0] n9115;
wire     [31:0] n9116;
wire     [31:0] n9117;
wire     [31:0] n9118;
wire     [31:0] n9119;
wire     [31:0] n9120;
wire     [31:0] n9121;
wire     [31:0] n9122;
wire     [31:0] n9123;
wire     [31:0] n9124;
wire     [31:0] n9125;
wire     [31:0] n9126;
wire     [31:0] n9127;
wire     [31:0] n9128;
wire     [31:0] n9129;
wire     [31:0] n9130;
wire     [31:0] n9131;
wire     [31:0] n9132;
wire     [31:0] n9133;
wire     [31:0] n9134;
wire     [31:0] n9135;
wire     [31:0] n9136;
wire     [31:0] n9137;
wire     [31:0] n9138;
wire     [31:0] n9139;
wire     [31:0] n9140;
wire     [31:0] n9141;
wire     [31:0] n9142;
wire     [31:0] n9143;
wire     [31:0] n9144;
wire     [31:0] n9145;
wire     [31:0] n9146;
wire     [31:0] n9147;
wire     [31:0] n9148;
wire     [31:0] n9149;
wire     [31:0] n9150;
wire     [31:0] n9151;
wire     [31:0] n9152;
wire     [31:0] n9153;
wire     [31:0] n9154;
wire     [31:0] n9155;
wire     [31:0] n9156;
wire     [31:0] n9157;
wire     [31:0] n9158;
wire     [31:0] n9159;
wire     [31:0] n9160;
wire     [31:0] n9161;
wire     [31:0] n9162;
wire     [31:0] n9163;
wire     [31:0] n9164;
wire     [31:0] n9165;
wire     [31:0] n9166;
wire     [31:0] n9167;
wire     [31:0] n9168;
wire     [31:0] n9169;
wire     [31:0] n9170;
wire     [31:0] n9171;
wire     [31:0] n9172;
wire     [31:0] n9173;
wire     [31:0] n9174;
wire     [31:0] n9175;
wire     [31:0] n9176;
wire     [31:0] n9177;
wire     [31:0] n9178;
wire     [31:0] n9179;
wire     [31:0] n9180;
wire     [31:0] n9181;
wire     [31:0] n9182;
wire     [31:0] n9183;
wire     [31:0] n9184;
wire     [31:0] n9185;
wire     [31:0] n9186;
wire     [31:0] n9187;
wire     [31:0] n9188;
wire     [31:0] n9189;
wire     [31:0] n9190;
wire     [31:0] n9191;
wire     [31:0] n9192;
wire     [31:0] n9193;
wire     [31:0] n9194;
wire     [31:0] n9195;
wire     [31:0] n9196;
wire     [31:0] n9197;
wire     [31:0] n9198;
wire     [31:0] n9199;
wire     [31:0] n9200;
wire     [31:0] n9201;
wire     [31:0] n9202;
wire     [31:0] n9203;
wire     [31:0] n9204;
wire     [31:0] n9205;
wire     [31:0] n9206;
wire     [31:0] n9207;
wire     [31:0] n9208;
wire     [31:0] n9209;
wire     [31:0] n9210;
wire     [31:0] n9211;
wire     [31:0] n9212;
wire     [31:0] n9213;
wire     [31:0] n9214;
wire     [31:0] n9215;
wire     [31:0] n9216;
wire     [31:0] n9217;
wire     [31:0] n9218;
wire     [31:0] n9219;
wire     [31:0] n9220;
wire     [31:0] n9221;
wire     [31:0] n9222;
wire     [31:0] n9223;
wire     [31:0] n9224;
wire     [31:0] n9225;
wire     [31:0] n9226;
wire     [31:0] n9227;
wire     [31:0] n9228;
wire     [31:0] n9229;
wire     [31:0] n9230;
wire     [31:0] n9231;
wire     [31:0] n9232;
wire     [31:0] n9233;
wire     [31:0] n9234;
wire     [31:0] n9235;
wire     [31:0] n9236;
wire     [31:0] n9237;
wire     [31:0] n9238;
wire     [31:0] n9239;
wire     [31:0] n9240;
wire     [31:0] n9241;
wire     [31:0] n9242;
wire     [31:0] n9243;
wire     [31:0] n9244;
wire     [31:0] n9245;
wire     [31:0] n9246;
wire     [31:0] n9247;
wire     [31:0] n9248;
wire     [31:0] n9249;
wire     [31:0] n9250;
wire     [31:0] n9251;
wire     [31:0] n9252;
wire     [31:0] n9253;
wire     [31:0] n9254;
wire     [31:0] n9255;
wire     [31:0] n9256;
wire     [31:0] n9257;
wire     [31:0] n9258;
wire     [31:0] n9259;
wire     [31:0] n9260;
wire     [31:0] n9261;
wire     [31:0] n9262;
wire     [31:0] n9263;
wire     [31:0] n9264;
wire     [31:0] n9265;
wire     [31:0] n9266;
wire     [31:0] n9267;
wire     [31:0] n9268;
wire     [31:0] n9269;
wire     [31:0] n9270;
wire     [31:0] n9271;
wire     [31:0] n9272;
wire     [31:0] n9273;
wire     [31:0] n9274;
wire     [31:0] n9275;
wire     [31:0] n9276;
wire     [31:0] n9277;
wire     [31:0] n9278;
wire     [31:0] n9279;
wire     [31:0] n9280;
wire     [31:0] n9281;
wire     [31:0] n9282;
wire     [31:0] n9283;
wire     [31:0] n9284;
wire     [31:0] n9285;
wire     [31:0] n9286;
wire     [31:0] n9287;
wire     [31:0] n9288;
wire     [31:0] n9289;
wire     [31:0] n9290;
wire     [31:0] n9291;
wire     [31:0] n9292;
wire     [31:0] n9293;
wire     [31:0] n9294;
wire     [31:0] n9295;
wire     [31:0] n9296;
wire     [31:0] n9297;
wire     [31:0] n9298;
wire     [31:0] n9299;
wire     [31:0] n9300;
wire     [31:0] n9301;
wire     [31:0] n9302;
wire     [31:0] n9303;
wire     [31:0] n9304;
wire     [31:0] n9305;
wire     [31:0] n9306;
wire     [31:0] n9307;
wire     [31:0] n9308;
wire     [31:0] n9309;
wire     [31:0] n9310;
wire     [31:0] n9311;
wire     [31:0] n9312;
wire     [31:0] n9313;
wire     [31:0] n9314;
wire     [31:0] n9315;
wire     [31:0] n9316;
wire     [31:0] n9317;
wire     [31:0] n9318;
wire     [31:0] n9319;
wire     [31:0] n9320;
wire     [31:0] n9321;
wire     [31:0] n9322;
wire     [31:0] n9323;
wire     [31:0] n9324;
wire     [31:0] n9325;
wire     [31:0] n9326;
wire     [31:0] n9327;
wire     [31:0] n9328;
wire     [31:0] n9329;
wire     [31:0] n9330;
wire     [31:0] n9331;
wire     [31:0] n9332;
wire     [31:0] n9333;
wire     [31:0] n9334;
wire     [31:0] n9335;
wire     [31:0] n9336;
wire     [31:0] n9337;
wire     [31:0] n9338;
wire     [31:0] n9339;
wire     [31:0] n9340;
wire     [31:0] n9341;
wire     [31:0] n9342;
wire     [31:0] n9343;
wire     [31:0] n9344;
wire     [31:0] n9345;
wire     [31:0] n9346;
wire     [31:0] n9347;
wire     [31:0] n9348;
wire     [31:0] n9349;
wire     [31:0] n9350;
wire     [31:0] n9351;
wire     [31:0] n9352;
wire     [31:0] n9353;
wire     [31:0] n9354;
wire     [31:0] n9355;
wire     [31:0] n9356;
wire     [31:0] n9357;
wire     [31:0] n9358;
wire     [31:0] n9359;
wire     [31:0] n9360;
wire     [31:0] n9361;
wire     [31:0] n9362;
wire     [31:0] n9363;
wire     [31:0] n9364;
wire     [31:0] n9365;
wire     [31:0] n9366;
wire     [31:0] n9367;
wire     [31:0] n9368;
wire     [31:0] n9369;
wire     [31:0] n9370;
wire     [31:0] n9371;
wire     [31:0] n9372;
wire     [31:0] n9373;
wire     [31:0] n9374;
wire     [31:0] n9375;
wire     [31:0] n9376;
wire     [31:0] n9377;
wire     [31:0] n9378;
wire     [31:0] n9379;
wire     [31:0] n9380;
wire     [31:0] n9381;
wire     [31:0] n9382;
wire     [31:0] n9383;
wire     [31:0] n9384;
wire     [31:0] n9385;
wire     [31:0] n9386;
wire     [31:0] n9387;
wire     [31:0] n9388;
wire     [31:0] n9389;
wire     [31:0] n9390;
wire            n9391;
wire            n9392;
wire     [31:0] n9393;
wire     [31:0] n9394;
wire     [31:0] n9395;
wire     [31:0] n9396;
wire     [31:0] n9397;
wire     [31:0] n9398;
wire     [31:0] n9399;
wire     [31:0] n9400;
wire     [31:0] n9401;
wire     [31:0] n9402;
wire     [31:0] n9403;
wire     [31:0] n9404;
wire     [31:0] n9405;
wire     [31:0] n9406;
wire     [31:0] n9407;
wire     [31:0] n9408;
wire     [31:0] n9409;
wire     [31:0] n9410;
wire     [31:0] n9411;
wire     [31:0] n9412;
wire     [31:0] n9413;
wire     [31:0] n9414;
wire     [31:0] n9415;
wire     [31:0] n9416;
wire     [31:0] n9417;
wire     [31:0] n9418;
wire     [31:0] n9419;
wire     [31:0] n9420;
wire     [31:0] n9421;
wire     [31:0] n9422;
wire     [31:0] n9423;
wire     [31:0] n9424;
wire     [31:0] n9425;
wire            n9426;
wire            n9427;
wire            n9428;
wire            n9429;
wire            n9430;
wire            n9431;
wire            n9432;
wire            n9433;
wire            n9434;
wire            n9435;
wire            n9436;
wire            n9437;
wire            n9438;
wire            n9439;
wire            n9440;
wire            n9441;
wire            n9442;
wire            n9443;
wire            n9444;
wire            n9445;
wire            n9446;
wire            n9447;
wire            n9448;
wire            n9449;
wire            n9450;
wire            n9451;
wire            n9452;
wire            n9453;
wire            n9454;
wire            n9455;
wire            n9456;
wire            n9457;
wire            n9458;
wire            n9459;
wire            n9460;
wire            n9461;
wire            n9462;
wire            n9463;
wire            n9464;
wire            n9465;
wire            n9466;
wire            n9467;
wire            n9468;
wire            n9469;
wire            n9470;
wire            n9471;
wire            n9472;
wire            n9473;
wire            n9474;
wire            n9475;
wire            n9476;
wire            n9477;
wire            n9478;
wire            n9479;
wire            n9480;
wire            n9481;
wire            n9482;
wire            n9483;
wire            n9484;
wire            n9485;
wire            n9486;
wire            n9487;
wire            n9488;
wire            n9489;
wire            n9490;
wire            n9491;
wire            n9492;
wire            n9493;
wire            n9494;
wire            n9495;
wire            n9496;
wire            n9497;
wire            n9498;
wire            n9499;
wire            n9500;
wire            n9501;
wire            n9502;
wire            n9503;
wire            n9504;
wire            n9505;
wire            n9506;
wire            n9507;
wire            n9508;
wire            n9509;
wire            n9510;
wire            n9511;
wire            n9512;
wire            n9513;
wire            n9514;
wire            n9515;
wire            n9516;
wire            n9517;
wire            n9518;
wire            n9519;
wire            n9520;
wire            n9521;
wire            n9522;
wire            n9523;
wire            n9524;
wire            n9525;
wire            n9526;
wire            n9527;
wire            n9528;
wire            n9529;
wire            n9530;
wire            n9531;
wire            n9532;
wire            n9533;
wire            n9534;
wire            n9535;
wire            n9536;
wire            n9537;
wire            n9538;
wire            n9539;
wire            n9540;
wire            n9541;
wire            n9542;
wire            n9543;
wire            n9544;
wire            n9545;
wire            n9546;
wire            n9547;
wire            n9548;
wire            n9549;
wire            n9550;
wire            n9551;
wire            n9552;
wire            n9553;
wire            n9554;
wire            n9555;
wire            n9556;
wire            n9557;
wire            n9558;
wire            n9559;
wire            n9560;
wire            n9561;
wire            n9562;
wire            n9563;
wire            n9564;
wire            n9565;
wire            n9566;
wire            n9567;
wire            n9568;
wire            n9569;
wire            n9570;
wire            n9571;
wire            n9572;
wire            n9573;
wire            n9574;
wire            n9575;
wire            n9576;
wire            n9577;
wire            n9578;
wire            n9579;
wire            n9580;
wire            n9581;
wire            n9582;
wire            n9583;
wire            n9584;
wire            n9585;
wire            n9586;
wire            n9587;
wire            n9588;
wire            n9589;
wire            n9590;
wire            n9591;
wire            n9592;
wire            n9593;
wire            n9594;
wire            n9595;
wire            n9596;
wire            n9597;
wire            n9598;
wire            n9599;
wire            n9600;
wire            n9601;
wire            n9602;
wire            n9603;
wire            n9604;
wire            n9605;
wire            n9606;
wire            n9607;
wire            n9608;
wire            n9609;
wire            n9610;
wire            n9611;
wire            n9612;
wire            n9613;
wire            n9614;
wire            n9615;
wire            n9616;
wire            n9617;
wire            n9618;
wire            n9619;
wire            n9620;
wire            n9621;
wire            n9622;
wire            n9623;
wire            n9624;
wire            n9625;
wire            n9626;
wire            n9627;
wire            n9628;
wire            n9629;
wire            n9630;
wire            n9631;
wire            n9632;
wire            n9633;
wire            n9634;
wire            n9635;
wire            n9636;
wire            n9637;
wire            n9638;
wire            n9639;
wire            n9640;
wire            n9641;
wire            n9642;
wire            n9643;
wire            n9644;
wire            n9645;
wire            n9646;
wire            n9647;
wire            n9648;
wire            n9649;
wire            n9650;
wire            n9651;
wire            n9652;
wire            n9653;
wire            n9654;
wire            n9655;
wire            n9656;
wire            n9657;
wire            n9658;
wire            n9659;
wire            n9660;
wire            n9661;
wire            n9662;
wire            n9663;
wire            n9664;
wire            n9665;
wire            n9666;
wire            n9667;
wire            n9668;
wire            n9669;
wire            n9670;
wire            n9671;
wire            n9672;
wire            n9673;
wire            n9674;
wire            n9675;
wire            n9676;
wire            n9677;
wire            n9678;
wire            n9679;
wire            n9680;
wire            n9681;
wire            n9682;
wire            n9683;
wire            n9684;
wire            n9685;
wire            n9686;
wire            n9687;
wire            n9688;
wire            n9689;
wire            n9690;
wire            n9691;
wire            n9692;
wire            n9693;
wire            n9694;
wire            n9695;
wire            n9696;
wire            n9697;
wire            n9698;
wire            n9699;
wire            n9700;
wire            n9701;
wire            n9702;
wire            n9703;
wire            n9704;
wire            n9705;
wire            n9706;
wire            n9707;
wire            n9708;
wire            n9709;
wire            n9710;
wire            n9711;
wire            n9712;
wire            n9713;
wire            n9714;
wire            n9715;
wire            n9716;
wire            n9717;
wire            n9718;
wire            n9719;
wire            n9720;
wire            n9721;
wire            n9722;
wire            n9723;
wire            n9724;
wire            n9725;
wire            n9726;
wire            n9727;
wire            n9728;
wire            n9729;
wire            n9730;
wire            n9731;
wire            n9732;
wire            n9733;
wire            n9734;
wire            n9735;
wire            n9736;
wire            n9737;
wire            n9738;
wire            n9739;
wire            n9740;
wire            n9741;
wire            n9742;
wire            n9743;
wire            n9744;
wire            n9745;
wire            n9746;
wire            n9747;
wire            n9748;
wire            n9749;
wire            n9750;
wire            n9751;
wire            n9752;
wire            n9753;
wire            n9754;
wire            n9755;
wire            n9756;
wire            n9757;
wire            n9758;
wire            n9759;
wire            n9760;
wire            n9761;
wire            n9762;
wire            n9763;
wire            n9764;
wire            n9765;
wire            n9766;
wire            n9767;
wire            n9768;
wire            n9769;
wire            n9770;
wire            n9771;
wire            n9772;
wire            n9773;
wire            n9774;
wire            n9775;
wire            n9776;
wire            n9777;
wire            n9778;
wire            n9779;
wire            n9780;
wire            n9781;
wire            n9782;
wire            n9783;
wire            n9784;
wire            n9785;
wire            n9786;
wire            n9787;
wire            n9788;
wire            n9789;
wire            n9790;
wire            n9791;
wire            n9792;
wire            n9793;
wire            n9794;
wire            n9795;
wire            n9796;
wire            n9797;
wire            n9798;
wire            n9799;
wire            n9800;
wire            n9801;
wire            n9802;
wire            n9803;
wire            n9804;
wire            n9805;
wire            n9806;
wire            n9807;
wire            n9808;
wire            n9809;
wire            n9810;
wire            n9811;
wire            n9812;
wire            n9813;
wire            n9814;
wire            n9815;
wire            n9816;
wire            n9817;
wire            n9818;
wire            n9819;
wire            n9820;
wire            n9821;
wire            n9822;
wire            n9823;
wire            n9824;
wire            n9825;
wire            n9826;
wire            n9827;
wire            n9828;
wire            n9829;
wire            n9830;
wire            n9831;
wire            n9832;
wire            n9833;
wire            n9834;
wire            n9835;
wire            n9836;
wire            n9837;
wire            n9838;
wire            n9839;
wire            n9840;
wire            n9841;
wire            n9842;
wire            n9843;
wire            n9844;
wire            n9845;
wire            n9846;
wire            n9847;
wire            n9848;
wire            n9849;
wire            n9850;
wire            n9851;
wire            n9852;
wire            n9853;
wire            n9854;
wire            n9855;
wire            n9856;
wire            n9857;
wire            n9858;
wire            n9859;
wire            n9860;
wire            n9861;
wire            n9862;
wire            n9863;
wire            n9864;
wire            n9865;
wire            n9866;
wire            n9867;
wire            n9868;
wire            n9869;
wire            n9870;
wire            n9871;
wire            n9872;
wire            n9873;
wire            n9874;
wire            n9875;
wire            n9876;
wire            n9877;
wire            n9878;
wire            n9879;
wire            n9880;
wire            n9881;
wire            n9882;
wire            n9883;
wire            n9884;
wire            n9885;
wire            n9886;
wire            n9887;
wire            n9888;
wire            n9889;
wire            n9890;
wire            n9891;
wire            n9892;
wire            n9893;
wire            n9894;
wire            n9895;
wire            n9896;
wire            n9897;
wire            n9898;
wire            n9899;
wire            n9900;
wire            n9901;
wire            n9902;
wire            n9903;
wire            n9904;
wire            n9905;
wire            n9906;
wire            n9907;
wire            n9908;
wire            n9909;
wire            n9910;
wire            n9911;
wire            n9912;
wire            n9913;
wire            n9914;
wire            n9915;
wire            n9916;
wire            n9917;
wire            n9918;
wire            n9919;
wire            n9920;
wire            n9921;
wire            n9922;
wire            n9923;
wire            n9924;
wire            n9925;
wire            n9926;
wire            n9927;
wire            n9928;
wire            n9929;
wire            n9930;
wire            n9931;
wire            n9932;
wire            n9933;
wire            n9934;
wire            n9935;
wire            n9936;
wire            n9937;
wire            n9938;
wire            n9939;
wire            n9940;
wire            n9941;
wire            n9942;
wire            n9943;
wire            n9944;
wire            n9945;
wire            n9946;
wire            n9947;
wire            n9948;
wire            n9949;
wire            n9950;
wire            n9951;
wire            n9952;
wire            n9953;
wire     [31:0] n9954;
wire     [31:0] n9955;
wire     [31:0] n9956;
wire     [31:0] n9957;
wire     [31:0] n9958;
wire     [31:0] n9959;
wire     [31:0] n9960;
wire     [31:0] n9961;
wire     [31:0] n9962;
wire     [31:0] n9963;
wire     [31:0] n9964;
wire     [31:0] n9965;
wire     [31:0] n9966;
wire     [31:0] n9967;
wire     [31:0] n9968;
wire     [31:0] n9969;
wire     [31:0] n9970;
wire     [31:0] n9971;
wire     [31:0] n9972;
wire     [31:0] n9973;
wire     [31:0] n9974;
wire     [31:0] n9975;
wire     [31:0] n9976;
wire     [31:0] n9977;
wire     [31:0] n9978;
wire     [31:0] n9979;
wire     [31:0] n9980;
wire     [31:0] n9981;
wire     [31:0] n9982;
wire     [31:0] n9983;
wire     [31:0] n9984;
wire     [31:0] n9985;
wire     [31:0] n9986;
wire     [31:0] n9987;
wire     [31:0] n9988;
wire     [31:0] n9989;
wire     [31:0] n9990;
wire     [31:0] n9991;
wire     [31:0] n9992;
wire     [31:0] n9993;
wire     [31:0] n9994;
wire     [31:0] n9995;
wire     [31:0] n9996;
wire     [31:0] n9997;
wire     [31:0] n9998;
wire     [31:0] n9999;
wire     [31:0] n10000;
wire     [31:0] n10001;
wire     [31:0] n10002;
wire     [31:0] n10003;
wire     [31:0] n10004;
wire     [31:0] n10005;
wire     [31:0] n10006;
wire     [31:0] n10007;
wire     [31:0] n10008;
wire     [31:0] n10009;
wire     [31:0] n10010;
wire     [31:0] n10011;
wire     [31:0] n10012;
wire     [31:0] n10013;
wire     [31:0] n10014;
wire     [31:0] n10015;
wire     [31:0] n10016;
wire     [31:0] n10017;
wire     [31:0] n10018;
wire     [31:0] n10019;
wire     [31:0] n10020;
wire     [31:0] n10021;
wire     [31:0] n10022;
wire     [31:0] n10023;
wire     [31:0] n10024;
wire     [31:0] n10025;
wire     [31:0] n10026;
wire     [31:0] n10027;
wire     [31:0] n10028;
wire     [31:0] n10029;
wire     [31:0] n10030;
wire     [31:0] n10031;
wire     [31:0] n10032;
wire     [31:0] n10033;
wire     [31:0] n10034;
wire     [31:0] n10035;
wire     [31:0] n10036;
wire     [31:0] n10037;
wire     [31:0] n10038;
wire     [31:0] n10039;
wire     [31:0] n10040;
wire     [31:0] n10041;
wire     [31:0] n10042;
wire     [31:0] n10043;
wire     [31:0] n10044;
wire     [31:0] n10045;
wire     [31:0] n10046;
wire     [31:0] n10047;
wire     [31:0] n10048;
wire     [31:0] n10049;
wire     [31:0] n10050;
wire     [31:0] n10051;
wire     [31:0] n10052;
wire     [31:0] n10053;
wire     [31:0] n10054;
wire     [31:0] n10055;
wire     [31:0] n10056;
wire     [31:0] n10057;
wire     [31:0] n10058;
wire     [31:0] n10059;
wire     [31:0] n10060;
wire     [31:0] n10061;
wire     [31:0] n10062;
wire     [31:0] n10063;
wire     [31:0] n10064;
wire     [31:0] n10065;
wire     [31:0] n10066;
wire     [31:0] n10067;
wire     [31:0] n10068;
wire     [31:0] n10069;
wire     [31:0] n10070;
wire     [31:0] n10071;
wire     [31:0] n10072;
wire     [31:0] n10073;
wire     [31:0] n10074;
wire     [31:0] n10075;
wire     [31:0] n10076;
wire     [31:0] n10077;
wire     [31:0] n10078;
wire     [31:0] n10079;
wire     [31:0] n10080;
wire     [31:0] n10081;
wire     [31:0] n10082;
wire     [31:0] n10083;
wire     [31:0] n10084;
wire     [31:0] n10085;
wire     [31:0] n10086;
wire     [31:0] n10087;
wire     [31:0] n10088;
wire     [31:0] n10089;
wire     [31:0] n10090;
wire     [31:0] n10091;
wire     [31:0] n10092;
wire     [31:0] n10093;
wire     [31:0] n10094;
wire     [31:0] n10095;
wire     [31:0] n10096;
wire     [31:0] n10097;
wire     [31:0] n10098;
wire     [31:0] n10099;
wire     [31:0] n10100;
wire     [31:0] n10101;
wire     [31:0] n10102;
wire     [31:0] n10103;
wire     [31:0] n10104;
wire     [31:0] n10105;
wire     [31:0] n10106;
wire     [31:0] n10107;
wire     [31:0] n10108;
wire     [31:0] n10109;
wire     [31:0] n10110;
wire     [31:0] n10111;
wire     [31:0] n10112;
wire     [31:0] n10113;
wire     [31:0] n10114;
wire     [31:0] n10115;
wire     [31:0] n10116;
wire     [31:0] n10117;
wire     [31:0] n10118;
wire     [31:0] n10119;
wire     [31:0] n10120;
wire     [31:0] n10121;
wire     [31:0] n10122;
wire     [31:0] n10123;
wire     [31:0] n10124;
wire     [31:0] n10125;
wire     [31:0] n10126;
wire     [31:0] n10127;
wire     [31:0] n10128;
wire     [31:0] n10129;
wire     [31:0] n10130;
wire     [31:0] n10131;
wire     [31:0] n10132;
wire     [31:0] n10133;
wire     [31:0] n10134;
wire     [31:0] n10135;
wire     [31:0] n10136;
wire     [31:0] n10137;
wire     [31:0] n10138;
wire     [31:0] n10139;
wire     [31:0] n10140;
wire     [31:0] n10141;
wire     [31:0] n10142;
wire     [31:0] n10143;
wire     [31:0] n10144;
wire     [31:0] n10145;
wire     [31:0] n10146;
wire     [31:0] n10147;
wire     [31:0] n10148;
wire     [31:0] n10149;
wire     [31:0] n10150;
wire     [31:0] n10151;
wire     [31:0] n10152;
wire     [31:0] n10153;
wire     [31:0] n10154;
wire     [31:0] n10155;
wire     [31:0] n10156;
wire     [31:0] n10157;
wire     [31:0] n10158;
wire     [31:0] n10159;
wire     [31:0] n10160;
wire     [31:0] n10161;
wire     [31:0] n10162;
wire     [31:0] n10163;
wire     [31:0] n10164;
wire     [31:0] n10165;
wire     [31:0] n10166;
wire     [31:0] n10167;
wire     [31:0] n10168;
wire     [31:0] n10169;
wire     [31:0] n10170;
wire     [31:0] n10171;
wire     [31:0] n10172;
wire     [31:0] n10173;
wire     [31:0] n10174;
wire     [31:0] n10175;
wire     [31:0] n10176;
wire     [31:0] n10177;
wire     [31:0] n10178;
wire     [31:0] n10179;
wire     [31:0] n10180;
wire     [31:0] n10181;
wire     [31:0] n10182;
wire     [31:0] n10183;
wire     [31:0] n10184;
wire     [31:0] n10185;
wire     [31:0] n10186;
wire     [31:0] n10187;
wire     [31:0] n10188;
wire     [31:0] n10189;
wire     [31:0] n10190;
wire     [31:0] n10191;
wire     [31:0] n10192;
wire     [31:0] n10193;
wire     [31:0] n10194;
wire     [31:0] n10195;
wire     [31:0] n10196;
wire     [31:0] n10197;
wire     [31:0] n10198;
wire     [31:0] n10199;
wire     [31:0] n10200;
wire     [31:0] n10201;
wire     [31:0] n10202;
wire     [31:0] n10203;
wire     [31:0] n10204;
wire     [31:0] n10205;
wire     [31:0] n10206;
wire     [31:0] n10207;
wire     [31:0] n10208;
wire     [31:0] n10209;
wire     [31:0] n10210;
wire     [31:0] n10211;
wire     [31:0] n10212;
wire     [31:0] n10213;
wire     [31:0] n10214;
wire     [31:0] n10215;
wire     [31:0] n10216;
wire     [31:0] n10217;
wire     [31:0] n10218;
wire     [31:0] n10219;
wire     [31:0] n10220;
wire     [31:0] n10221;
wire     [31:0] n10222;
wire     [31:0] n10223;
wire     [31:0] n10224;
wire     [31:0] n10225;
wire     [31:0] n10226;
wire     [31:0] n10227;
wire     [31:0] n10228;
wire     [31:0] n10229;
wire     [31:0] n10230;
wire     [31:0] n10231;
wire     [31:0] n10232;
wire     [31:0] n10233;
wire     [31:0] n10234;
wire     [31:0] n10235;
wire     [31:0] n10236;
wire     [31:0] n10237;
wire     [31:0] n10238;
wire     [31:0] n10239;
wire     [31:0] n10240;
wire     [31:0] n10241;
wire     [31:0] n10242;
wire     [31:0] n10243;
wire     [31:0] n10244;
wire     [31:0] n10245;
wire     [31:0] n10246;
wire     [31:0] n10247;
wire     [31:0] n10248;
wire     [31:0] n10249;
wire     [31:0] n10250;
wire     [31:0] n10251;
wire     [31:0] n10252;
wire     [31:0] n10253;
wire     [31:0] n10254;
wire     [31:0] n10255;
wire     [31:0] n10256;
wire     [31:0] n10257;
wire     [31:0] n10258;
wire     [31:0] n10259;
wire     [31:0] n10260;
wire     [31:0] n10261;
wire     [31:0] n10262;
wire     [31:0] n10263;
wire     [31:0] n10264;
wire     [31:0] n10265;
wire     [31:0] n10266;
wire     [31:0] n10267;
wire     [31:0] n10268;
wire     [31:0] n10269;
wire     [31:0] n10270;
wire     [31:0] n10271;
wire     [31:0] n10272;
wire     [31:0] n10273;
wire     [31:0] n10274;
wire     [31:0] n10275;
wire     [31:0] n10276;
wire     [31:0] n10277;
wire     [31:0] n10278;
wire     [31:0] n10279;
wire     [31:0] n10280;
wire     [31:0] n10281;
wire     [31:0] n10282;
wire     [31:0] n10283;
wire     [31:0] n10284;
wire     [31:0] n10285;
wire     [31:0] n10286;
wire     [31:0] n10287;
wire     [31:0] n10288;
wire     [31:0] n10289;
wire     [31:0] n10290;
wire     [31:0] n10291;
wire     [31:0] n10292;
wire     [31:0] n10293;
wire     [31:0] n10294;
wire     [31:0] n10295;
wire     [31:0] n10296;
wire     [31:0] n10297;
wire     [31:0] n10298;
wire     [31:0] n10299;
wire     [31:0] n10300;
wire     [31:0] n10301;
wire     [31:0] n10302;
wire     [31:0] n10303;
wire     [31:0] n10304;
wire     [31:0] n10305;
wire     [31:0] n10306;
wire     [31:0] n10307;
wire     [31:0] n10308;
wire     [31:0] n10309;
wire     [31:0] n10310;
wire     [31:0] n10311;
wire     [31:0] n10312;
wire     [31:0] n10313;
wire     [31:0] n10314;
wire     [31:0] n10315;
wire     [31:0] n10316;
wire     [31:0] n10317;
wire     [31:0] n10318;
wire     [31:0] n10319;
wire     [31:0] n10320;
wire     [31:0] n10321;
wire     [31:0] n10322;
wire     [31:0] n10323;
wire     [31:0] n10324;
wire     [31:0] n10325;
wire     [31:0] n10326;
wire     [31:0] n10327;
wire     [31:0] n10328;
wire     [31:0] n10329;
wire     [31:0] n10330;
wire     [31:0] n10331;
wire     [31:0] n10332;
wire     [31:0] n10333;
wire     [31:0] n10334;
wire     [31:0] n10335;
wire     [31:0] n10336;
wire     [31:0] n10337;
wire     [31:0] n10338;
wire     [31:0] n10339;
wire     [31:0] n10340;
wire     [31:0] n10341;
wire     [31:0] n10342;
wire     [31:0] n10343;
wire     [31:0] n10344;
wire     [31:0] n10345;
wire     [31:0] n10346;
wire     [31:0] n10347;
wire     [31:0] n10348;
wire     [31:0] n10349;
wire     [31:0] n10350;
wire     [31:0] n10351;
wire     [31:0] n10352;
wire     [31:0] n10353;
wire     [31:0] n10354;
wire     [31:0] n10355;
wire     [31:0] n10356;
wire     [31:0] n10357;
wire     [31:0] n10358;
wire     [31:0] n10359;
wire     [31:0] n10360;
wire     [31:0] n10361;
wire     [31:0] n10362;
wire     [31:0] n10363;
wire     [31:0] n10364;
wire     [31:0] n10365;
wire     [31:0] n10366;
wire     [31:0] n10367;
wire     [31:0] n10368;
wire     [31:0] n10369;
wire     [31:0] n10370;
wire     [31:0] n10371;
wire     [31:0] n10372;
wire     [31:0] n10373;
wire     [31:0] n10374;
wire     [31:0] n10375;
wire     [31:0] n10376;
wire     [31:0] n10377;
wire     [31:0] n10378;
wire     [31:0] n10379;
wire     [31:0] n10380;
wire     [31:0] n10381;
wire     [31:0] n10382;
wire     [31:0] n10383;
wire     [31:0] n10384;
wire     [31:0] n10385;
wire     [31:0] n10386;
wire     [31:0] n10387;
wire     [31:0] n10388;
wire     [31:0] n10389;
wire     [31:0] n10390;
wire     [31:0] n10391;
wire     [31:0] n10392;
wire     [31:0] n10393;
wire     [31:0] n10394;
wire     [31:0] n10395;
wire     [31:0] n10396;
wire     [31:0] n10397;
wire     [31:0] n10398;
wire     [31:0] n10399;
wire     [31:0] n10400;
wire     [31:0] n10401;
wire     [31:0] n10402;
wire     [31:0] n10403;
wire     [31:0] n10404;
wire     [31:0] n10405;
wire     [31:0] n10406;
wire     [31:0] n10407;
wire     [31:0] n10408;
wire     [31:0] n10409;
wire     [31:0] n10410;
wire     [31:0] n10411;
wire     [31:0] n10412;
wire     [31:0] n10413;
wire     [31:0] n10414;
wire     [31:0] n10415;
wire     [31:0] n10416;
wire     [31:0] n10417;
wire     [31:0] n10418;
wire     [31:0] n10419;
wire     [31:0] n10420;
wire     [31:0] n10421;
wire     [31:0] n10422;
wire     [31:0] n10423;
wire     [31:0] n10424;
wire     [31:0] n10425;
wire     [31:0] n10426;
wire     [31:0] n10427;
wire     [31:0] n10428;
wire     [31:0] n10429;
wire     [31:0] n10430;
wire     [31:0] n10431;
wire     [31:0] n10432;
wire     [31:0] n10433;
wire     [31:0] n10434;
wire     [31:0] n10435;
wire     [31:0] n10436;
wire     [31:0] n10437;
wire     [31:0] n10438;
wire     [31:0] n10439;
wire     [31:0] n10440;
wire     [31:0] n10441;
wire     [31:0] n10442;
wire     [31:0] n10443;
wire     [31:0] n10444;
wire     [31:0] n10445;
wire     [31:0] n10446;
wire     [31:0] n10447;
wire     [31:0] n10448;
wire     [31:0] n10449;
wire     [31:0] n10450;
wire     [31:0] n10451;
wire     [31:0] n10452;
wire     [31:0] n10453;
wire     [31:0] n10454;
wire     [31:0] n10455;
wire     [31:0] n10456;
wire     [31:0] n10457;
wire     [31:0] n10458;
wire     [31:0] n10459;
wire     [31:0] n10460;
wire     [31:0] n10461;
wire     [31:0] n10462;
wire     [31:0] n10463;
wire     [31:0] n10464;
wire     [31:0] n10465;
wire     [31:0] n10466;
wire     [31:0] n10467;
wire     [31:0] n10468;
wire     [31:0] n10469;
wire     [31:0] n10470;
wire     [31:0] n10471;
wire     [31:0] n10472;
wire     [31:0] n10473;
wire     [31:0] n10474;
wire     [31:0] n10475;
wire            n10476;
wire            n10477;
wire            n10478;
wire            n10479;
wire            n10480;
wire            n10481;
wire            n10482;
wire            n10483;
wire            n10484;
wire            n10485;
wire            n10486;
wire            n10487;
wire            n10488;
wire            n10489;
wire            n10490;
wire            n10491;
wire            n10492;
wire            n10493;
wire            n10494;
wire            n10495;
wire            n10496;
wire            n10497;
wire            n10498;
wire            n10499;
wire            n10500;
wire            n10501;
wire            n10502;
wire            n10503;
wire            n10504;
wire            n10505;
wire            n10506;
wire            n10507;
wire            n10508;
wire            n10509;
wire            n10510;
wire            n10511;
wire            n10512;
wire            n10513;
wire            n10514;
wire            n10515;
wire            n10516;
wire            n10517;
wire            n10518;
wire            n10519;
wire            n10520;
wire            n10521;
wire            n10522;
wire            n10523;
wire            n10524;
wire            n10525;
wire            n10526;
wire            n10527;
wire            n10528;
wire            n10529;
wire            n10530;
wire            n10531;
wire            n10532;
wire            n10533;
wire            n10534;
wire            n10535;
wire            n10536;
wire            n10537;
wire            n10538;
wire            n10539;
wire            n10540;
wire            n10541;
wire            n10542;
wire            n10543;
wire            n10544;
wire            n10545;
wire            n10546;
wire            n10547;
wire            n10548;
wire            n10549;
wire            n10550;
wire            n10551;
wire            n10552;
wire            n10553;
wire            n10554;
wire            n10555;
wire            n10556;
wire            n10557;
wire            n10558;
wire            n10559;
wire            n10560;
wire            n10561;
wire            n10562;
wire            n10563;
wire            n10564;
wire            n10565;
wire            n10566;
wire            n10567;
wire            n10568;
wire            n10569;
wire            n10570;
wire            n10571;
wire            n10572;
wire            n10573;
wire            n10574;
wire            n10575;
wire            n10576;
wire            n10577;
wire            n10578;
wire            n10579;
wire            n10580;
wire            n10581;
wire            n10582;
wire            n10583;
wire            n10584;
wire            n10585;
wire            n10586;
wire            n10587;
wire            n10588;
wire            n10589;
wire            n10590;
wire            n10591;
wire            n10592;
wire            n10593;
wire            n10594;
wire            n10595;
wire            n10596;
wire            n10597;
wire            n10598;
wire            n10599;
wire            n10600;
wire            n10601;
wire            n10602;
wire            n10603;
wire            n10604;
wire            n10605;
wire            n10606;
wire            n10607;
wire            n10608;
wire            n10609;
wire            n10610;
wire            n10611;
wire            n10612;
wire            n10613;
wire            n10614;
wire            n10615;
wire            n10616;
wire            n10617;
wire            n10618;
wire            n10619;
wire            n10620;
wire            n10621;
wire            n10622;
wire            n10623;
wire            n10624;
wire            n10625;
wire            n10626;
wire            n10627;
wire            n10628;
wire            n10629;
wire            n10630;
wire            n10631;
wire            n10632;
wire            n10633;
wire            n10634;
wire            n10635;
wire            n10636;
wire            n10637;
wire            n10638;
wire            n10639;
wire            n10640;
wire            n10641;
wire            n10642;
wire            n10643;
wire            n10644;
wire            n10645;
wire            n10646;
wire            n10647;
wire            n10648;
wire            n10649;
wire            n10650;
wire            n10651;
wire            n10652;
wire            n10653;
wire            n10654;
wire            n10655;
wire            n10656;
wire            n10657;
wire            n10658;
wire            n10659;
wire            n10660;
wire            n10661;
wire            n10662;
wire            n10663;
wire            n10664;
wire            n10665;
wire            n10666;
wire            n10667;
wire            n10668;
wire            n10669;
wire            n10670;
wire            n10671;
wire            n10672;
wire            n10673;
wire            n10674;
wire            n10675;
wire            n10676;
wire            n10677;
wire            n10678;
wire            n10679;
wire            n10680;
wire            n10681;
wire            n10682;
wire            n10683;
wire            n10684;
wire            n10685;
wire            n10686;
wire            n10687;
wire            n10688;
wire            n10689;
wire            n10690;
wire            n10691;
wire            n10692;
wire            n10693;
wire            n10694;
wire            n10695;
wire            n10696;
wire            n10697;
wire            n10698;
wire            n10699;
wire            n10700;
wire            n10701;
wire            n10702;
wire            n10703;
wire            n10704;
wire            n10705;
wire            n10706;
wire            n10707;
wire            n10708;
wire            n10709;
wire            n10710;
wire            n10711;
wire            n10712;
wire            n10713;
wire            n10714;
wire            n10715;
wire            n10716;
wire            n10717;
wire            n10718;
wire            n10719;
wire            n10720;
wire            n10721;
wire            n10722;
wire            n10723;
wire            n10724;
wire            n10725;
wire            n10726;
wire            n10727;
wire            n10728;
wire            n10729;
wire            n10730;
wire            n10731;
wire            n10732;
wire            n10733;
wire            n10734;
wire            n10735;
wire            n10736;
wire            n10737;
wire            n10738;
wire            n10739;
wire            n10740;
wire            n10741;
wire            n10742;
wire            n10743;
wire            n10744;
wire            n10745;
wire            n10746;
wire            n10747;
wire            n10748;
wire            n10749;
wire            n10750;
wire            n10751;
wire            n10752;
wire            n10753;
wire            n10754;
wire            n10755;
wire            n10756;
wire            n10757;
wire            n10758;
wire            n10759;
wire            n10760;
wire            n10761;
wire            n10762;
wire            n10763;
wire            n10764;
wire            n10765;
wire            n10766;
wire            n10767;
wire            n10768;
wire            n10769;
wire            n10770;
wire            n10771;
wire            n10772;
wire            n10773;
wire            n10774;
wire            n10775;
wire            n10776;
wire            n10777;
wire            n10778;
wire            n10779;
wire            n10780;
wire            n10781;
wire            n10782;
wire            n10783;
wire            n10784;
wire            n10785;
wire            n10786;
wire            n10787;
wire            n10788;
wire            n10789;
wire            n10790;
wire            n10791;
wire            n10792;
wire            n10793;
wire            n10794;
wire            n10795;
wire            n10796;
wire            n10797;
wire            n10798;
wire            n10799;
wire            n10800;
wire            n10801;
wire            n10802;
wire            n10803;
wire            n10804;
wire            n10805;
wire            n10806;
wire            n10807;
wire            n10808;
wire            n10809;
wire            n10810;
wire            n10811;
wire            n10812;
wire            n10813;
wire            n10814;
wire            n10815;
wire            n10816;
wire            n10817;
wire            n10818;
wire            n10819;
wire            n10820;
wire            n10821;
wire            n10822;
wire            n10823;
wire            n10824;
wire            n10825;
wire            n10826;
wire            n10827;
wire            n10828;
wire            n10829;
wire            n10830;
wire            n10831;
wire            n10832;
wire            n10833;
wire            n10834;
wire            n10835;
wire            n10836;
wire            n10837;
wire            n10838;
wire            n10839;
wire            n10840;
wire            n10841;
wire            n10842;
wire            n10843;
wire            n10844;
wire            n10845;
wire            n10846;
wire            n10847;
wire            n10848;
wire            n10849;
wire            n10850;
wire            n10851;
wire            n10852;
wire            n10853;
wire            n10854;
wire            n10855;
wire            n10856;
wire            n10857;
wire            n10858;
wire            n10859;
wire            n10860;
wire            n10861;
wire            n10862;
wire            n10863;
wire            n10864;
wire            n10865;
wire            n10866;
wire            n10867;
wire            n10868;
wire            n10869;
wire            n10870;
wire            n10871;
wire            n10872;
wire            n10873;
wire            n10874;
wire            n10875;
wire            n10876;
wire            n10877;
wire            n10878;
wire            n10879;
wire            n10880;
wire            n10881;
wire            n10882;
wire            n10883;
wire            n10884;
wire            n10885;
wire            n10886;
wire            n10887;
wire            n10888;
wire            n10889;
wire            n10890;
wire            n10891;
wire            n10892;
wire            n10893;
wire            n10894;
wire            n10895;
wire            n10896;
wire            n10897;
wire            n10898;
wire            n10899;
wire            n10900;
wire            n10901;
wire            n10902;
wire            n10903;
wire            n10904;
wire            n10905;
wire            n10906;
wire            n10907;
wire            n10908;
wire            n10909;
wire            n10910;
wire            n10911;
wire            n10912;
wire            n10913;
wire            n10914;
wire            n10915;
wire            n10916;
wire            n10917;
wire            n10918;
wire            n10919;
wire            n10920;
wire            n10921;
wire            n10922;
wire            n10923;
wire            n10924;
wire            n10925;
wire            n10926;
wire            n10927;
wire            n10928;
wire            n10929;
wire            n10930;
wire            n10931;
wire            n10932;
wire            n10933;
wire            n10934;
wire            n10935;
wire            n10936;
wire            n10937;
wire            n10938;
wire            n10939;
wire            n10940;
wire            n10941;
wire            n10942;
wire            n10943;
wire            n10944;
wire            n10945;
wire            n10946;
wire            n10947;
wire            n10948;
wire            n10949;
wire            n10950;
wire            n10951;
wire            n10952;
wire            n10953;
wire            n10954;
wire            n10955;
wire            n10956;
wire            n10957;
wire            n10958;
wire            n10959;
wire            n10960;
wire            n10961;
wire            n10962;
wire            n10963;
wire            n10964;
wire            n10965;
wire            n10966;
wire            n10967;
wire            n10968;
wire            n10969;
wire            n10970;
wire            n10971;
wire            n10972;
wire            n10973;
wire            n10974;
wire            n10975;
wire            n10976;
wire            n10977;
wire            n10978;
wire            n10979;
wire            n10980;
wire            n10981;
wire            n10982;
wire            n10983;
wire            n10984;
wire            n10985;
wire            n10986;
wire            n10987;
wire     [31:0] n10988;
wire     [31:0] n10989;
wire     [31:0] n10990;
wire     [31:0] n10991;
wire     [31:0] n10992;
wire     [31:0] n10993;
wire     [31:0] n10994;
wire     [31:0] n10995;
wire     [31:0] n10996;
wire     [31:0] n10997;
wire     [31:0] n10998;
wire     [31:0] n10999;
wire     [31:0] n11000;
wire     [31:0] n11001;
wire     [31:0] n11002;
wire     [31:0] n11003;
wire     [31:0] n11004;
wire     [31:0] n11005;
wire     [31:0] n11006;
wire     [31:0] n11007;
wire     [31:0] n11008;
wire     [31:0] n11009;
wire     [31:0] n11010;
wire     [31:0] n11011;
wire     [31:0] n11012;
wire     [31:0] n11013;
wire     [31:0] n11014;
wire     [31:0] n11015;
wire     [31:0] n11016;
wire     [31:0] n11017;
wire     [31:0] n11018;
wire     [31:0] n11019;
wire     [31:0] n11020;
wire     [31:0] n11021;
wire     [31:0] n11022;
wire     [31:0] n11023;
wire     [31:0] n11024;
wire     [31:0] n11025;
wire     [31:0] n11026;
wire     [31:0] n11027;
wire     [31:0] n11028;
wire     [31:0] n11029;
wire     [31:0] n11030;
wire     [31:0] n11031;
wire     [31:0] n11032;
wire     [31:0] n11033;
wire     [31:0] n11034;
wire     [31:0] n11035;
wire     [31:0] n11036;
wire     [31:0] n11037;
wire     [31:0] n11038;
wire     [31:0] n11039;
wire     [31:0] n11040;
wire     [31:0] n11041;
wire     [31:0] n11042;
wire     [31:0] n11043;
wire     [31:0] n11044;
wire     [31:0] n11045;
wire     [31:0] n11046;
wire     [31:0] n11047;
wire     [31:0] n11048;
wire     [31:0] n11049;
wire     [31:0] n11050;
wire     [31:0] n11051;
wire     [31:0] n11052;
wire     [31:0] n11053;
wire     [31:0] n11054;
wire     [31:0] n11055;
wire     [31:0] n11056;
wire     [31:0] n11057;
wire     [31:0] n11058;
wire     [31:0] n11059;
wire     [31:0] n11060;
wire     [31:0] n11061;
wire     [31:0] n11062;
wire     [31:0] n11063;
wire     [31:0] n11064;
wire     [31:0] n11065;
wire     [31:0] n11066;
wire     [31:0] n11067;
wire     [31:0] n11068;
wire     [31:0] n11069;
wire     [31:0] n11070;
wire     [31:0] n11071;
wire     [31:0] n11072;
wire     [31:0] n11073;
wire     [31:0] n11074;
wire     [31:0] n11075;
wire     [31:0] n11076;
wire     [31:0] n11077;
wire     [31:0] n11078;
wire     [31:0] n11079;
wire     [31:0] n11080;
wire     [31:0] n11081;
wire     [31:0] n11082;
wire     [31:0] n11083;
wire     [31:0] n11084;
wire     [31:0] n11085;
wire     [31:0] n11086;
wire     [31:0] n11087;
wire     [31:0] n11088;
wire     [31:0] n11089;
wire     [31:0] n11090;
wire     [31:0] n11091;
wire     [31:0] n11092;
wire     [31:0] n11093;
wire     [31:0] n11094;
wire     [31:0] n11095;
wire     [31:0] n11096;
wire     [31:0] n11097;
wire     [31:0] n11098;
wire     [31:0] n11099;
wire     [31:0] n11100;
wire     [31:0] n11101;
wire     [31:0] n11102;
wire     [31:0] n11103;
wire     [31:0] n11104;
wire     [31:0] n11105;
wire     [31:0] n11106;
wire     [31:0] n11107;
wire     [31:0] n11108;
wire     [31:0] n11109;
wire     [31:0] n11110;
wire     [31:0] n11111;
wire     [31:0] n11112;
wire     [31:0] n11113;
wire     [31:0] n11114;
wire     [31:0] n11115;
wire     [31:0] n11116;
wire     [31:0] n11117;
wire     [31:0] n11118;
wire     [31:0] n11119;
wire     [31:0] n11120;
wire     [31:0] n11121;
wire     [31:0] n11122;
wire     [31:0] n11123;
wire     [31:0] n11124;
wire     [31:0] n11125;
wire     [31:0] n11126;
wire     [31:0] n11127;
wire     [31:0] n11128;
wire     [31:0] n11129;
wire     [31:0] n11130;
wire     [31:0] n11131;
wire     [31:0] n11132;
wire     [31:0] n11133;
wire     [31:0] n11134;
wire     [31:0] n11135;
wire     [31:0] n11136;
wire     [31:0] n11137;
wire     [31:0] n11138;
wire     [31:0] n11139;
wire     [31:0] n11140;
wire     [31:0] n11141;
wire     [31:0] n11142;
wire     [31:0] n11143;
wire     [31:0] n11144;
wire     [31:0] n11145;
wire     [31:0] n11146;
wire     [31:0] n11147;
wire     [31:0] n11148;
wire     [31:0] n11149;
wire     [31:0] n11150;
wire     [31:0] n11151;
wire     [31:0] n11152;
wire     [31:0] n11153;
wire     [31:0] n11154;
wire     [31:0] n11155;
wire     [31:0] n11156;
wire     [31:0] n11157;
wire     [31:0] n11158;
wire     [31:0] n11159;
wire     [31:0] n11160;
wire     [31:0] n11161;
wire     [31:0] n11162;
wire     [31:0] n11163;
wire     [31:0] n11164;
wire     [31:0] n11165;
wire     [31:0] n11166;
wire     [31:0] n11167;
wire     [31:0] n11168;
wire     [31:0] n11169;
wire     [31:0] n11170;
wire     [31:0] n11171;
wire     [31:0] n11172;
wire     [31:0] n11173;
wire     [31:0] n11174;
wire     [31:0] n11175;
wire     [31:0] n11176;
wire     [31:0] n11177;
wire     [31:0] n11178;
wire     [31:0] n11179;
wire     [31:0] n11180;
wire     [31:0] n11181;
wire     [31:0] n11182;
wire     [31:0] n11183;
wire     [31:0] n11184;
wire     [31:0] n11185;
wire     [31:0] n11186;
wire     [31:0] n11187;
wire     [31:0] n11188;
wire     [31:0] n11189;
wire     [31:0] n11190;
wire     [31:0] n11191;
wire     [31:0] n11192;
wire     [31:0] n11193;
wire     [31:0] n11194;
wire     [31:0] n11195;
wire     [31:0] n11196;
wire     [31:0] n11197;
wire     [31:0] n11198;
wire     [31:0] n11199;
wire     [31:0] n11200;
wire     [31:0] n11201;
wire     [31:0] n11202;
wire     [31:0] n11203;
wire     [31:0] n11204;
wire     [31:0] n11205;
wire     [31:0] n11206;
wire     [31:0] n11207;
wire     [31:0] n11208;
wire     [31:0] n11209;
wire     [31:0] n11210;
wire     [31:0] n11211;
wire     [31:0] n11212;
wire     [31:0] n11213;
wire     [31:0] n11214;
wire     [31:0] n11215;
wire     [31:0] n11216;
wire     [31:0] n11217;
wire     [31:0] n11218;
wire     [31:0] n11219;
wire     [31:0] n11220;
wire     [31:0] n11221;
wire     [31:0] n11222;
wire     [31:0] n11223;
wire     [31:0] n11224;
wire     [31:0] n11225;
wire     [31:0] n11226;
wire     [31:0] n11227;
wire     [31:0] n11228;
wire     [31:0] n11229;
wire     [31:0] n11230;
wire     [31:0] n11231;
wire     [31:0] n11232;
wire     [31:0] n11233;
wire     [31:0] n11234;
wire     [31:0] n11235;
wire     [31:0] n11236;
wire     [31:0] n11237;
wire     [31:0] n11238;
wire     [31:0] n11239;
wire     [31:0] n11240;
wire     [31:0] n11241;
wire     [31:0] n11242;
wire     [31:0] n11243;
wire     [31:0] n11244;
wire     [31:0] n11245;
wire     [31:0] n11246;
wire     [31:0] n11247;
wire     [31:0] n11248;
wire     [31:0] n11249;
wire     [31:0] n11250;
wire     [31:0] n11251;
wire     [31:0] n11252;
wire     [31:0] n11253;
wire     [31:0] n11254;
wire     [31:0] n11255;
wire     [31:0] n11256;
wire     [31:0] n11257;
wire     [31:0] n11258;
wire     [31:0] n11259;
wire     [31:0] n11260;
wire     [31:0] n11261;
wire     [31:0] n11262;
wire     [31:0] n11263;
wire     [31:0] n11264;
wire     [31:0] n11265;
wire     [31:0] n11266;
wire     [31:0] n11267;
wire     [31:0] n11268;
wire     [31:0] n11269;
wire     [31:0] n11270;
wire     [31:0] n11271;
wire     [31:0] n11272;
wire     [31:0] n11273;
wire     [31:0] n11274;
wire     [31:0] n11275;
wire     [31:0] n11276;
wire     [31:0] n11277;
wire     [31:0] n11278;
wire     [31:0] n11279;
wire     [31:0] n11280;
wire     [31:0] n11281;
wire     [31:0] n11282;
wire     [31:0] n11283;
wire     [31:0] n11284;
wire     [31:0] n11285;
wire     [31:0] n11286;
wire     [31:0] n11287;
wire     [31:0] n11288;
wire     [31:0] n11289;
wire     [31:0] n11290;
wire     [31:0] n11291;
wire     [31:0] n11292;
wire     [31:0] n11293;
wire     [31:0] n11294;
wire     [31:0] n11295;
wire     [31:0] n11296;
wire     [31:0] n11297;
wire     [31:0] n11298;
wire     [31:0] n11299;
wire     [31:0] n11300;
wire     [31:0] n11301;
wire     [31:0] n11302;
wire     [31:0] n11303;
wire     [31:0] n11304;
wire     [31:0] n11305;
wire     [31:0] n11306;
wire     [31:0] n11307;
wire     [31:0] n11308;
wire     [31:0] n11309;
wire     [31:0] n11310;
wire     [31:0] n11311;
wire     [31:0] n11312;
wire     [31:0] n11313;
wire     [31:0] n11314;
wire     [31:0] n11315;
wire     [31:0] n11316;
wire     [31:0] n11317;
wire     [31:0] n11318;
wire     [31:0] n11319;
wire     [31:0] n11320;
wire     [31:0] n11321;
wire     [31:0] n11322;
wire     [31:0] n11323;
wire     [31:0] n11324;
wire     [31:0] n11325;
wire     [31:0] n11326;
wire     [31:0] n11327;
wire     [31:0] n11328;
wire     [31:0] n11329;
wire     [31:0] n11330;
wire     [31:0] n11331;
wire     [31:0] n11332;
wire     [31:0] n11333;
wire     [31:0] n11334;
wire     [31:0] n11335;
wire     [31:0] n11336;
wire     [31:0] n11337;
wire     [31:0] n11338;
wire     [31:0] n11339;
wire     [31:0] n11340;
wire     [31:0] n11341;
wire     [31:0] n11342;
wire     [31:0] n11343;
wire     [31:0] n11344;
wire     [31:0] n11345;
wire     [31:0] n11346;
wire     [31:0] n11347;
wire     [31:0] n11348;
wire     [31:0] n11349;
wire     [31:0] n11350;
wire     [31:0] n11351;
wire     [31:0] n11352;
wire     [31:0] n11353;
wire     [31:0] n11354;
wire     [31:0] n11355;
wire     [31:0] n11356;
wire     [31:0] n11357;
wire     [31:0] n11358;
wire     [31:0] n11359;
wire     [31:0] n11360;
wire     [31:0] n11361;
wire     [31:0] n11362;
wire     [31:0] n11363;
wire     [31:0] n11364;
wire     [31:0] n11365;
wire     [31:0] n11366;
wire     [31:0] n11367;
wire     [31:0] n11368;
wire     [31:0] n11369;
wire     [31:0] n11370;
wire     [31:0] n11371;
wire     [31:0] n11372;
wire     [31:0] n11373;
wire     [31:0] n11374;
wire     [31:0] n11375;
wire     [31:0] n11376;
wire     [31:0] n11377;
wire     [31:0] n11378;
wire     [31:0] n11379;
wire     [31:0] n11380;
wire     [31:0] n11381;
wire     [31:0] n11382;
wire     [31:0] n11383;
wire     [31:0] n11384;
wire     [31:0] n11385;
wire     [31:0] n11386;
wire     [31:0] n11387;
wire     [31:0] n11388;
wire     [31:0] n11389;
wire     [31:0] n11390;
wire     [31:0] n11391;
wire     [31:0] n11392;
wire     [31:0] n11393;
wire     [31:0] n11394;
wire     [31:0] n11395;
wire     [31:0] n11396;
wire     [31:0] n11397;
wire     [31:0] n11398;
wire     [31:0] n11399;
wire     [31:0] n11400;
wire     [31:0] n11401;
wire     [31:0] n11402;
wire     [31:0] n11403;
wire     [31:0] n11404;
wire     [31:0] n11405;
wire     [31:0] n11406;
wire     [31:0] n11407;
wire     [31:0] n11408;
wire     [31:0] n11409;
wire     [31:0] n11410;
wire     [31:0] n11411;
wire     [31:0] n11412;
wire     [31:0] n11413;
wire     [31:0] n11414;
wire     [31:0] n11415;
wire     [31:0] n11416;
wire     [31:0] n11417;
wire     [31:0] n11418;
wire     [31:0] n11419;
wire     [31:0] n11420;
wire     [31:0] n11421;
wire     [31:0] n11422;
wire     [31:0] n11423;
wire     [31:0] n11424;
wire     [31:0] n11425;
wire     [31:0] n11426;
wire     [31:0] n11427;
wire     [31:0] n11428;
wire     [31:0] n11429;
wire     [31:0] n11430;
wire     [31:0] n11431;
wire     [31:0] n11432;
wire     [31:0] n11433;
wire     [31:0] n11434;
wire     [31:0] n11435;
wire     [31:0] n11436;
wire     [31:0] n11437;
wire     [31:0] n11438;
wire     [31:0] n11439;
wire     [31:0] n11440;
wire     [31:0] n11441;
wire     [31:0] n11442;
wire     [31:0] n11443;
wire     [31:0] n11444;
wire     [31:0] n11445;
wire     [31:0] n11446;
wire     [31:0] n11447;
wire     [31:0] n11448;
wire     [31:0] n11449;
wire     [31:0] n11450;
wire     [31:0] n11451;
wire     [31:0] n11452;
wire     [31:0] n11453;
wire     [31:0] n11454;
wire     [31:0] n11455;
wire     [31:0] n11456;
wire     [31:0] n11457;
wire     [31:0] n11458;
wire     [31:0] n11459;
wire     [31:0] n11460;
wire     [31:0] n11461;
wire     [31:0] n11462;
wire     [31:0] n11463;
wire     [31:0] n11464;
wire     [31:0] n11465;
wire     [31:0] n11466;
wire     [31:0] n11467;
wire     [31:0] n11468;
wire     [31:0] n11469;
wire     [31:0] n11470;
wire     [31:0] n11471;
wire     [31:0] n11472;
wire     [31:0] n11473;
wire     [31:0] n11474;
wire     [31:0] n11475;
wire     [31:0] n11476;
wire     [31:0] n11477;
wire     [31:0] n11478;
wire     [31:0] n11479;
wire     [31:0] n11480;
wire     [31:0] n11481;
wire     [31:0] n11482;
wire     [31:0] n11483;
wire     [31:0] n11484;
wire     [31:0] n11485;
wire     [31:0] n11486;
wire     [31:0] n11487;
wire     [31:0] n11488;
wire     [31:0] n11489;
wire     [31:0] n11490;
wire     [31:0] n11491;
wire     [31:0] n11492;
wire     [31:0] n11493;
wire     [31:0] n11494;
wire     [31:0] n11495;
wire     [31:0] n11496;
wire     [31:0] n11497;
wire     [31:0] n11498;
wire     [31:0] n11499;
wire     [31:0] n11500;
wire     [31:0] n11501;
wire     [31:0] n11502;
wire     [31:0] n11503;
wire     [31:0] n11504;
wire     [31:0] n11505;
wire     [31:0] n11506;
wire     [31:0] n11507;
wire     [31:0] n11508;
wire     [31:0] n11509;
wire            n11510;
wire            n11511;
wire     [31:0] n11512;
wire     [31:0] n11513;
wire     [31:0] n11514;
wire     [31:0] n11515;
wire     [31:0] n11516;
wire     [31:0] n11517;
wire     [31:0] n11518;
wire     [31:0] n11519;
wire     [31:0] n11520;
wire     [31:0] n11521;
wire     [31:0] n11522;
wire     [31:0] n11523;
wire     [31:0] n11524;
wire     [31:0] n11525;
wire     [31:0] n11526;
wire     [31:0] n11527;
wire     [31:0] n11528;
wire     [31:0] n11529;
wire     [31:0] n11530;
wire     [31:0] n11531;
wire     [31:0] n11532;
wire     [31:0] n11533;
wire     [31:0] n11534;
wire     [31:0] n11535;
wire     [31:0] n11536;
wire     [31:0] n11537;
wire     [31:0] n11538;
wire     [31:0] n11539;
wire     [31:0] n11540;
wire     [31:0] n11541;
wire     [31:0] n11542;
wire     [31:0] n11543;
wire     [31:0] n11544;
wire            n11545;
wire            n11546;
wire            n11547;
wire            n11548;
wire            n11549;
wire            n11550;
wire            n11551;
wire            n11552;
wire            n11553;
wire            n11554;
wire            n11555;
wire            n11556;
wire            n11557;
wire            n11558;
wire            n11559;
wire            n11560;
wire            n11561;
wire            n11562;
wire            n11563;
wire            n11564;
wire            n11565;
wire            n11566;
wire            n11567;
wire            n11568;
wire            n11569;
wire            n11570;
wire            n11571;
wire            n11572;
wire            n11573;
wire            n11574;
wire            n11575;
wire            n11576;
wire            n11577;
wire            n11578;
wire            n11579;
wire            n11580;
wire            n11581;
wire            n11582;
wire            n11583;
wire            n11584;
wire            n11585;
wire            n11586;
wire            n11587;
wire            n11588;
wire            n11589;
wire            n11590;
wire            n11591;
wire            n11592;
wire            n11593;
wire            n11594;
wire            n11595;
wire            n11596;
wire            n11597;
wire            n11598;
wire            n11599;
wire            n11600;
wire            n11601;
wire            n11602;
wire            n11603;
wire            n11604;
wire            n11605;
wire            n11606;
wire            n11607;
wire            n11608;
wire            n11609;
wire            n11610;
wire            n11611;
wire            n11612;
wire            n11613;
wire            n11614;
wire            n11615;
wire            n11616;
wire            n11617;
wire            n11618;
wire            n11619;
wire            n11620;
wire            n11621;
wire            n11622;
wire            n11623;
wire            n11624;
wire            n11625;
wire            n11626;
wire            n11627;
wire            n11628;
wire            n11629;
wire            n11630;
wire            n11631;
wire            n11632;
wire            n11633;
wire            n11634;
wire            n11635;
wire            n11636;
wire            n11637;
wire            n11638;
wire            n11639;
wire            n11640;
wire            n11641;
wire            n11642;
wire            n11643;
wire            n11644;
wire            n11645;
wire            n11646;
wire            n11647;
wire            n11648;
wire            n11649;
wire            n11650;
wire            n11651;
wire            n11652;
wire            n11653;
wire            n11654;
wire            n11655;
wire            n11656;
wire            n11657;
wire            n11658;
wire            n11659;
wire            n11660;
wire            n11661;
wire            n11662;
wire            n11663;
wire            n11664;
wire            n11665;
wire            n11666;
wire            n11667;
wire            n11668;
wire            n11669;
wire            n11670;
wire            n11671;
wire            n11672;
wire            n11673;
wire            n11674;
wire            n11675;
wire            n11676;
wire            n11677;
wire            n11678;
wire            n11679;
wire            n11680;
wire            n11681;
wire            n11682;
wire            n11683;
wire            n11684;
wire            n11685;
wire            n11686;
wire            n11687;
wire            n11688;
wire            n11689;
wire            n11690;
wire            n11691;
wire            n11692;
wire            n11693;
wire            n11694;
wire            n11695;
wire            n11696;
wire            n11697;
wire            n11698;
wire            n11699;
wire            n11700;
wire            n11701;
wire            n11702;
wire            n11703;
wire            n11704;
wire            n11705;
wire            n11706;
wire            n11707;
wire            n11708;
wire            n11709;
wire            n11710;
wire            n11711;
wire            n11712;
wire            n11713;
wire            n11714;
wire            n11715;
wire            n11716;
wire            n11717;
wire            n11718;
wire            n11719;
wire            n11720;
wire            n11721;
wire            n11722;
wire            n11723;
wire            n11724;
wire            n11725;
wire            n11726;
wire            n11727;
wire            n11728;
wire            n11729;
wire            n11730;
wire            n11731;
wire            n11732;
wire            n11733;
wire            n11734;
wire            n11735;
wire            n11736;
wire            n11737;
wire            n11738;
wire            n11739;
wire            n11740;
wire            n11741;
wire            n11742;
wire            n11743;
wire            n11744;
wire            n11745;
wire            n11746;
wire            n11747;
wire            n11748;
wire            n11749;
wire            n11750;
wire            n11751;
wire            n11752;
wire            n11753;
wire            n11754;
wire            n11755;
wire            n11756;
wire            n11757;
wire            n11758;
wire            n11759;
wire            n11760;
wire            n11761;
wire            n11762;
wire            n11763;
wire            n11764;
wire            n11765;
wire            n11766;
wire            n11767;
wire            n11768;
wire            n11769;
wire            n11770;
wire            n11771;
wire            n11772;
wire            n11773;
wire            n11774;
wire            n11775;
wire            n11776;
wire            n11777;
wire            n11778;
wire            n11779;
wire            n11780;
wire            n11781;
wire            n11782;
wire            n11783;
wire            n11784;
wire            n11785;
wire            n11786;
wire            n11787;
wire            n11788;
wire            n11789;
wire            n11790;
wire            n11791;
wire            n11792;
wire            n11793;
wire            n11794;
wire            n11795;
wire            n11796;
wire            n11797;
wire            n11798;
wire            n11799;
wire            n11800;
wire            n11801;
wire            n11802;
wire            n11803;
wire            n11804;
wire            n11805;
wire            n11806;
wire            n11807;
wire            n11808;
wire            n11809;
wire            n11810;
wire            n11811;
wire            n11812;
wire            n11813;
wire            n11814;
wire            n11815;
wire            n11816;
wire            n11817;
wire            n11818;
wire            n11819;
wire            n11820;
wire            n11821;
wire            n11822;
wire            n11823;
wire            n11824;
wire            n11825;
wire            n11826;
wire            n11827;
wire            n11828;
wire            n11829;
wire            n11830;
wire            n11831;
wire            n11832;
wire            n11833;
wire            n11834;
wire            n11835;
wire            n11836;
wire            n11837;
wire            n11838;
wire            n11839;
wire            n11840;
wire            n11841;
wire            n11842;
wire            n11843;
wire            n11844;
wire            n11845;
wire            n11846;
wire            n11847;
wire            n11848;
wire            n11849;
wire            n11850;
wire            n11851;
wire            n11852;
wire            n11853;
wire            n11854;
wire            n11855;
wire            n11856;
wire            n11857;
wire            n11858;
wire            n11859;
wire            n11860;
wire            n11861;
wire            n11862;
wire            n11863;
wire            n11864;
wire            n11865;
wire            n11866;
wire            n11867;
wire            n11868;
wire            n11869;
wire            n11870;
wire            n11871;
wire            n11872;
wire            n11873;
wire            n11874;
wire            n11875;
wire            n11876;
wire            n11877;
wire            n11878;
wire            n11879;
wire            n11880;
wire            n11881;
wire            n11882;
wire            n11883;
wire            n11884;
wire            n11885;
wire            n11886;
wire            n11887;
wire            n11888;
wire            n11889;
wire            n11890;
wire            n11891;
wire            n11892;
wire            n11893;
wire            n11894;
wire            n11895;
wire            n11896;
wire            n11897;
wire            n11898;
wire            n11899;
wire            n11900;
wire            n11901;
wire            n11902;
wire            n11903;
wire            n11904;
wire            n11905;
wire            n11906;
wire            n11907;
wire            n11908;
wire            n11909;
wire            n11910;
wire            n11911;
wire            n11912;
wire            n11913;
wire            n11914;
wire            n11915;
wire            n11916;
wire            n11917;
wire            n11918;
wire            n11919;
wire            n11920;
wire            n11921;
wire            n11922;
wire            n11923;
wire            n11924;
wire            n11925;
wire            n11926;
wire            n11927;
wire            n11928;
wire            n11929;
wire            n11930;
wire            n11931;
wire            n11932;
wire            n11933;
wire            n11934;
wire            n11935;
wire            n11936;
wire            n11937;
wire            n11938;
wire            n11939;
wire            n11940;
wire            n11941;
wire            n11942;
wire            n11943;
wire            n11944;
wire            n11945;
wire            n11946;
wire            n11947;
wire            n11948;
wire            n11949;
wire            n11950;
wire            n11951;
wire            n11952;
wire            n11953;
wire            n11954;
wire            n11955;
wire            n11956;
wire            n11957;
wire            n11958;
wire            n11959;
wire            n11960;
wire            n11961;
wire            n11962;
wire            n11963;
wire            n11964;
wire            n11965;
wire            n11966;
wire            n11967;
wire            n11968;
wire            n11969;
wire            n11970;
wire            n11971;
wire            n11972;
wire            n11973;
wire            n11974;
wire            n11975;
wire            n11976;
wire            n11977;
wire            n11978;
wire            n11979;
wire            n11980;
wire            n11981;
wire            n11982;
wire            n11983;
wire            n11984;
wire            n11985;
wire            n11986;
wire            n11987;
wire            n11988;
wire            n11989;
wire            n11990;
wire            n11991;
wire            n11992;
wire            n11993;
wire            n11994;
wire            n11995;
wire            n11996;
wire            n11997;
wire            n11998;
wire            n11999;
wire            n12000;
wire            n12001;
wire            n12002;
wire            n12003;
wire            n12004;
wire            n12005;
wire            n12006;
wire            n12007;
wire            n12008;
wire            n12009;
wire            n12010;
wire            n12011;
wire            n12012;
wire            n12013;
wire            n12014;
wire            n12015;
wire            n12016;
wire            n12017;
wire            n12018;
wire            n12019;
wire            n12020;
wire            n12021;
wire            n12022;
wire            n12023;
wire            n12024;
wire            n12025;
wire            n12026;
wire            n12027;
wire            n12028;
wire            n12029;
wire            n12030;
wire            n12031;
wire            n12032;
wire            n12033;
wire            n12034;
wire            n12035;
wire            n12036;
wire            n12037;
wire            n12038;
wire            n12039;
wire            n12040;
wire            n12041;
wire            n12042;
wire            n12043;
wire            n12044;
wire            n12045;
wire            n12046;
wire            n12047;
wire            n12048;
wire            n12049;
wire            n12050;
wire            n12051;
wire            n12052;
wire            n12053;
wire            n12054;
wire            n12055;
wire            n12056;
wire            n12057;
wire            n12058;
wire            n12059;
wire            n12060;
wire            n12061;
wire            n12062;
wire            n12063;
wire            n12064;
wire            n12065;
wire            n12066;
wire            n12067;
wire            n12068;
wire            n12069;
wire            n12070;
wire            n12071;
wire            n12072;
wire     [31:0] n12073;
wire     [31:0] n12074;
wire     [31:0] n12075;
wire     [31:0] n12076;
wire     [31:0] n12077;
wire     [31:0] n12078;
wire     [31:0] n12079;
wire     [31:0] n12080;
wire     [31:0] n12081;
wire     [31:0] n12082;
wire     [31:0] n12083;
wire     [31:0] n12084;
wire     [31:0] n12085;
wire     [31:0] n12086;
wire     [31:0] n12087;
wire     [31:0] n12088;
wire     [31:0] n12089;
wire     [31:0] n12090;
wire     [31:0] n12091;
wire     [31:0] n12092;
wire     [31:0] n12093;
wire     [31:0] n12094;
wire     [31:0] n12095;
wire     [31:0] n12096;
wire     [31:0] n12097;
wire     [31:0] n12098;
wire     [31:0] n12099;
wire     [31:0] n12100;
wire     [31:0] n12101;
wire     [31:0] n12102;
wire     [31:0] n12103;
wire     [31:0] n12104;
wire     [31:0] n12105;
wire     [31:0] n12106;
wire     [31:0] n12107;
wire     [31:0] n12108;
wire     [31:0] n12109;
wire     [31:0] n12110;
wire     [31:0] n12111;
wire     [31:0] n12112;
wire     [31:0] n12113;
wire     [31:0] n12114;
wire     [31:0] n12115;
wire     [31:0] n12116;
wire     [31:0] n12117;
wire     [31:0] n12118;
wire     [31:0] n12119;
wire     [31:0] n12120;
wire     [31:0] n12121;
wire     [31:0] n12122;
wire     [31:0] n12123;
wire     [31:0] n12124;
wire     [31:0] n12125;
wire     [31:0] n12126;
wire     [31:0] n12127;
wire     [31:0] n12128;
wire     [31:0] n12129;
wire     [31:0] n12130;
wire     [31:0] n12131;
wire     [31:0] n12132;
wire     [31:0] n12133;
wire     [31:0] n12134;
wire     [31:0] n12135;
wire     [31:0] n12136;
wire     [31:0] n12137;
wire     [31:0] n12138;
wire     [31:0] n12139;
wire     [31:0] n12140;
wire     [31:0] n12141;
wire     [31:0] n12142;
wire     [31:0] n12143;
wire     [31:0] n12144;
wire     [31:0] n12145;
wire     [31:0] n12146;
wire     [31:0] n12147;
wire     [31:0] n12148;
wire     [31:0] n12149;
wire     [31:0] n12150;
wire     [31:0] n12151;
wire     [31:0] n12152;
wire     [31:0] n12153;
wire     [31:0] n12154;
wire     [31:0] n12155;
wire     [31:0] n12156;
wire     [31:0] n12157;
wire     [31:0] n12158;
wire     [31:0] n12159;
wire     [31:0] n12160;
wire     [31:0] n12161;
wire     [31:0] n12162;
wire     [31:0] n12163;
wire     [31:0] n12164;
wire     [31:0] n12165;
wire     [31:0] n12166;
wire     [31:0] n12167;
wire     [31:0] n12168;
wire     [31:0] n12169;
wire     [31:0] n12170;
wire     [31:0] n12171;
wire     [31:0] n12172;
wire     [31:0] n12173;
wire     [31:0] n12174;
wire     [31:0] n12175;
wire     [31:0] n12176;
wire     [31:0] n12177;
wire     [31:0] n12178;
wire     [31:0] n12179;
wire     [31:0] n12180;
wire     [31:0] n12181;
wire     [31:0] n12182;
wire     [31:0] n12183;
wire     [31:0] n12184;
wire     [31:0] n12185;
wire     [31:0] n12186;
wire     [31:0] n12187;
wire     [31:0] n12188;
wire     [31:0] n12189;
wire     [31:0] n12190;
wire     [31:0] n12191;
wire     [31:0] n12192;
wire     [31:0] n12193;
wire     [31:0] n12194;
wire     [31:0] n12195;
wire     [31:0] n12196;
wire     [31:0] n12197;
wire     [31:0] n12198;
wire     [31:0] n12199;
wire     [31:0] n12200;
wire     [31:0] n12201;
wire     [31:0] n12202;
wire     [31:0] n12203;
wire     [31:0] n12204;
wire     [31:0] n12205;
wire     [31:0] n12206;
wire     [31:0] n12207;
wire     [31:0] n12208;
wire     [31:0] n12209;
wire     [31:0] n12210;
wire     [31:0] n12211;
wire     [31:0] n12212;
wire     [31:0] n12213;
wire     [31:0] n12214;
wire     [31:0] n12215;
wire     [31:0] n12216;
wire     [31:0] n12217;
wire     [31:0] n12218;
wire     [31:0] n12219;
wire     [31:0] n12220;
wire     [31:0] n12221;
wire     [31:0] n12222;
wire     [31:0] n12223;
wire     [31:0] n12224;
wire     [31:0] n12225;
wire     [31:0] n12226;
wire     [31:0] n12227;
wire     [31:0] n12228;
wire     [31:0] n12229;
wire     [31:0] n12230;
wire     [31:0] n12231;
wire     [31:0] n12232;
wire     [31:0] n12233;
wire     [31:0] n12234;
wire     [31:0] n12235;
wire     [31:0] n12236;
wire     [31:0] n12237;
wire     [31:0] n12238;
wire     [31:0] n12239;
wire     [31:0] n12240;
wire     [31:0] n12241;
wire     [31:0] n12242;
wire     [31:0] n12243;
wire     [31:0] n12244;
wire     [31:0] n12245;
wire     [31:0] n12246;
wire     [31:0] n12247;
wire     [31:0] n12248;
wire     [31:0] n12249;
wire     [31:0] n12250;
wire     [31:0] n12251;
wire     [31:0] n12252;
wire     [31:0] n12253;
wire     [31:0] n12254;
wire     [31:0] n12255;
wire     [31:0] n12256;
wire     [31:0] n12257;
wire     [31:0] n12258;
wire     [31:0] n12259;
wire     [31:0] n12260;
wire     [31:0] n12261;
wire     [31:0] n12262;
wire     [31:0] n12263;
wire     [31:0] n12264;
wire     [31:0] n12265;
wire     [31:0] n12266;
wire     [31:0] n12267;
wire     [31:0] n12268;
wire     [31:0] n12269;
wire     [31:0] n12270;
wire     [31:0] n12271;
wire     [31:0] n12272;
wire     [31:0] n12273;
wire     [31:0] n12274;
wire     [31:0] n12275;
wire     [31:0] n12276;
wire     [31:0] n12277;
wire     [31:0] n12278;
wire     [31:0] n12279;
wire     [31:0] n12280;
wire     [31:0] n12281;
wire     [31:0] n12282;
wire     [31:0] n12283;
wire     [31:0] n12284;
wire     [31:0] n12285;
wire     [31:0] n12286;
wire     [31:0] n12287;
wire     [31:0] n12288;
wire     [31:0] n12289;
wire     [31:0] n12290;
wire     [31:0] n12291;
wire     [31:0] n12292;
wire     [31:0] n12293;
wire     [31:0] n12294;
wire     [31:0] n12295;
wire     [31:0] n12296;
wire     [31:0] n12297;
wire     [31:0] n12298;
wire     [31:0] n12299;
wire     [31:0] n12300;
wire     [31:0] n12301;
wire     [31:0] n12302;
wire     [31:0] n12303;
wire     [31:0] n12304;
wire     [31:0] n12305;
wire     [31:0] n12306;
wire     [31:0] n12307;
wire     [31:0] n12308;
wire     [31:0] n12309;
wire     [31:0] n12310;
wire     [31:0] n12311;
wire     [31:0] n12312;
wire     [31:0] n12313;
wire     [31:0] n12314;
wire     [31:0] n12315;
wire     [31:0] n12316;
wire     [31:0] n12317;
wire     [31:0] n12318;
wire     [31:0] n12319;
wire     [31:0] n12320;
wire     [31:0] n12321;
wire     [31:0] n12322;
wire     [31:0] n12323;
wire     [31:0] n12324;
wire     [31:0] n12325;
wire     [31:0] n12326;
wire     [31:0] n12327;
wire     [31:0] n12328;
wire     [31:0] n12329;
wire     [31:0] n12330;
wire     [31:0] n12331;
wire     [31:0] n12332;
wire     [31:0] n12333;
wire     [31:0] n12334;
wire     [31:0] n12335;
wire     [31:0] n12336;
wire     [31:0] n12337;
wire     [31:0] n12338;
wire     [31:0] n12339;
wire     [31:0] n12340;
wire     [31:0] n12341;
wire     [31:0] n12342;
wire     [31:0] n12343;
wire     [31:0] n12344;
wire     [31:0] n12345;
wire     [31:0] n12346;
wire     [31:0] n12347;
wire     [31:0] n12348;
wire     [31:0] n12349;
wire     [31:0] n12350;
wire     [31:0] n12351;
wire     [31:0] n12352;
wire     [31:0] n12353;
wire     [31:0] n12354;
wire     [31:0] n12355;
wire     [31:0] n12356;
wire     [31:0] n12357;
wire     [31:0] n12358;
wire     [31:0] n12359;
wire     [31:0] n12360;
wire     [31:0] n12361;
wire     [31:0] n12362;
wire     [31:0] n12363;
wire     [31:0] n12364;
wire     [31:0] n12365;
wire     [31:0] n12366;
wire     [31:0] n12367;
wire     [31:0] n12368;
wire     [31:0] n12369;
wire     [31:0] n12370;
wire     [31:0] n12371;
wire     [31:0] n12372;
wire     [31:0] n12373;
wire     [31:0] n12374;
wire     [31:0] n12375;
wire     [31:0] n12376;
wire     [31:0] n12377;
wire     [31:0] n12378;
wire     [31:0] n12379;
wire     [31:0] n12380;
wire     [31:0] n12381;
wire     [31:0] n12382;
wire     [31:0] n12383;
wire     [31:0] n12384;
wire     [31:0] n12385;
wire     [31:0] n12386;
wire     [31:0] n12387;
wire     [31:0] n12388;
wire     [31:0] n12389;
wire     [31:0] n12390;
wire     [31:0] n12391;
wire     [31:0] n12392;
wire     [31:0] n12393;
wire     [31:0] n12394;
wire     [31:0] n12395;
wire     [31:0] n12396;
wire     [31:0] n12397;
wire     [31:0] n12398;
wire     [31:0] n12399;
wire     [31:0] n12400;
wire     [31:0] n12401;
wire     [31:0] n12402;
wire     [31:0] n12403;
wire     [31:0] n12404;
wire     [31:0] n12405;
wire     [31:0] n12406;
wire     [31:0] n12407;
wire     [31:0] n12408;
wire     [31:0] n12409;
wire     [31:0] n12410;
wire     [31:0] n12411;
wire     [31:0] n12412;
wire     [31:0] n12413;
wire     [31:0] n12414;
wire     [31:0] n12415;
wire     [31:0] n12416;
wire     [31:0] n12417;
wire     [31:0] n12418;
wire     [31:0] n12419;
wire     [31:0] n12420;
wire     [31:0] n12421;
wire     [31:0] n12422;
wire     [31:0] n12423;
wire     [31:0] n12424;
wire     [31:0] n12425;
wire     [31:0] n12426;
wire     [31:0] n12427;
wire     [31:0] n12428;
wire     [31:0] n12429;
wire     [31:0] n12430;
wire     [31:0] n12431;
wire     [31:0] n12432;
wire     [31:0] n12433;
wire     [31:0] n12434;
wire     [31:0] n12435;
wire     [31:0] n12436;
wire     [31:0] n12437;
wire     [31:0] n12438;
wire     [31:0] n12439;
wire     [31:0] n12440;
wire     [31:0] n12441;
wire     [31:0] n12442;
wire     [31:0] n12443;
wire     [31:0] n12444;
wire     [31:0] n12445;
wire     [31:0] n12446;
wire     [31:0] n12447;
wire     [31:0] n12448;
wire     [31:0] n12449;
wire     [31:0] n12450;
wire     [31:0] n12451;
wire     [31:0] n12452;
wire     [31:0] n12453;
wire     [31:0] n12454;
wire     [31:0] n12455;
wire     [31:0] n12456;
wire     [31:0] n12457;
wire     [31:0] n12458;
wire     [31:0] n12459;
wire     [31:0] n12460;
wire     [31:0] n12461;
wire     [31:0] n12462;
wire     [31:0] n12463;
wire     [31:0] n12464;
wire     [31:0] n12465;
wire     [31:0] n12466;
wire     [31:0] n12467;
wire     [31:0] n12468;
wire     [31:0] n12469;
wire     [31:0] n12470;
wire     [31:0] n12471;
wire     [31:0] n12472;
wire     [31:0] n12473;
wire     [31:0] n12474;
wire     [31:0] n12475;
wire     [31:0] n12476;
wire     [31:0] n12477;
wire     [31:0] n12478;
wire     [31:0] n12479;
wire     [31:0] n12480;
wire     [31:0] n12481;
wire     [31:0] n12482;
wire     [31:0] n12483;
wire     [31:0] n12484;
wire     [31:0] n12485;
wire     [31:0] n12486;
wire     [31:0] n12487;
wire     [31:0] n12488;
wire     [31:0] n12489;
wire     [31:0] n12490;
wire     [31:0] n12491;
wire     [31:0] n12492;
wire     [31:0] n12493;
wire     [31:0] n12494;
wire     [31:0] n12495;
wire     [31:0] n12496;
wire     [31:0] n12497;
wire     [31:0] n12498;
wire     [31:0] n12499;
wire     [31:0] n12500;
wire     [31:0] n12501;
wire     [31:0] n12502;
wire     [31:0] n12503;
wire     [31:0] n12504;
wire     [31:0] n12505;
wire     [31:0] n12506;
wire     [31:0] n12507;
wire     [31:0] n12508;
wire     [31:0] n12509;
wire     [31:0] n12510;
wire     [31:0] n12511;
wire     [31:0] n12512;
wire     [31:0] n12513;
wire     [31:0] n12514;
wire     [31:0] n12515;
wire     [31:0] n12516;
wire     [31:0] n12517;
wire     [31:0] n12518;
wire     [31:0] n12519;
wire     [31:0] n12520;
wire     [31:0] n12521;
wire     [31:0] n12522;
wire     [31:0] n12523;
wire     [31:0] n12524;
wire     [31:0] n12525;
wire     [31:0] n12526;
wire     [31:0] n12527;
wire     [31:0] n12528;
wire     [31:0] n12529;
wire     [31:0] n12530;
wire     [31:0] n12531;
wire     [31:0] n12532;
wire     [31:0] n12533;
wire     [31:0] n12534;
wire     [31:0] n12535;
wire     [31:0] n12536;
wire     [31:0] n12537;
wire     [31:0] n12538;
wire     [31:0] n12539;
wire     [31:0] n12540;
wire     [31:0] n12541;
wire     [31:0] n12542;
wire     [31:0] n12543;
wire     [31:0] n12544;
wire     [31:0] n12545;
wire     [31:0] n12546;
wire     [31:0] n12547;
wire     [31:0] n12548;
wire     [31:0] n12549;
wire     [31:0] n12550;
wire     [31:0] n12551;
wire     [31:0] n12552;
wire     [31:0] n12553;
wire     [31:0] n12554;
wire     [31:0] n12555;
wire     [31:0] n12556;
wire     [31:0] n12557;
wire     [31:0] n12558;
wire     [31:0] n12559;
wire     [31:0] n12560;
wire     [31:0] n12561;
wire     [31:0] n12562;
wire     [31:0] n12563;
wire     [31:0] n12564;
wire     [31:0] n12565;
wire     [31:0] n12566;
wire     [31:0] n12567;
wire     [31:0] n12568;
wire     [31:0] n12569;
wire     [31:0] n12570;
wire     [31:0] n12571;
wire     [31:0] n12572;
wire     [31:0] n12573;
wire     [31:0] n12574;
wire     [31:0] n12575;
wire     [31:0] n12576;
wire     [31:0] n12577;
wire     [31:0] n12578;
wire     [31:0] n12579;
wire     [31:0] n12580;
wire     [31:0] n12581;
wire     [31:0] n12582;
wire     [31:0] n12583;
wire     [31:0] n12584;
wire     [31:0] n12585;
wire     [31:0] n12586;
wire     [31:0] n12587;
wire     [31:0] n12588;
wire     [31:0] n12589;
wire     [31:0] n12590;
wire     [31:0] n12591;
wire     [31:0] n12592;
wire     [31:0] n12593;
wire     [31:0] n12594;
wire            n12595;
wire            n12596;
wire            n12597;
wire            n12598;
wire            n12599;
wire            n12600;
wire            n12601;
wire            n12602;
wire            n12603;
wire            n12604;
wire            n12605;
wire            n12606;
wire            n12607;
wire            n12608;
wire            n12609;
wire            n12610;
wire            n12611;
wire            n12612;
wire            n12613;
wire            n12614;
wire            n12615;
wire            n12616;
wire            n12617;
wire            n12618;
wire            n12619;
wire            n12620;
wire            n12621;
wire            n12622;
wire            n12623;
wire            n12624;
wire            n12625;
wire            n12626;
wire            n12627;
wire            n12628;
wire            n12629;
wire            n12630;
wire            n12631;
wire            n12632;
wire            n12633;
wire            n12634;
wire            n12635;
wire            n12636;
wire            n12637;
wire            n12638;
wire            n12639;
wire            n12640;
wire            n12641;
wire            n12642;
wire            n12643;
wire            n12644;
wire            n12645;
wire            n12646;
wire            n12647;
wire            n12648;
wire            n12649;
wire            n12650;
wire            n12651;
wire            n12652;
wire            n12653;
wire            n12654;
wire            n12655;
wire            n12656;
wire            n12657;
wire            n12658;
wire            n12659;
wire            n12660;
wire            n12661;
wire            n12662;
wire            n12663;
wire            n12664;
wire            n12665;
wire            n12666;
wire            n12667;
wire            n12668;
wire            n12669;
wire            n12670;
wire            n12671;
wire            n12672;
wire            n12673;
wire            n12674;
wire            n12675;
wire            n12676;
wire            n12677;
wire            n12678;
wire            n12679;
wire            n12680;
wire            n12681;
wire            n12682;
wire            n12683;
wire            n12684;
wire            n12685;
wire            n12686;
wire            n12687;
wire            n12688;
wire            n12689;
wire            n12690;
wire            n12691;
wire            n12692;
wire            n12693;
wire            n12694;
wire            n12695;
wire            n12696;
wire            n12697;
wire            n12698;
wire            n12699;
wire            n12700;
wire            n12701;
wire            n12702;
wire            n12703;
wire            n12704;
wire            n12705;
wire            n12706;
wire            n12707;
wire            n12708;
wire            n12709;
wire            n12710;
wire            n12711;
wire            n12712;
wire            n12713;
wire            n12714;
wire            n12715;
wire            n12716;
wire            n12717;
wire            n12718;
wire            n12719;
wire            n12720;
wire            n12721;
wire            n12722;
wire            n12723;
wire            n12724;
wire            n12725;
wire            n12726;
wire            n12727;
wire            n12728;
wire            n12729;
wire            n12730;
wire            n12731;
wire            n12732;
wire            n12733;
wire            n12734;
wire            n12735;
wire            n12736;
wire            n12737;
wire            n12738;
wire            n12739;
wire            n12740;
wire            n12741;
wire            n12742;
wire            n12743;
wire            n12744;
wire            n12745;
wire            n12746;
wire            n12747;
wire            n12748;
wire            n12749;
wire            n12750;
wire            n12751;
wire            n12752;
wire            n12753;
wire            n12754;
wire            n12755;
wire            n12756;
wire            n12757;
wire            n12758;
wire            n12759;
wire            n12760;
wire            n12761;
wire            n12762;
wire            n12763;
wire            n12764;
wire            n12765;
wire            n12766;
wire            n12767;
wire            n12768;
wire            n12769;
wire            n12770;
wire            n12771;
wire            n12772;
wire            n12773;
wire            n12774;
wire            n12775;
wire            n12776;
wire            n12777;
wire            n12778;
wire            n12779;
wire            n12780;
wire            n12781;
wire            n12782;
wire            n12783;
wire            n12784;
wire            n12785;
wire            n12786;
wire            n12787;
wire            n12788;
wire            n12789;
wire            n12790;
wire            n12791;
wire            n12792;
wire            n12793;
wire            n12794;
wire            n12795;
wire            n12796;
wire            n12797;
wire            n12798;
wire            n12799;
wire            n12800;
wire            n12801;
wire            n12802;
wire            n12803;
wire            n12804;
wire            n12805;
wire            n12806;
wire            n12807;
wire            n12808;
wire            n12809;
wire            n12810;
wire            n12811;
wire            n12812;
wire            n12813;
wire            n12814;
wire            n12815;
wire            n12816;
wire            n12817;
wire            n12818;
wire            n12819;
wire            n12820;
wire            n12821;
wire            n12822;
wire            n12823;
wire            n12824;
wire            n12825;
wire            n12826;
wire            n12827;
wire            n12828;
wire            n12829;
wire            n12830;
wire            n12831;
wire            n12832;
wire            n12833;
wire            n12834;
wire            n12835;
wire            n12836;
wire            n12837;
wire            n12838;
wire            n12839;
wire            n12840;
wire            n12841;
wire            n12842;
wire            n12843;
wire            n12844;
wire            n12845;
wire            n12846;
wire            n12847;
wire            n12848;
wire            n12849;
wire            n12850;
wire            n12851;
wire            n12852;
wire            n12853;
wire            n12854;
wire            n12855;
wire            n12856;
wire            n12857;
wire            n12858;
wire            n12859;
wire            n12860;
wire            n12861;
wire            n12862;
wire            n12863;
wire            n12864;
wire            n12865;
wire            n12866;
wire            n12867;
wire            n12868;
wire            n12869;
wire            n12870;
wire            n12871;
wire            n12872;
wire            n12873;
wire            n12874;
wire            n12875;
wire            n12876;
wire            n12877;
wire            n12878;
wire            n12879;
wire            n12880;
wire            n12881;
wire            n12882;
wire            n12883;
wire            n12884;
wire            n12885;
wire            n12886;
wire            n12887;
wire            n12888;
wire            n12889;
wire            n12890;
wire            n12891;
wire            n12892;
wire            n12893;
wire            n12894;
wire            n12895;
wire            n12896;
wire            n12897;
wire            n12898;
wire            n12899;
wire            n12900;
wire            n12901;
wire            n12902;
wire            n12903;
wire            n12904;
wire            n12905;
wire            n12906;
wire            n12907;
wire            n12908;
wire            n12909;
wire            n12910;
wire            n12911;
wire            n12912;
wire            n12913;
wire            n12914;
wire            n12915;
wire            n12916;
wire            n12917;
wire            n12918;
wire            n12919;
wire            n12920;
wire            n12921;
wire            n12922;
wire            n12923;
wire            n12924;
wire            n12925;
wire            n12926;
wire            n12927;
wire            n12928;
wire            n12929;
wire            n12930;
wire            n12931;
wire            n12932;
wire            n12933;
wire            n12934;
wire            n12935;
wire            n12936;
wire            n12937;
wire            n12938;
wire            n12939;
wire            n12940;
wire            n12941;
wire            n12942;
wire            n12943;
wire            n12944;
wire            n12945;
wire            n12946;
wire            n12947;
wire            n12948;
wire            n12949;
wire            n12950;
wire            n12951;
wire            n12952;
wire            n12953;
wire            n12954;
wire            n12955;
wire            n12956;
wire            n12957;
wire            n12958;
wire            n12959;
wire            n12960;
wire            n12961;
wire            n12962;
wire            n12963;
wire            n12964;
wire            n12965;
wire            n12966;
wire            n12967;
wire            n12968;
wire            n12969;
wire            n12970;
wire            n12971;
wire            n12972;
wire            n12973;
wire            n12974;
wire            n12975;
wire            n12976;
wire            n12977;
wire            n12978;
wire            n12979;
wire            n12980;
wire            n12981;
wire            n12982;
wire            n12983;
wire            n12984;
wire            n12985;
wire            n12986;
wire            n12987;
wire            n12988;
wire            n12989;
wire            n12990;
wire            n12991;
wire            n12992;
wire            n12993;
wire            n12994;
wire            n12995;
wire            n12996;
wire            n12997;
wire            n12998;
wire            n12999;
wire            n13000;
wire            n13001;
wire            n13002;
wire            n13003;
wire            n13004;
wire            n13005;
wire            n13006;
wire            n13007;
wire            n13008;
wire            n13009;
wire            n13010;
wire            n13011;
wire            n13012;
wire            n13013;
wire            n13014;
wire            n13015;
wire            n13016;
wire            n13017;
wire            n13018;
wire            n13019;
wire            n13020;
wire            n13021;
wire            n13022;
wire            n13023;
wire            n13024;
wire            n13025;
wire            n13026;
wire            n13027;
wire            n13028;
wire            n13029;
wire            n13030;
wire            n13031;
wire            n13032;
wire            n13033;
wire            n13034;
wire            n13035;
wire            n13036;
wire            n13037;
wire            n13038;
wire            n13039;
wire            n13040;
wire            n13041;
wire            n13042;
wire            n13043;
wire            n13044;
wire            n13045;
wire            n13046;
wire            n13047;
wire            n13048;
wire            n13049;
wire            n13050;
wire            n13051;
wire            n13052;
wire            n13053;
wire            n13054;
wire            n13055;
wire            n13056;
wire            n13057;
wire            n13058;
wire            n13059;
wire            n13060;
wire            n13061;
wire            n13062;
wire            n13063;
wire            n13064;
wire            n13065;
wire            n13066;
wire            n13067;
wire            n13068;
wire            n13069;
wire            n13070;
wire            n13071;
wire            n13072;
wire            n13073;
wire            n13074;
wire            n13075;
wire            n13076;
wire            n13077;
wire            n13078;
wire            n13079;
wire            n13080;
wire            n13081;
wire            n13082;
wire            n13083;
wire            n13084;
wire            n13085;
wire            n13086;
wire            n13087;
wire            n13088;
wire            n13089;
wire            n13090;
wire            n13091;
wire            n13092;
wire            n13093;
wire            n13094;
wire            n13095;
wire            n13096;
wire            n13097;
wire            n13098;
wire            n13099;
wire            n13100;
wire            n13101;
wire            n13102;
wire            n13103;
wire            n13104;
wire            n13105;
wire            n13106;
wire     [31:0] n13107;
wire     [31:0] n13108;
wire     [31:0] n13109;
wire     [31:0] n13110;
wire     [31:0] n13111;
wire     [31:0] n13112;
wire     [31:0] n13113;
wire     [31:0] n13114;
wire     [31:0] n13115;
wire     [31:0] n13116;
wire     [31:0] n13117;
wire     [31:0] n13118;
wire     [31:0] n13119;
wire     [31:0] n13120;
wire     [31:0] n13121;
wire     [31:0] n13122;
wire     [31:0] n13123;
wire     [31:0] n13124;
wire     [31:0] n13125;
wire     [31:0] n13126;
wire     [31:0] n13127;
wire     [31:0] n13128;
wire     [31:0] n13129;
wire     [31:0] n13130;
wire     [31:0] n13131;
wire     [31:0] n13132;
wire     [31:0] n13133;
wire     [31:0] n13134;
wire     [31:0] n13135;
wire     [31:0] n13136;
wire     [31:0] n13137;
wire     [31:0] n13138;
wire     [31:0] n13139;
wire     [31:0] n13140;
wire     [31:0] n13141;
wire     [31:0] n13142;
wire     [31:0] n13143;
wire     [31:0] n13144;
wire     [31:0] n13145;
wire     [31:0] n13146;
wire     [31:0] n13147;
wire     [31:0] n13148;
wire     [31:0] n13149;
wire     [31:0] n13150;
wire     [31:0] n13151;
wire     [31:0] n13152;
wire     [31:0] n13153;
wire     [31:0] n13154;
wire     [31:0] n13155;
wire     [31:0] n13156;
wire     [31:0] n13157;
wire     [31:0] n13158;
wire     [31:0] n13159;
wire     [31:0] n13160;
wire     [31:0] n13161;
wire     [31:0] n13162;
wire     [31:0] n13163;
wire     [31:0] n13164;
wire     [31:0] n13165;
wire     [31:0] n13166;
wire     [31:0] n13167;
wire     [31:0] n13168;
wire     [31:0] n13169;
wire     [31:0] n13170;
wire     [31:0] n13171;
wire     [31:0] n13172;
wire     [31:0] n13173;
wire     [31:0] n13174;
wire     [31:0] n13175;
wire     [31:0] n13176;
wire     [31:0] n13177;
wire     [31:0] n13178;
wire     [31:0] n13179;
wire     [31:0] n13180;
wire     [31:0] n13181;
wire     [31:0] n13182;
wire     [31:0] n13183;
wire     [31:0] n13184;
wire     [31:0] n13185;
wire     [31:0] n13186;
wire     [31:0] n13187;
wire     [31:0] n13188;
wire     [31:0] n13189;
wire     [31:0] n13190;
wire     [31:0] n13191;
wire     [31:0] n13192;
wire     [31:0] n13193;
wire     [31:0] n13194;
wire     [31:0] n13195;
wire     [31:0] n13196;
wire     [31:0] n13197;
wire     [31:0] n13198;
wire     [31:0] n13199;
wire     [31:0] n13200;
wire     [31:0] n13201;
wire     [31:0] n13202;
wire     [31:0] n13203;
wire     [31:0] n13204;
wire     [31:0] n13205;
wire     [31:0] n13206;
wire     [31:0] n13207;
wire     [31:0] n13208;
wire     [31:0] n13209;
wire     [31:0] n13210;
wire     [31:0] n13211;
wire     [31:0] n13212;
wire     [31:0] n13213;
wire     [31:0] n13214;
wire     [31:0] n13215;
wire     [31:0] n13216;
wire     [31:0] n13217;
wire     [31:0] n13218;
wire     [31:0] n13219;
wire     [31:0] n13220;
wire     [31:0] n13221;
wire     [31:0] n13222;
wire     [31:0] n13223;
wire     [31:0] n13224;
wire     [31:0] n13225;
wire     [31:0] n13226;
wire     [31:0] n13227;
wire     [31:0] n13228;
wire     [31:0] n13229;
wire     [31:0] n13230;
wire     [31:0] n13231;
wire     [31:0] n13232;
wire     [31:0] n13233;
wire     [31:0] n13234;
wire     [31:0] n13235;
wire     [31:0] n13236;
wire     [31:0] n13237;
wire     [31:0] n13238;
wire     [31:0] n13239;
wire     [31:0] n13240;
wire     [31:0] n13241;
wire     [31:0] n13242;
wire     [31:0] n13243;
wire     [31:0] n13244;
wire     [31:0] n13245;
wire     [31:0] n13246;
wire     [31:0] n13247;
wire     [31:0] n13248;
wire     [31:0] n13249;
wire     [31:0] n13250;
wire     [31:0] n13251;
wire     [31:0] n13252;
wire     [31:0] n13253;
wire     [31:0] n13254;
wire     [31:0] n13255;
wire     [31:0] n13256;
wire     [31:0] n13257;
wire     [31:0] n13258;
wire     [31:0] n13259;
wire     [31:0] n13260;
wire     [31:0] n13261;
wire     [31:0] n13262;
wire     [31:0] n13263;
wire     [31:0] n13264;
wire     [31:0] n13265;
wire     [31:0] n13266;
wire     [31:0] n13267;
wire     [31:0] n13268;
wire     [31:0] n13269;
wire     [31:0] n13270;
wire     [31:0] n13271;
wire     [31:0] n13272;
wire     [31:0] n13273;
wire     [31:0] n13274;
wire     [31:0] n13275;
wire     [31:0] n13276;
wire     [31:0] n13277;
wire     [31:0] n13278;
wire     [31:0] n13279;
wire     [31:0] n13280;
wire     [31:0] n13281;
wire     [31:0] n13282;
wire     [31:0] n13283;
wire     [31:0] n13284;
wire     [31:0] n13285;
wire     [31:0] n13286;
wire     [31:0] n13287;
wire     [31:0] n13288;
wire     [31:0] n13289;
wire     [31:0] n13290;
wire     [31:0] n13291;
wire     [31:0] n13292;
wire     [31:0] n13293;
wire     [31:0] n13294;
wire     [31:0] n13295;
wire     [31:0] n13296;
wire     [31:0] n13297;
wire     [31:0] n13298;
wire     [31:0] n13299;
wire     [31:0] n13300;
wire     [31:0] n13301;
wire     [31:0] n13302;
wire     [31:0] n13303;
wire     [31:0] n13304;
wire     [31:0] n13305;
wire     [31:0] n13306;
wire     [31:0] n13307;
wire     [31:0] n13308;
wire     [31:0] n13309;
wire     [31:0] n13310;
wire     [31:0] n13311;
wire     [31:0] n13312;
wire     [31:0] n13313;
wire     [31:0] n13314;
wire     [31:0] n13315;
wire     [31:0] n13316;
wire     [31:0] n13317;
wire     [31:0] n13318;
wire     [31:0] n13319;
wire     [31:0] n13320;
wire     [31:0] n13321;
wire     [31:0] n13322;
wire     [31:0] n13323;
wire     [31:0] n13324;
wire     [31:0] n13325;
wire     [31:0] n13326;
wire     [31:0] n13327;
wire     [31:0] n13328;
wire     [31:0] n13329;
wire     [31:0] n13330;
wire     [31:0] n13331;
wire     [31:0] n13332;
wire     [31:0] n13333;
wire     [31:0] n13334;
wire     [31:0] n13335;
wire     [31:0] n13336;
wire     [31:0] n13337;
wire     [31:0] n13338;
wire     [31:0] n13339;
wire     [31:0] n13340;
wire     [31:0] n13341;
wire     [31:0] n13342;
wire     [31:0] n13343;
wire     [31:0] n13344;
wire     [31:0] n13345;
wire     [31:0] n13346;
wire     [31:0] n13347;
wire     [31:0] n13348;
wire     [31:0] n13349;
wire     [31:0] n13350;
wire     [31:0] n13351;
wire     [31:0] n13352;
wire     [31:0] n13353;
wire     [31:0] n13354;
wire     [31:0] n13355;
wire     [31:0] n13356;
wire     [31:0] n13357;
wire     [31:0] n13358;
wire     [31:0] n13359;
wire     [31:0] n13360;
wire     [31:0] n13361;
wire     [31:0] n13362;
wire     [31:0] n13363;
wire     [31:0] n13364;
wire     [31:0] n13365;
wire     [31:0] n13366;
wire     [31:0] n13367;
wire     [31:0] n13368;
wire     [31:0] n13369;
wire     [31:0] n13370;
wire     [31:0] n13371;
wire     [31:0] n13372;
wire     [31:0] n13373;
wire     [31:0] n13374;
wire     [31:0] n13375;
wire     [31:0] n13376;
wire     [31:0] n13377;
wire     [31:0] n13378;
wire     [31:0] n13379;
wire     [31:0] n13380;
wire     [31:0] n13381;
wire     [31:0] n13382;
wire     [31:0] n13383;
wire     [31:0] n13384;
wire     [31:0] n13385;
wire     [31:0] n13386;
wire     [31:0] n13387;
wire     [31:0] n13388;
wire     [31:0] n13389;
wire     [31:0] n13390;
wire     [31:0] n13391;
wire     [31:0] n13392;
wire     [31:0] n13393;
wire     [31:0] n13394;
wire     [31:0] n13395;
wire     [31:0] n13396;
wire     [31:0] n13397;
wire     [31:0] n13398;
wire     [31:0] n13399;
wire     [31:0] n13400;
wire     [31:0] n13401;
wire     [31:0] n13402;
wire     [31:0] n13403;
wire     [31:0] n13404;
wire     [31:0] n13405;
wire     [31:0] n13406;
wire     [31:0] n13407;
wire     [31:0] n13408;
wire     [31:0] n13409;
wire     [31:0] n13410;
wire     [31:0] n13411;
wire     [31:0] n13412;
wire     [31:0] n13413;
wire     [31:0] n13414;
wire     [31:0] n13415;
wire     [31:0] n13416;
wire     [31:0] n13417;
wire     [31:0] n13418;
wire     [31:0] n13419;
wire     [31:0] n13420;
wire     [31:0] n13421;
wire     [31:0] n13422;
wire     [31:0] n13423;
wire     [31:0] n13424;
wire     [31:0] n13425;
wire     [31:0] n13426;
wire     [31:0] n13427;
wire     [31:0] n13428;
wire     [31:0] n13429;
wire     [31:0] n13430;
wire     [31:0] n13431;
wire     [31:0] n13432;
wire     [31:0] n13433;
wire     [31:0] n13434;
wire     [31:0] n13435;
wire     [31:0] n13436;
wire     [31:0] n13437;
wire     [31:0] n13438;
wire     [31:0] n13439;
wire     [31:0] n13440;
wire     [31:0] n13441;
wire     [31:0] n13442;
wire     [31:0] n13443;
wire     [31:0] n13444;
wire     [31:0] n13445;
wire     [31:0] n13446;
wire     [31:0] n13447;
wire     [31:0] n13448;
wire     [31:0] n13449;
wire     [31:0] n13450;
wire     [31:0] n13451;
wire     [31:0] n13452;
wire     [31:0] n13453;
wire     [31:0] n13454;
wire     [31:0] n13455;
wire     [31:0] n13456;
wire     [31:0] n13457;
wire     [31:0] n13458;
wire     [31:0] n13459;
wire     [31:0] n13460;
wire     [31:0] n13461;
wire     [31:0] n13462;
wire     [31:0] n13463;
wire     [31:0] n13464;
wire     [31:0] n13465;
wire     [31:0] n13466;
wire     [31:0] n13467;
wire     [31:0] n13468;
wire     [31:0] n13469;
wire     [31:0] n13470;
wire     [31:0] n13471;
wire     [31:0] n13472;
wire     [31:0] n13473;
wire     [31:0] n13474;
wire     [31:0] n13475;
wire     [31:0] n13476;
wire     [31:0] n13477;
wire     [31:0] n13478;
wire     [31:0] n13479;
wire     [31:0] n13480;
wire     [31:0] n13481;
wire     [31:0] n13482;
wire     [31:0] n13483;
wire     [31:0] n13484;
wire     [31:0] n13485;
wire     [31:0] n13486;
wire     [31:0] n13487;
wire     [31:0] n13488;
wire     [31:0] n13489;
wire     [31:0] n13490;
wire     [31:0] n13491;
wire     [31:0] n13492;
wire     [31:0] n13493;
wire     [31:0] n13494;
wire     [31:0] n13495;
wire     [31:0] n13496;
wire     [31:0] n13497;
wire     [31:0] n13498;
wire     [31:0] n13499;
wire     [31:0] n13500;
wire     [31:0] n13501;
wire     [31:0] n13502;
wire     [31:0] n13503;
wire     [31:0] n13504;
wire     [31:0] n13505;
wire     [31:0] n13506;
wire     [31:0] n13507;
wire     [31:0] n13508;
wire     [31:0] n13509;
wire     [31:0] n13510;
wire     [31:0] n13511;
wire     [31:0] n13512;
wire     [31:0] n13513;
wire     [31:0] n13514;
wire     [31:0] n13515;
wire     [31:0] n13516;
wire     [31:0] n13517;
wire     [31:0] n13518;
wire     [31:0] n13519;
wire     [31:0] n13520;
wire     [31:0] n13521;
wire     [31:0] n13522;
wire     [31:0] n13523;
wire     [31:0] n13524;
wire     [31:0] n13525;
wire     [31:0] n13526;
wire     [31:0] n13527;
wire     [31:0] n13528;
wire     [31:0] n13529;
wire     [31:0] n13530;
wire     [31:0] n13531;
wire     [31:0] n13532;
wire     [31:0] n13533;
wire     [31:0] n13534;
wire     [31:0] n13535;
wire     [31:0] n13536;
wire     [31:0] n13537;
wire     [31:0] n13538;
wire     [31:0] n13539;
wire     [31:0] n13540;
wire     [31:0] n13541;
wire     [31:0] n13542;
wire     [31:0] n13543;
wire     [31:0] n13544;
wire     [31:0] n13545;
wire     [31:0] n13546;
wire     [31:0] n13547;
wire     [31:0] n13548;
wire     [31:0] n13549;
wire     [31:0] n13550;
wire     [31:0] n13551;
wire     [31:0] n13552;
wire     [31:0] n13553;
wire     [31:0] n13554;
wire     [31:0] n13555;
wire     [31:0] n13556;
wire     [31:0] n13557;
wire     [31:0] n13558;
wire     [31:0] n13559;
wire     [31:0] n13560;
wire     [31:0] n13561;
wire     [31:0] n13562;
wire     [31:0] n13563;
wire     [31:0] n13564;
wire     [31:0] n13565;
wire     [31:0] n13566;
wire     [31:0] n13567;
wire     [31:0] n13568;
wire     [31:0] n13569;
wire     [31:0] n13570;
wire     [31:0] n13571;
wire     [31:0] n13572;
wire     [31:0] n13573;
wire     [31:0] n13574;
wire     [31:0] n13575;
wire     [31:0] n13576;
wire     [31:0] n13577;
wire     [31:0] n13578;
wire     [31:0] n13579;
wire     [31:0] n13580;
wire     [31:0] n13581;
wire     [31:0] n13582;
wire     [31:0] n13583;
wire     [31:0] n13584;
wire     [31:0] n13585;
wire     [31:0] n13586;
wire     [31:0] n13587;
wire     [31:0] n13588;
wire     [31:0] n13589;
wire     [31:0] n13590;
wire     [31:0] n13591;
wire     [31:0] n13592;
wire     [31:0] n13593;
wire     [31:0] n13594;
wire     [31:0] n13595;
wire     [31:0] n13596;
wire     [31:0] n13597;
wire     [31:0] n13598;
wire     [31:0] n13599;
wire     [31:0] n13600;
wire     [31:0] n13601;
wire     [31:0] n13602;
wire     [31:0] n13603;
wire     [31:0] n13604;
wire     [31:0] n13605;
wire     [31:0] n13606;
wire     [31:0] n13607;
wire     [31:0] n13608;
wire     [31:0] n13609;
wire     [31:0] n13610;
wire     [31:0] n13611;
wire     [31:0] n13612;
wire     [31:0] n13613;
wire     [31:0] n13614;
wire     [31:0] n13615;
wire     [31:0] n13616;
wire     [31:0] n13617;
wire     [31:0] n13618;
wire     [31:0] n13619;
wire     [31:0] n13620;
wire     [31:0] n13621;
wire     [31:0] n13622;
wire     [31:0] n13623;
wire     [31:0] n13624;
wire     [31:0] n13625;
wire     [31:0] n13626;
wire     [31:0] n13627;
wire     [31:0] n13628;
wire            n13629;
wire            n13630;
wire     [31:0] n13631;
wire     [31:0] n13632;
wire     [31:0] n13633;
wire     [31:0] n13634;
wire     [31:0] n13635;
wire     [31:0] n13636;
wire     [31:0] n13637;
wire     [31:0] n13638;
wire     [31:0] n13639;
wire     [31:0] n13640;
wire     [31:0] n13641;
wire     [31:0] n13642;
wire     [31:0] n13643;
wire     [31:0] n13644;
wire     [31:0] n13645;
wire     [31:0] n13646;
wire     [31:0] n13647;
wire     [31:0] n13648;
wire     [31:0] n13649;
wire     [31:0] n13650;
wire     [31:0] n13651;
wire     [31:0] n13652;
wire     [31:0] n13653;
wire     [31:0] n13654;
wire     [31:0] n13655;
wire     [31:0] n13656;
wire     [31:0] n13657;
wire     [31:0] n13658;
wire     [31:0] n13659;
wire     [31:0] n13660;
wire     [31:0] n13661;
wire     [31:0] n13662;
wire     [31:0] n13663;
wire            n13664;
wire            n13665;
wire            n13666;
wire            n13667;
wire            n13668;
wire            n13669;
wire            n13670;
wire            n13671;
wire            n13672;
wire            n13673;
wire            n13674;
wire            n13675;
wire            n13676;
wire            n13677;
wire            n13678;
wire            n13679;
wire            n13680;
wire            n13681;
wire            n13682;
wire            n13683;
wire            n13684;
wire            n13685;
wire            n13686;
wire            n13687;
wire            n13688;
wire            n13689;
wire            n13690;
wire            n13691;
wire            n13692;
wire            n13693;
wire            n13694;
wire            n13695;
wire            n13696;
wire            n13697;
wire            n13698;
wire            n13699;
wire            n13700;
wire            n13701;
wire            n13702;
wire            n13703;
wire            n13704;
wire            n13705;
wire            n13706;
wire            n13707;
wire            n13708;
wire            n13709;
wire            n13710;
wire            n13711;
wire            n13712;
wire            n13713;
wire            n13714;
wire            n13715;
wire            n13716;
wire            n13717;
wire            n13718;
wire            n13719;
wire            n13720;
wire            n13721;
wire            n13722;
wire            n13723;
wire            n13724;
wire            n13725;
wire            n13726;
wire            n13727;
wire            n13728;
wire            n13729;
wire            n13730;
wire            n13731;
wire            n13732;
wire            n13733;
wire            n13734;
wire            n13735;
wire            n13736;
wire            n13737;
wire            n13738;
wire            n13739;
wire            n13740;
wire            n13741;
wire            n13742;
wire            n13743;
wire            n13744;
wire            n13745;
wire            n13746;
wire            n13747;
wire            n13748;
wire            n13749;
wire            n13750;
wire            n13751;
wire            n13752;
wire            n13753;
wire            n13754;
wire            n13755;
wire            n13756;
wire            n13757;
wire            n13758;
wire            n13759;
wire            n13760;
wire            n13761;
wire            n13762;
wire            n13763;
wire            n13764;
wire            n13765;
wire            n13766;
wire            n13767;
wire            n13768;
wire            n13769;
wire            n13770;
wire            n13771;
wire            n13772;
wire            n13773;
wire            n13774;
wire            n13775;
wire            n13776;
wire            n13777;
wire            n13778;
wire            n13779;
wire            n13780;
wire            n13781;
wire            n13782;
wire            n13783;
wire            n13784;
wire            n13785;
wire            n13786;
wire            n13787;
wire            n13788;
wire            n13789;
wire            n13790;
wire            n13791;
wire            n13792;
wire            n13793;
wire            n13794;
wire            n13795;
wire            n13796;
wire            n13797;
wire            n13798;
wire            n13799;
wire            n13800;
wire            n13801;
wire            n13802;
wire            n13803;
wire            n13804;
wire            n13805;
wire            n13806;
wire            n13807;
wire            n13808;
wire            n13809;
wire            n13810;
wire            n13811;
wire            n13812;
wire            n13813;
wire            n13814;
wire            n13815;
wire            n13816;
wire            n13817;
wire            n13818;
wire            n13819;
wire            n13820;
wire            n13821;
wire            n13822;
wire            n13823;
wire            n13824;
wire            n13825;
wire            n13826;
wire            n13827;
wire            n13828;
wire            n13829;
wire            n13830;
wire            n13831;
wire            n13832;
wire            n13833;
wire            n13834;
wire            n13835;
wire            n13836;
wire            n13837;
wire            n13838;
wire            n13839;
wire            n13840;
wire            n13841;
wire            n13842;
wire            n13843;
wire            n13844;
wire            n13845;
wire            n13846;
wire            n13847;
wire            n13848;
wire            n13849;
wire            n13850;
wire            n13851;
wire            n13852;
wire            n13853;
wire            n13854;
wire            n13855;
wire            n13856;
wire            n13857;
wire            n13858;
wire            n13859;
wire            n13860;
wire            n13861;
wire            n13862;
wire            n13863;
wire            n13864;
wire            n13865;
wire            n13866;
wire            n13867;
wire            n13868;
wire            n13869;
wire            n13870;
wire            n13871;
wire            n13872;
wire            n13873;
wire            n13874;
wire            n13875;
wire            n13876;
wire            n13877;
wire            n13878;
wire            n13879;
wire            n13880;
wire            n13881;
wire            n13882;
wire            n13883;
wire            n13884;
wire            n13885;
wire            n13886;
wire            n13887;
wire            n13888;
wire            n13889;
wire            n13890;
wire            n13891;
wire            n13892;
wire            n13893;
wire            n13894;
wire            n13895;
wire            n13896;
wire            n13897;
wire            n13898;
wire            n13899;
wire            n13900;
wire            n13901;
wire            n13902;
wire            n13903;
wire            n13904;
wire            n13905;
wire            n13906;
wire            n13907;
wire            n13908;
wire            n13909;
wire            n13910;
wire            n13911;
wire            n13912;
wire            n13913;
wire            n13914;
wire            n13915;
wire            n13916;
wire            n13917;
wire            n13918;
wire            n13919;
wire            n13920;
wire            n13921;
wire            n13922;
wire            n13923;
wire            n13924;
wire            n13925;
wire            n13926;
wire            n13927;
wire            n13928;
wire            n13929;
wire            n13930;
wire            n13931;
wire            n13932;
wire            n13933;
wire            n13934;
wire            n13935;
wire            n13936;
wire            n13937;
wire            n13938;
wire            n13939;
wire            n13940;
wire            n13941;
wire            n13942;
wire            n13943;
wire            n13944;
wire            n13945;
wire            n13946;
wire            n13947;
wire            n13948;
wire            n13949;
wire            n13950;
wire            n13951;
wire            n13952;
wire            n13953;
wire            n13954;
wire            n13955;
wire            n13956;
wire            n13957;
wire            n13958;
wire            n13959;
wire            n13960;
wire            n13961;
wire            n13962;
wire            n13963;
wire            n13964;
wire            n13965;
wire            n13966;
wire            n13967;
wire            n13968;
wire            n13969;
wire            n13970;
wire            n13971;
wire            n13972;
wire            n13973;
wire            n13974;
wire            n13975;
wire            n13976;
wire            n13977;
wire            n13978;
wire            n13979;
wire            n13980;
wire            n13981;
wire            n13982;
wire            n13983;
wire            n13984;
wire            n13985;
wire            n13986;
wire            n13987;
wire            n13988;
wire            n13989;
wire            n13990;
wire            n13991;
wire            n13992;
wire            n13993;
wire            n13994;
wire            n13995;
wire            n13996;
wire            n13997;
wire            n13998;
wire            n13999;
wire            n14000;
wire            n14001;
wire            n14002;
wire            n14003;
wire            n14004;
wire            n14005;
wire            n14006;
wire            n14007;
wire            n14008;
wire            n14009;
wire            n14010;
wire            n14011;
wire            n14012;
wire            n14013;
wire            n14014;
wire            n14015;
wire            n14016;
wire            n14017;
wire            n14018;
wire            n14019;
wire            n14020;
wire            n14021;
wire            n14022;
wire            n14023;
wire            n14024;
wire            n14025;
wire            n14026;
wire            n14027;
wire            n14028;
wire            n14029;
wire            n14030;
wire            n14031;
wire            n14032;
wire            n14033;
wire            n14034;
wire            n14035;
wire            n14036;
wire            n14037;
wire            n14038;
wire            n14039;
wire            n14040;
wire            n14041;
wire            n14042;
wire            n14043;
wire            n14044;
wire            n14045;
wire            n14046;
wire            n14047;
wire            n14048;
wire            n14049;
wire            n14050;
wire            n14051;
wire            n14052;
wire            n14053;
wire            n14054;
wire            n14055;
wire            n14056;
wire            n14057;
wire            n14058;
wire            n14059;
wire            n14060;
wire            n14061;
wire            n14062;
wire            n14063;
wire            n14064;
wire            n14065;
wire            n14066;
wire            n14067;
wire            n14068;
wire            n14069;
wire            n14070;
wire            n14071;
wire            n14072;
wire            n14073;
wire            n14074;
wire            n14075;
wire            n14076;
wire            n14077;
wire            n14078;
wire            n14079;
wire            n14080;
wire            n14081;
wire            n14082;
wire            n14083;
wire            n14084;
wire            n14085;
wire            n14086;
wire            n14087;
wire            n14088;
wire            n14089;
wire            n14090;
wire            n14091;
wire            n14092;
wire            n14093;
wire            n14094;
wire            n14095;
wire            n14096;
wire            n14097;
wire            n14098;
wire            n14099;
wire            n14100;
wire            n14101;
wire            n14102;
wire            n14103;
wire            n14104;
wire            n14105;
wire            n14106;
wire            n14107;
wire            n14108;
wire            n14109;
wire            n14110;
wire            n14111;
wire            n14112;
wire            n14113;
wire            n14114;
wire            n14115;
wire            n14116;
wire            n14117;
wire            n14118;
wire            n14119;
wire            n14120;
wire            n14121;
wire            n14122;
wire            n14123;
wire            n14124;
wire            n14125;
wire            n14126;
wire            n14127;
wire            n14128;
wire            n14129;
wire            n14130;
wire            n14131;
wire            n14132;
wire            n14133;
wire            n14134;
wire            n14135;
wire            n14136;
wire            n14137;
wire            n14138;
wire            n14139;
wire            n14140;
wire            n14141;
wire            n14142;
wire            n14143;
wire            n14144;
wire            n14145;
wire            n14146;
wire            n14147;
wire            n14148;
wire            n14149;
wire            n14150;
wire            n14151;
wire            n14152;
wire            n14153;
wire            n14154;
wire            n14155;
wire            n14156;
wire            n14157;
wire            n14158;
wire            n14159;
wire            n14160;
wire            n14161;
wire            n14162;
wire            n14163;
wire            n14164;
wire            n14165;
wire            n14166;
wire            n14167;
wire            n14168;
wire            n14169;
wire            n14170;
wire            n14171;
wire            n14172;
wire            n14173;
wire            n14174;
wire            n14175;
wire            n14176;
wire            n14177;
wire            n14178;
wire            n14179;
wire            n14180;
wire            n14181;
wire            n14182;
wire            n14183;
wire            n14184;
wire            n14185;
wire            n14186;
wire            n14187;
wire            n14188;
wire            n14189;
wire            n14190;
wire            n14191;
wire     [31:0] n14192;
wire     [31:0] n14193;
wire     [31:0] n14194;
wire     [31:0] n14195;
wire     [31:0] n14196;
wire     [31:0] n14197;
wire     [31:0] n14198;
wire     [31:0] n14199;
wire     [31:0] n14200;
wire     [31:0] n14201;
wire     [31:0] n14202;
wire     [31:0] n14203;
wire     [31:0] n14204;
wire     [31:0] n14205;
wire     [31:0] n14206;
wire     [31:0] n14207;
wire     [31:0] n14208;
wire     [31:0] n14209;
wire     [31:0] n14210;
wire     [31:0] n14211;
wire     [31:0] n14212;
wire     [31:0] n14213;
wire     [31:0] n14214;
wire     [31:0] n14215;
wire     [31:0] n14216;
wire     [31:0] n14217;
wire     [31:0] n14218;
wire     [31:0] n14219;
wire     [31:0] n14220;
wire     [31:0] n14221;
wire     [31:0] n14222;
wire     [31:0] n14223;
wire     [31:0] n14224;
wire     [31:0] n14225;
wire     [31:0] n14226;
wire     [31:0] n14227;
wire     [31:0] n14228;
wire     [31:0] n14229;
wire     [31:0] n14230;
wire     [31:0] n14231;
wire     [31:0] n14232;
wire     [31:0] n14233;
wire     [31:0] n14234;
wire     [31:0] n14235;
wire     [31:0] n14236;
wire     [31:0] n14237;
wire     [31:0] n14238;
wire     [31:0] n14239;
wire     [31:0] n14240;
wire     [31:0] n14241;
wire     [31:0] n14242;
wire     [31:0] n14243;
wire     [31:0] n14244;
wire     [31:0] n14245;
wire     [31:0] n14246;
wire     [31:0] n14247;
wire     [31:0] n14248;
wire     [31:0] n14249;
wire     [31:0] n14250;
wire     [31:0] n14251;
wire     [31:0] n14252;
wire     [31:0] n14253;
wire     [31:0] n14254;
wire     [31:0] n14255;
wire     [31:0] n14256;
wire     [31:0] n14257;
wire     [31:0] n14258;
wire     [31:0] n14259;
wire     [31:0] n14260;
wire     [31:0] n14261;
wire     [31:0] n14262;
wire     [31:0] n14263;
wire     [31:0] n14264;
wire     [31:0] n14265;
wire     [31:0] n14266;
wire     [31:0] n14267;
wire     [31:0] n14268;
wire     [31:0] n14269;
wire     [31:0] n14270;
wire     [31:0] n14271;
wire     [31:0] n14272;
wire     [31:0] n14273;
wire     [31:0] n14274;
wire     [31:0] n14275;
wire     [31:0] n14276;
wire     [31:0] n14277;
wire     [31:0] n14278;
wire     [31:0] n14279;
wire     [31:0] n14280;
wire     [31:0] n14281;
wire     [31:0] n14282;
wire     [31:0] n14283;
wire     [31:0] n14284;
wire     [31:0] n14285;
wire     [31:0] n14286;
wire     [31:0] n14287;
wire     [31:0] n14288;
wire     [31:0] n14289;
wire     [31:0] n14290;
wire     [31:0] n14291;
wire     [31:0] n14292;
wire     [31:0] n14293;
wire     [31:0] n14294;
wire     [31:0] n14295;
wire     [31:0] n14296;
wire     [31:0] n14297;
wire     [31:0] n14298;
wire     [31:0] n14299;
wire     [31:0] n14300;
wire     [31:0] n14301;
wire     [31:0] n14302;
wire     [31:0] n14303;
wire     [31:0] n14304;
wire     [31:0] n14305;
wire     [31:0] n14306;
wire     [31:0] n14307;
wire     [31:0] n14308;
wire     [31:0] n14309;
wire     [31:0] n14310;
wire     [31:0] n14311;
wire     [31:0] n14312;
wire     [31:0] n14313;
wire     [31:0] n14314;
wire     [31:0] n14315;
wire     [31:0] n14316;
wire     [31:0] n14317;
wire     [31:0] n14318;
wire     [31:0] n14319;
wire     [31:0] n14320;
wire     [31:0] n14321;
wire     [31:0] n14322;
wire     [31:0] n14323;
wire     [31:0] n14324;
wire     [31:0] n14325;
wire     [31:0] n14326;
wire     [31:0] n14327;
wire     [31:0] n14328;
wire     [31:0] n14329;
wire     [31:0] n14330;
wire     [31:0] n14331;
wire     [31:0] n14332;
wire     [31:0] n14333;
wire     [31:0] n14334;
wire     [31:0] n14335;
wire     [31:0] n14336;
wire     [31:0] n14337;
wire     [31:0] n14338;
wire     [31:0] n14339;
wire     [31:0] n14340;
wire     [31:0] n14341;
wire     [31:0] n14342;
wire     [31:0] n14343;
wire     [31:0] n14344;
wire     [31:0] n14345;
wire     [31:0] n14346;
wire     [31:0] n14347;
wire     [31:0] n14348;
wire     [31:0] n14349;
wire     [31:0] n14350;
wire     [31:0] n14351;
wire     [31:0] n14352;
wire     [31:0] n14353;
wire     [31:0] n14354;
wire     [31:0] n14355;
wire     [31:0] n14356;
wire     [31:0] n14357;
wire     [31:0] n14358;
wire     [31:0] n14359;
wire     [31:0] n14360;
wire     [31:0] n14361;
wire     [31:0] n14362;
wire     [31:0] n14363;
wire     [31:0] n14364;
wire     [31:0] n14365;
wire     [31:0] n14366;
wire     [31:0] n14367;
wire     [31:0] n14368;
wire     [31:0] n14369;
wire     [31:0] n14370;
wire     [31:0] n14371;
wire     [31:0] n14372;
wire     [31:0] n14373;
wire     [31:0] n14374;
wire     [31:0] n14375;
wire     [31:0] n14376;
wire     [31:0] n14377;
wire     [31:0] n14378;
wire     [31:0] n14379;
wire     [31:0] n14380;
wire     [31:0] n14381;
wire     [31:0] n14382;
wire     [31:0] n14383;
wire     [31:0] n14384;
wire     [31:0] n14385;
wire     [31:0] n14386;
wire     [31:0] n14387;
wire     [31:0] n14388;
wire     [31:0] n14389;
wire     [31:0] n14390;
wire     [31:0] n14391;
wire     [31:0] n14392;
wire     [31:0] n14393;
wire     [31:0] n14394;
wire     [31:0] n14395;
wire     [31:0] n14396;
wire     [31:0] n14397;
wire     [31:0] n14398;
wire     [31:0] n14399;
wire     [31:0] n14400;
wire     [31:0] n14401;
wire     [31:0] n14402;
wire     [31:0] n14403;
wire     [31:0] n14404;
wire     [31:0] n14405;
wire     [31:0] n14406;
wire     [31:0] n14407;
wire     [31:0] n14408;
wire     [31:0] n14409;
wire     [31:0] n14410;
wire     [31:0] n14411;
wire     [31:0] n14412;
wire     [31:0] n14413;
wire     [31:0] n14414;
wire     [31:0] n14415;
wire     [31:0] n14416;
wire     [31:0] n14417;
wire     [31:0] n14418;
wire     [31:0] n14419;
wire     [31:0] n14420;
wire     [31:0] n14421;
wire     [31:0] n14422;
wire     [31:0] n14423;
wire     [31:0] n14424;
wire     [31:0] n14425;
wire     [31:0] n14426;
wire     [31:0] n14427;
wire     [31:0] n14428;
wire     [31:0] n14429;
wire     [31:0] n14430;
wire     [31:0] n14431;
wire     [31:0] n14432;
wire     [31:0] n14433;
wire     [31:0] n14434;
wire     [31:0] n14435;
wire     [31:0] n14436;
wire     [31:0] n14437;
wire     [31:0] n14438;
wire     [31:0] n14439;
wire     [31:0] n14440;
wire     [31:0] n14441;
wire     [31:0] n14442;
wire     [31:0] n14443;
wire     [31:0] n14444;
wire     [31:0] n14445;
wire     [31:0] n14446;
wire     [31:0] n14447;
wire     [31:0] n14448;
wire     [31:0] n14449;
wire     [31:0] n14450;
wire     [31:0] n14451;
wire     [31:0] n14452;
wire     [31:0] n14453;
wire     [31:0] n14454;
wire     [31:0] n14455;
wire     [31:0] n14456;
wire     [31:0] n14457;
wire     [31:0] n14458;
wire     [31:0] n14459;
wire     [31:0] n14460;
wire     [31:0] n14461;
wire     [31:0] n14462;
wire     [31:0] n14463;
wire     [31:0] n14464;
wire     [31:0] n14465;
wire     [31:0] n14466;
wire     [31:0] n14467;
wire     [31:0] n14468;
wire     [31:0] n14469;
wire     [31:0] n14470;
wire     [31:0] n14471;
wire     [31:0] n14472;
wire     [31:0] n14473;
wire     [31:0] n14474;
wire     [31:0] n14475;
wire     [31:0] n14476;
wire     [31:0] n14477;
wire     [31:0] n14478;
wire     [31:0] n14479;
wire     [31:0] n14480;
wire     [31:0] n14481;
wire     [31:0] n14482;
wire     [31:0] n14483;
wire     [31:0] n14484;
wire     [31:0] n14485;
wire     [31:0] n14486;
wire     [31:0] n14487;
wire     [31:0] n14488;
wire     [31:0] n14489;
wire     [31:0] n14490;
wire     [31:0] n14491;
wire     [31:0] n14492;
wire     [31:0] n14493;
wire     [31:0] n14494;
wire     [31:0] n14495;
wire     [31:0] n14496;
wire     [31:0] n14497;
wire     [31:0] n14498;
wire     [31:0] n14499;
wire     [31:0] n14500;
wire     [31:0] n14501;
wire     [31:0] n14502;
wire     [31:0] n14503;
wire     [31:0] n14504;
wire     [31:0] n14505;
wire     [31:0] n14506;
wire     [31:0] n14507;
wire     [31:0] n14508;
wire     [31:0] n14509;
wire     [31:0] n14510;
wire     [31:0] n14511;
wire     [31:0] n14512;
wire     [31:0] n14513;
wire     [31:0] n14514;
wire     [31:0] n14515;
wire     [31:0] n14516;
wire     [31:0] n14517;
wire     [31:0] n14518;
wire     [31:0] n14519;
wire     [31:0] n14520;
wire     [31:0] n14521;
wire     [31:0] n14522;
wire     [31:0] n14523;
wire     [31:0] n14524;
wire     [31:0] n14525;
wire     [31:0] n14526;
wire     [31:0] n14527;
wire     [31:0] n14528;
wire     [31:0] n14529;
wire     [31:0] n14530;
wire     [31:0] n14531;
wire     [31:0] n14532;
wire     [31:0] n14533;
wire     [31:0] n14534;
wire     [31:0] n14535;
wire     [31:0] n14536;
wire     [31:0] n14537;
wire     [31:0] n14538;
wire     [31:0] n14539;
wire     [31:0] n14540;
wire     [31:0] n14541;
wire     [31:0] n14542;
wire     [31:0] n14543;
wire     [31:0] n14544;
wire     [31:0] n14545;
wire     [31:0] n14546;
wire     [31:0] n14547;
wire     [31:0] n14548;
wire     [31:0] n14549;
wire     [31:0] n14550;
wire     [31:0] n14551;
wire     [31:0] n14552;
wire     [31:0] n14553;
wire     [31:0] n14554;
wire     [31:0] n14555;
wire     [31:0] n14556;
wire     [31:0] n14557;
wire     [31:0] n14558;
wire     [31:0] n14559;
wire     [31:0] n14560;
wire     [31:0] n14561;
wire     [31:0] n14562;
wire     [31:0] n14563;
wire     [31:0] n14564;
wire     [31:0] n14565;
wire     [31:0] n14566;
wire     [31:0] n14567;
wire     [31:0] n14568;
wire     [31:0] n14569;
wire     [31:0] n14570;
wire     [31:0] n14571;
wire     [31:0] n14572;
wire     [31:0] n14573;
wire     [31:0] n14574;
wire     [31:0] n14575;
wire     [31:0] n14576;
wire     [31:0] n14577;
wire     [31:0] n14578;
wire     [31:0] n14579;
wire     [31:0] n14580;
wire     [31:0] n14581;
wire     [31:0] n14582;
wire     [31:0] n14583;
wire     [31:0] n14584;
wire     [31:0] n14585;
wire     [31:0] n14586;
wire     [31:0] n14587;
wire     [31:0] n14588;
wire     [31:0] n14589;
wire     [31:0] n14590;
wire     [31:0] n14591;
wire     [31:0] n14592;
wire     [31:0] n14593;
wire     [31:0] n14594;
wire     [31:0] n14595;
wire     [31:0] n14596;
wire     [31:0] n14597;
wire     [31:0] n14598;
wire     [31:0] n14599;
wire     [31:0] n14600;
wire     [31:0] n14601;
wire     [31:0] n14602;
wire     [31:0] n14603;
wire     [31:0] n14604;
wire     [31:0] n14605;
wire     [31:0] n14606;
wire     [31:0] n14607;
wire     [31:0] n14608;
wire     [31:0] n14609;
wire     [31:0] n14610;
wire     [31:0] n14611;
wire     [31:0] n14612;
wire     [31:0] n14613;
wire     [31:0] n14614;
wire     [31:0] n14615;
wire     [31:0] n14616;
wire     [31:0] n14617;
wire     [31:0] n14618;
wire     [31:0] n14619;
wire     [31:0] n14620;
wire     [31:0] n14621;
wire     [31:0] n14622;
wire     [31:0] n14623;
wire     [31:0] n14624;
wire     [31:0] n14625;
wire     [31:0] n14626;
wire     [31:0] n14627;
wire     [31:0] n14628;
wire     [31:0] n14629;
wire     [31:0] n14630;
wire     [31:0] n14631;
wire     [31:0] n14632;
wire     [31:0] n14633;
wire     [31:0] n14634;
wire     [31:0] n14635;
wire     [31:0] n14636;
wire     [31:0] n14637;
wire     [31:0] n14638;
wire     [31:0] n14639;
wire     [31:0] n14640;
wire     [31:0] n14641;
wire     [31:0] n14642;
wire     [31:0] n14643;
wire     [31:0] n14644;
wire     [31:0] n14645;
wire     [31:0] n14646;
wire     [31:0] n14647;
wire     [31:0] n14648;
wire     [31:0] n14649;
wire     [31:0] n14650;
wire     [31:0] n14651;
wire     [31:0] n14652;
wire     [31:0] n14653;
wire     [31:0] n14654;
wire     [31:0] n14655;
wire     [31:0] n14656;
wire     [31:0] n14657;
wire     [31:0] n14658;
wire     [31:0] n14659;
wire     [31:0] n14660;
wire     [31:0] n14661;
wire     [31:0] n14662;
wire     [31:0] n14663;
wire     [31:0] n14664;
wire     [31:0] n14665;
wire     [31:0] n14666;
wire     [31:0] n14667;
wire     [31:0] n14668;
wire     [31:0] n14669;
wire     [31:0] n14670;
wire     [31:0] n14671;
wire     [31:0] n14672;
wire     [31:0] n14673;
wire     [31:0] n14674;
wire     [31:0] n14675;
wire     [31:0] n14676;
wire     [31:0] n14677;
wire     [31:0] n14678;
wire     [31:0] n14679;
wire     [31:0] n14680;
wire     [31:0] n14681;
wire     [31:0] n14682;
wire     [31:0] n14683;
wire     [31:0] n14684;
wire     [31:0] n14685;
wire     [31:0] n14686;
wire     [31:0] n14687;
wire     [31:0] n14688;
wire     [31:0] n14689;
wire     [31:0] n14690;
wire     [31:0] n14691;
wire     [31:0] n14692;
wire     [31:0] n14693;
wire     [31:0] n14694;
wire     [31:0] n14695;
wire     [31:0] n14696;
wire     [31:0] n14697;
wire     [31:0] n14698;
wire     [31:0] n14699;
wire     [31:0] n14700;
wire     [31:0] n14701;
wire     [31:0] n14702;
wire     [31:0] n14703;
wire     [31:0] n14704;
wire     [31:0] n14705;
wire     [31:0] n14706;
wire     [31:0] n14707;
wire     [31:0] n14708;
wire     [31:0] n14709;
wire     [31:0] n14710;
wire     [31:0] n14711;
wire     [31:0] n14712;
wire     [31:0] n14713;
wire            n14714;
wire            n14715;
wire            n14716;
wire            n14717;
wire            n14718;
wire            n14719;
wire            n14720;
wire            n14721;
wire            n14722;
wire            n14723;
wire            n14724;
wire            n14725;
wire            n14726;
wire            n14727;
wire            n14728;
wire            n14729;
wire            n14730;
wire            n14731;
wire            n14732;
wire            n14733;
wire            n14734;
wire            n14735;
wire            n14736;
wire            n14737;
wire            n14738;
wire            n14739;
wire            n14740;
wire            n14741;
wire            n14742;
wire            n14743;
wire            n14744;
wire            n14745;
wire            n14746;
wire            n14747;
wire            n14748;
wire            n14749;
wire            n14750;
wire            n14751;
wire            n14752;
wire            n14753;
wire            n14754;
wire            n14755;
wire            n14756;
wire            n14757;
wire            n14758;
wire            n14759;
wire            n14760;
wire            n14761;
wire            n14762;
wire            n14763;
wire            n14764;
wire            n14765;
wire            n14766;
wire            n14767;
wire            n14768;
wire            n14769;
wire            n14770;
wire            n14771;
wire            n14772;
wire            n14773;
wire            n14774;
wire            n14775;
wire            n14776;
wire            n14777;
wire            n14778;
wire            n14779;
wire            n14780;
wire            n14781;
wire            n14782;
wire            n14783;
wire            n14784;
wire            n14785;
wire            n14786;
wire            n14787;
wire            n14788;
wire            n14789;
wire            n14790;
wire            n14791;
wire            n14792;
wire            n14793;
wire            n14794;
wire            n14795;
wire            n14796;
wire            n14797;
wire            n14798;
wire            n14799;
wire            n14800;
wire            n14801;
wire            n14802;
wire            n14803;
wire            n14804;
wire            n14805;
wire            n14806;
wire            n14807;
wire            n14808;
wire            n14809;
wire            n14810;
wire            n14811;
wire            n14812;
wire            n14813;
wire            n14814;
wire            n14815;
wire            n14816;
wire            n14817;
wire            n14818;
wire            n14819;
wire            n14820;
wire            n14821;
wire            n14822;
wire            n14823;
wire            n14824;
wire            n14825;
wire            n14826;
wire            n14827;
wire            n14828;
wire            n14829;
wire            n14830;
wire            n14831;
wire            n14832;
wire            n14833;
wire            n14834;
wire            n14835;
wire            n14836;
wire            n14837;
wire            n14838;
wire            n14839;
wire            n14840;
wire            n14841;
wire            n14842;
wire            n14843;
wire            n14844;
wire            n14845;
wire            n14846;
wire            n14847;
wire            n14848;
wire            n14849;
wire            n14850;
wire            n14851;
wire            n14852;
wire            n14853;
wire            n14854;
wire            n14855;
wire            n14856;
wire            n14857;
wire            n14858;
wire            n14859;
wire            n14860;
wire            n14861;
wire            n14862;
wire            n14863;
wire            n14864;
wire            n14865;
wire            n14866;
wire            n14867;
wire            n14868;
wire            n14869;
wire            n14870;
wire            n14871;
wire            n14872;
wire            n14873;
wire            n14874;
wire            n14875;
wire            n14876;
wire            n14877;
wire            n14878;
wire            n14879;
wire            n14880;
wire            n14881;
wire            n14882;
wire            n14883;
wire            n14884;
wire            n14885;
wire            n14886;
wire            n14887;
wire            n14888;
wire            n14889;
wire            n14890;
wire            n14891;
wire            n14892;
wire            n14893;
wire            n14894;
wire            n14895;
wire            n14896;
wire            n14897;
wire            n14898;
wire            n14899;
wire            n14900;
wire            n14901;
wire            n14902;
wire            n14903;
wire            n14904;
wire            n14905;
wire            n14906;
wire            n14907;
wire            n14908;
wire            n14909;
wire            n14910;
wire            n14911;
wire            n14912;
wire            n14913;
wire            n14914;
wire            n14915;
wire            n14916;
wire            n14917;
wire            n14918;
wire            n14919;
wire            n14920;
wire            n14921;
wire            n14922;
wire            n14923;
wire            n14924;
wire            n14925;
wire            n14926;
wire            n14927;
wire            n14928;
wire            n14929;
wire            n14930;
wire            n14931;
wire            n14932;
wire            n14933;
wire            n14934;
wire            n14935;
wire            n14936;
wire            n14937;
wire            n14938;
wire            n14939;
wire            n14940;
wire            n14941;
wire            n14942;
wire            n14943;
wire            n14944;
wire            n14945;
wire            n14946;
wire            n14947;
wire            n14948;
wire            n14949;
wire            n14950;
wire            n14951;
wire            n14952;
wire            n14953;
wire            n14954;
wire            n14955;
wire            n14956;
wire            n14957;
wire            n14958;
wire            n14959;
wire            n14960;
wire            n14961;
wire            n14962;
wire            n14963;
wire            n14964;
wire            n14965;
wire            n14966;
wire            n14967;
wire            n14968;
wire            n14969;
wire            n14970;
wire            n14971;
wire            n14972;
wire            n14973;
wire            n14974;
wire            n14975;
wire            n14976;
wire            n14977;
wire            n14978;
wire            n14979;
wire            n14980;
wire            n14981;
wire            n14982;
wire            n14983;
wire            n14984;
wire            n14985;
wire            n14986;
wire            n14987;
wire            n14988;
wire            n14989;
wire            n14990;
wire            n14991;
wire            n14992;
wire            n14993;
wire            n14994;
wire            n14995;
wire            n14996;
wire            n14997;
wire            n14998;
wire            n14999;
wire            n15000;
wire            n15001;
wire            n15002;
wire            n15003;
wire            n15004;
wire            n15005;
wire            n15006;
wire            n15007;
wire            n15008;
wire            n15009;
wire            n15010;
wire            n15011;
wire            n15012;
wire            n15013;
wire            n15014;
wire            n15015;
wire            n15016;
wire            n15017;
wire            n15018;
wire            n15019;
wire            n15020;
wire            n15021;
wire            n15022;
wire            n15023;
wire            n15024;
wire            n15025;
wire            n15026;
wire            n15027;
wire            n15028;
wire            n15029;
wire            n15030;
wire            n15031;
wire            n15032;
wire            n15033;
wire            n15034;
wire            n15035;
wire            n15036;
wire            n15037;
wire            n15038;
wire            n15039;
wire            n15040;
wire            n15041;
wire            n15042;
wire            n15043;
wire            n15044;
wire            n15045;
wire            n15046;
wire            n15047;
wire            n15048;
wire            n15049;
wire            n15050;
wire            n15051;
wire            n15052;
wire            n15053;
wire            n15054;
wire            n15055;
wire            n15056;
wire            n15057;
wire            n15058;
wire            n15059;
wire            n15060;
wire            n15061;
wire            n15062;
wire            n15063;
wire            n15064;
wire            n15065;
wire            n15066;
wire            n15067;
wire            n15068;
wire            n15069;
wire            n15070;
wire            n15071;
wire            n15072;
wire            n15073;
wire            n15074;
wire            n15075;
wire            n15076;
wire            n15077;
wire            n15078;
wire            n15079;
wire            n15080;
wire            n15081;
wire            n15082;
wire            n15083;
wire            n15084;
wire            n15085;
wire            n15086;
wire            n15087;
wire            n15088;
wire            n15089;
wire            n15090;
wire            n15091;
wire            n15092;
wire            n15093;
wire            n15094;
wire            n15095;
wire            n15096;
wire            n15097;
wire            n15098;
wire            n15099;
wire            n15100;
wire            n15101;
wire            n15102;
wire            n15103;
wire            n15104;
wire            n15105;
wire            n15106;
wire            n15107;
wire            n15108;
wire            n15109;
wire            n15110;
wire            n15111;
wire            n15112;
wire            n15113;
wire            n15114;
wire            n15115;
wire            n15116;
wire            n15117;
wire            n15118;
wire            n15119;
wire            n15120;
wire            n15121;
wire            n15122;
wire            n15123;
wire            n15124;
wire            n15125;
wire            n15126;
wire            n15127;
wire            n15128;
wire            n15129;
wire            n15130;
wire            n15131;
wire            n15132;
wire            n15133;
wire            n15134;
wire            n15135;
wire            n15136;
wire            n15137;
wire            n15138;
wire            n15139;
wire            n15140;
wire            n15141;
wire            n15142;
wire            n15143;
wire            n15144;
wire            n15145;
wire            n15146;
wire            n15147;
wire            n15148;
wire            n15149;
wire            n15150;
wire            n15151;
wire            n15152;
wire            n15153;
wire            n15154;
wire            n15155;
wire            n15156;
wire            n15157;
wire            n15158;
wire            n15159;
wire            n15160;
wire            n15161;
wire            n15162;
wire            n15163;
wire            n15164;
wire            n15165;
wire            n15166;
wire            n15167;
wire            n15168;
wire            n15169;
wire            n15170;
wire            n15171;
wire            n15172;
wire            n15173;
wire            n15174;
wire            n15175;
wire            n15176;
wire            n15177;
wire            n15178;
wire            n15179;
wire            n15180;
wire            n15181;
wire            n15182;
wire            n15183;
wire            n15184;
wire            n15185;
wire            n15186;
wire            n15187;
wire            n15188;
wire            n15189;
wire            n15190;
wire            n15191;
wire            n15192;
wire            n15193;
wire            n15194;
wire            n15195;
wire            n15196;
wire            n15197;
wire            n15198;
wire            n15199;
wire            n15200;
wire            n15201;
wire            n15202;
wire            n15203;
wire            n15204;
wire            n15205;
wire            n15206;
wire            n15207;
wire            n15208;
wire            n15209;
wire            n15210;
wire            n15211;
wire            n15212;
wire            n15213;
wire            n15214;
wire            n15215;
wire            n15216;
wire            n15217;
wire            n15218;
wire            n15219;
wire            n15220;
wire            n15221;
wire            n15222;
wire            n15223;
wire            n15224;
wire            n15225;
wire     [31:0] n15226;
wire     [31:0] n15227;
wire     [31:0] n15228;
wire     [31:0] n15229;
wire     [31:0] n15230;
wire     [31:0] n15231;
wire     [31:0] n15232;
wire     [31:0] n15233;
wire     [31:0] n15234;
wire     [31:0] n15235;
wire     [31:0] n15236;
wire     [31:0] n15237;
wire     [31:0] n15238;
wire     [31:0] n15239;
wire     [31:0] n15240;
wire     [31:0] n15241;
wire     [31:0] n15242;
wire     [31:0] n15243;
wire     [31:0] n15244;
wire     [31:0] n15245;
wire     [31:0] n15246;
wire     [31:0] n15247;
wire     [31:0] n15248;
wire     [31:0] n15249;
wire     [31:0] n15250;
wire     [31:0] n15251;
wire     [31:0] n15252;
wire     [31:0] n15253;
wire     [31:0] n15254;
wire     [31:0] n15255;
wire     [31:0] n15256;
wire     [31:0] n15257;
wire     [31:0] n15258;
wire     [31:0] n15259;
wire     [31:0] n15260;
wire     [31:0] n15261;
wire     [31:0] n15262;
wire     [31:0] n15263;
wire     [31:0] n15264;
wire     [31:0] n15265;
wire     [31:0] n15266;
wire     [31:0] n15267;
wire     [31:0] n15268;
wire     [31:0] n15269;
wire     [31:0] n15270;
wire     [31:0] n15271;
wire     [31:0] n15272;
wire     [31:0] n15273;
wire     [31:0] n15274;
wire     [31:0] n15275;
wire     [31:0] n15276;
wire     [31:0] n15277;
wire     [31:0] n15278;
wire     [31:0] n15279;
wire     [31:0] n15280;
wire     [31:0] n15281;
wire     [31:0] n15282;
wire     [31:0] n15283;
wire     [31:0] n15284;
wire     [31:0] n15285;
wire     [31:0] n15286;
wire     [31:0] n15287;
wire     [31:0] n15288;
wire     [31:0] n15289;
wire     [31:0] n15290;
wire     [31:0] n15291;
wire     [31:0] n15292;
wire     [31:0] n15293;
wire     [31:0] n15294;
wire     [31:0] n15295;
wire     [31:0] n15296;
wire     [31:0] n15297;
wire     [31:0] n15298;
wire     [31:0] n15299;
wire     [31:0] n15300;
wire     [31:0] n15301;
wire     [31:0] n15302;
wire     [31:0] n15303;
wire     [31:0] n15304;
wire     [31:0] n15305;
wire     [31:0] n15306;
wire     [31:0] n15307;
wire     [31:0] n15308;
wire     [31:0] n15309;
wire     [31:0] n15310;
wire     [31:0] n15311;
wire     [31:0] n15312;
wire     [31:0] n15313;
wire     [31:0] n15314;
wire     [31:0] n15315;
wire     [31:0] n15316;
wire     [31:0] n15317;
wire     [31:0] n15318;
wire     [31:0] n15319;
wire     [31:0] n15320;
wire     [31:0] n15321;
wire     [31:0] n15322;
wire     [31:0] n15323;
wire     [31:0] n15324;
wire     [31:0] n15325;
wire     [31:0] n15326;
wire     [31:0] n15327;
wire     [31:0] n15328;
wire     [31:0] n15329;
wire     [31:0] n15330;
wire     [31:0] n15331;
wire     [31:0] n15332;
wire     [31:0] n15333;
wire     [31:0] n15334;
wire     [31:0] n15335;
wire     [31:0] n15336;
wire     [31:0] n15337;
wire     [31:0] n15338;
wire     [31:0] n15339;
wire     [31:0] n15340;
wire     [31:0] n15341;
wire     [31:0] n15342;
wire     [31:0] n15343;
wire     [31:0] n15344;
wire     [31:0] n15345;
wire     [31:0] n15346;
wire     [31:0] n15347;
wire     [31:0] n15348;
wire     [31:0] n15349;
wire     [31:0] n15350;
wire     [31:0] n15351;
wire     [31:0] n15352;
wire     [31:0] n15353;
wire     [31:0] n15354;
wire     [31:0] n15355;
wire     [31:0] n15356;
wire     [31:0] n15357;
wire     [31:0] n15358;
wire     [31:0] n15359;
wire     [31:0] n15360;
wire     [31:0] n15361;
wire     [31:0] n15362;
wire     [31:0] n15363;
wire     [31:0] n15364;
wire     [31:0] n15365;
wire     [31:0] n15366;
wire     [31:0] n15367;
wire     [31:0] n15368;
wire     [31:0] n15369;
wire     [31:0] n15370;
wire     [31:0] n15371;
wire     [31:0] n15372;
wire     [31:0] n15373;
wire     [31:0] n15374;
wire     [31:0] n15375;
wire     [31:0] n15376;
wire     [31:0] n15377;
wire     [31:0] n15378;
wire     [31:0] n15379;
wire     [31:0] n15380;
wire     [31:0] n15381;
wire     [31:0] n15382;
wire     [31:0] n15383;
wire     [31:0] n15384;
wire     [31:0] n15385;
wire     [31:0] n15386;
wire     [31:0] n15387;
wire     [31:0] n15388;
wire     [31:0] n15389;
wire     [31:0] n15390;
wire     [31:0] n15391;
wire     [31:0] n15392;
wire     [31:0] n15393;
wire     [31:0] n15394;
wire     [31:0] n15395;
wire     [31:0] n15396;
wire     [31:0] n15397;
wire     [31:0] n15398;
wire     [31:0] n15399;
wire     [31:0] n15400;
wire     [31:0] n15401;
wire     [31:0] n15402;
wire     [31:0] n15403;
wire     [31:0] n15404;
wire     [31:0] n15405;
wire     [31:0] n15406;
wire     [31:0] n15407;
wire     [31:0] n15408;
wire     [31:0] n15409;
wire     [31:0] n15410;
wire     [31:0] n15411;
wire     [31:0] n15412;
wire     [31:0] n15413;
wire     [31:0] n15414;
wire     [31:0] n15415;
wire     [31:0] n15416;
wire     [31:0] n15417;
wire     [31:0] n15418;
wire     [31:0] n15419;
wire     [31:0] n15420;
wire     [31:0] n15421;
wire     [31:0] n15422;
wire     [31:0] n15423;
wire     [31:0] n15424;
wire     [31:0] n15425;
wire     [31:0] n15426;
wire     [31:0] n15427;
wire     [31:0] n15428;
wire     [31:0] n15429;
wire     [31:0] n15430;
wire     [31:0] n15431;
wire     [31:0] n15432;
wire     [31:0] n15433;
wire     [31:0] n15434;
wire     [31:0] n15435;
wire     [31:0] n15436;
wire     [31:0] n15437;
wire     [31:0] n15438;
wire     [31:0] n15439;
wire     [31:0] n15440;
wire     [31:0] n15441;
wire     [31:0] n15442;
wire     [31:0] n15443;
wire     [31:0] n15444;
wire     [31:0] n15445;
wire     [31:0] n15446;
wire     [31:0] n15447;
wire     [31:0] n15448;
wire     [31:0] n15449;
wire     [31:0] n15450;
wire     [31:0] n15451;
wire     [31:0] n15452;
wire     [31:0] n15453;
wire     [31:0] n15454;
wire     [31:0] n15455;
wire     [31:0] n15456;
wire     [31:0] n15457;
wire     [31:0] n15458;
wire     [31:0] n15459;
wire     [31:0] n15460;
wire     [31:0] n15461;
wire     [31:0] n15462;
wire     [31:0] n15463;
wire     [31:0] n15464;
wire     [31:0] n15465;
wire     [31:0] n15466;
wire     [31:0] n15467;
wire     [31:0] n15468;
wire     [31:0] n15469;
wire     [31:0] n15470;
wire     [31:0] n15471;
wire     [31:0] n15472;
wire     [31:0] n15473;
wire     [31:0] n15474;
wire     [31:0] n15475;
wire     [31:0] n15476;
wire     [31:0] n15477;
wire     [31:0] n15478;
wire     [31:0] n15479;
wire     [31:0] n15480;
wire     [31:0] n15481;
wire     [31:0] n15482;
wire     [31:0] n15483;
wire     [31:0] n15484;
wire     [31:0] n15485;
wire     [31:0] n15486;
wire     [31:0] n15487;
wire     [31:0] n15488;
wire     [31:0] n15489;
wire     [31:0] n15490;
wire     [31:0] n15491;
wire     [31:0] n15492;
wire     [31:0] n15493;
wire     [31:0] n15494;
wire     [31:0] n15495;
wire     [31:0] n15496;
wire     [31:0] n15497;
wire     [31:0] n15498;
wire     [31:0] n15499;
wire     [31:0] n15500;
wire     [31:0] n15501;
wire     [31:0] n15502;
wire     [31:0] n15503;
wire     [31:0] n15504;
wire     [31:0] n15505;
wire     [31:0] n15506;
wire     [31:0] n15507;
wire     [31:0] n15508;
wire     [31:0] n15509;
wire     [31:0] n15510;
wire     [31:0] n15511;
wire     [31:0] n15512;
wire     [31:0] n15513;
wire     [31:0] n15514;
wire     [31:0] n15515;
wire     [31:0] n15516;
wire     [31:0] n15517;
wire     [31:0] n15518;
wire     [31:0] n15519;
wire     [31:0] n15520;
wire     [31:0] n15521;
wire     [31:0] n15522;
wire     [31:0] n15523;
wire     [31:0] n15524;
wire     [31:0] n15525;
wire     [31:0] n15526;
wire     [31:0] n15527;
wire     [31:0] n15528;
wire     [31:0] n15529;
wire     [31:0] n15530;
wire     [31:0] n15531;
wire     [31:0] n15532;
wire     [31:0] n15533;
wire     [31:0] n15534;
wire     [31:0] n15535;
wire     [31:0] n15536;
wire     [31:0] n15537;
wire     [31:0] n15538;
wire     [31:0] n15539;
wire     [31:0] n15540;
wire     [31:0] n15541;
wire     [31:0] n15542;
wire     [31:0] n15543;
wire     [31:0] n15544;
wire     [31:0] n15545;
wire     [31:0] n15546;
wire     [31:0] n15547;
wire     [31:0] n15548;
wire     [31:0] n15549;
wire     [31:0] n15550;
wire     [31:0] n15551;
wire     [31:0] n15552;
wire     [31:0] n15553;
wire     [31:0] n15554;
wire     [31:0] n15555;
wire     [31:0] n15556;
wire     [31:0] n15557;
wire     [31:0] n15558;
wire     [31:0] n15559;
wire     [31:0] n15560;
wire     [31:0] n15561;
wire     [31:0] n15562;
wire     [31:0] n15563;
wire     [31:0] n15564;
wire     [31:0] n15565;
wire     [31:0] n15566;
wire     [31:0] n15567;
wire     [31:0] n15568;
wire     [31:0] n15569;
wire     [31:0] n15570;
wire     [31:0] n15571;
wire     [31:0] n15572;
wire     [31:0] n15573;
wire     [31:0] n15574;
wire     [31:0] n15575;
wire     [31:0] n15576;
wire     [31:0] n15577;
wire     [31:0] n15578;
wire     [31:0] n15579;
wire     [31:0] n15580;
wire     [31:0] n15581;
wire     [31:0] n15582;
wire     [31:0] n15583;
wire     [31:0] n15584;
wire     [31:0] n15585;
wire     [31:0] n15586;
wire     [31:0] n15587;
wire     [31:0] n15588;
wire     [31:0] n15589;
wire     [31:0] n15590;
wire     [31:0] n15591;
wire     [31:0] n15592;
wire     [31:0] n15593;
wire     [31:0] n15594;
wire     [31:0] n15595;
wire     [31:0] n15596;
wire     [31:0] n15597;
wire     [31:0] n15598;
wire     [31:0] n15599;
wire     [31:0] n15600;
wire     [31:0] n15601;
wire     [31:0] n15602;
wire     [31:0] n15603;
wire     [31:0] n15604;
wire     [31:0] n15605;
wire     [31:0] n15606;
wire     [31:0] n15607;
wire     [31:0] n15608;
wire     [31:0] n15609;
wire     [31:0] n15610;
wire     [31:0] n15611;
wire     [31:0] n15612;
wire     [31:0] n15613;
wire     [31:0] n15614;
wire     [31:0] n15615;
wire     [31:0] n15616;
wire     [31:0] n15617;
wire     [31:0] n15618;
wire     [31:0] n15619;
wire     [31:0] n15620;
wire     [31:0] n15621;
wire     [31:0] n15622;
wire     [31:0] n15623;
wire     [31:0] n15624;
wire     [31:0] n15625;
wire     [31:0] n15626;
wire     [31:0] n15627;
wire     [31:0] n15628;
wire     [31:0] n15629;
wire     [31:0] n15630;
wire     [31:0] n15631;
wire     [31:0] n15632;
wire     [31:0] n15633;
wire     [31:0] n15634;
wire     [31:0] n15635;
wire     [31:0] n15636;
wire     [31:0] n15637;
wire     [31:0] n15638;
wire     [31:0] n15639;
wire     [31:0] n15640;
wire     [31:0] n15641;
wire     [31:0] n15642;
wire     [31:0] n15643;
wire     [31:0] n15644;
wire     [31:0] n15645;
wire     [31:0] n15646;
wire     [31:0] n15647;
wire     [31:0] n15648;
wire     [31:0] n15649;
wire     [31:0] n15650;
wire     [31:0] n15651;
wire     [31:0] n15652;
wire     [31:0] n15653;
wire     [31:0] n15654;
wire     [31:0] n15655;
wire     [31:0] n15656;
wire     [31:0] n15657;
wire     [31:0] n15658;
wire     [31:0] n15659;
wire     [31:0] n15660;
wire     [31:0] n15661;
wire     [31:0] n15662;
wire     [31:0] n15663;
wire     [31:0] n15664;
wire     [31:0] n15665;
wire     [31:0] n15666;
wire     [31:0] n15667;
wire     [31:0] n15668;
wire     [31:0] n15669;
wire     [31:0] n15670;
wire     [31:0] n15671;
wire     [31:0] n15672;
wire     [31:0] n15673;
wire     [31:0] n15674;
wire     [31:0] n15675;
wire     [31:0] n15676;
wire     [31:0] n15677;
wire     [31:0] n15678;
wire     [31:0] n15679;
wire     [31:0] n15680;
wire     [31:0] n15681;
wire     [31:0] n15682;
wire     [31:0] n15683;
wire     [31:0] n15684;
wire     [31:0] n15685;
wire     [31:0] n15686;
wire     [31:0] n15687;
wire     [31:0] n15688;
wire     [31:0] n15689;
wire     [31:0] n15690;
wire     [31:0] n15691;
wire     [31:0] n15692;
wire     [31:0] n15693;
wire     [31:0] n15694;
wire     [31:0] n15695;
wire     [31:0] n15696;
wire     [31:0] n15697;
wire     [31:0] n15698;
wire     [31:0] n15699;
wire     [31:0] n15700;
wire     [31:0] n15701;
wire     [31:0] n15702;
wire     [31:0] n15703;
wire     [31:0] n15704;
wire     [31:0] n15705;
wire     [31:0] n15706;
wire     [31:0] n15707;
wire     [31:0] n15708;
wire     [31:0] n15709;
wire     [31:0] n15710;
wire     [31:0] n15711;
wire     [31:0] n15712;
wire     [31:0] n15713;
wire     [31:0] n15714;
wire     [31:0] n15715;
wire     [31:0] n15716;
wire     [31:0] n15717;
wire     [31:0] n15718;
wire     [31:0] n15719;
wire     [31:0] n15720;
wire     [31:0] n15721;
wire     [31:0] n15722;
wire     [31:0] n15723;
wire     [31:0] n15724;
wire     [31:0] n15725;
wire     [31:0] n15726;
wire     [31:0] n15727;
wire     [31:0] n15728;
wire     [31:0] n15729;
wire     [31:0] n15730;
wire     [31:0] n15731;
wire     [31:0] n15732;
wire     [31:0] n15733;
wire     [31:0] n15734;
wire     [31:0] n15735;
wire     [31:0] n15736;
wire     [31:0] n15737;
wire     [31:0] n15738;
wire     [31:0] n15739;
wire     [31:0] n15740;
wire     [31:0] n15741;
wire     [31:0] n15742;
wire     [31:0] n15743;
wire     [31:0] n15744;
wire     [31:0] n15745;
wire     [31:0] n15746;
wire     [31:0] n15747;
wire            n15748;
wire            n15749;
wire     [31:0] n15750;
wire     [31:0] n15751;
wire     [31:0] n15752;
wire     [31:0] n15753;
wire     [31:0] n15754;
wire     [31:0] n15755;
wire     [31:0] n15756;
wire     [31:0] n15757;
wire     [31:0] n15758;
wire     [31:0] n15759;
wire     [31:0] n15760;
wire     [31:0] n15761;
wire     [31:0] n15762;
wire     [31:0] n15763;
wire     [31:0] n15764;
wire     [31:0] n15765;
wire     [31:0] n15766;
wire     [31:0] n15767;
wire     [31:0] n15768;
wire     [31:0] n15769;
wire     [31:0] n15770;
wire     [31:0] n15771;
wire     [31:0] n15772;
wire     [31:0] n15773;
wire     [31:0] n15774;
wire     [31:0] n15775;
wire     [31:0] n15776;
wire     [31:0] n15777;
wire     [31:0] n15778;
wire     [31:0] n15779;
wire     [31:0] n15780;
wire     [31:0] n15781;
wire     [31:0] n15782;
wire            n15783;
wire            n15784;
wire            n15785;
wire            n15786;
wire            n15787;
wire            n15788;
wire            n15789;
wire            n15790;
wire            n15791;
wire            n15792;
wire            n15793;
wire            n15794;
wire            n15795;
wire            n15796;
wire            n15797;
wire            n15798;
wire            n15799;
wire            n15800;
wire            n15801;
wire            n15802;
wire            n15803;
wire            n15804;
wire            n15805;
wire            n15806;
wire            n15807;
wire            n15808;
wire            n15809;
wire            n15810;
wire            n15811;
wire            n15812;
wire            n15813;
wire            n15814;
wire            n15815;
wire            n15816;
wire            n15817;
wire            n15818;
wire            n15819;
wire            n15820;
wire            n15821;
wire            n15822;
wire            n15823;
wire            n15824;
wire            n15825;
wire            n15826;
wire            n15827;
wire            n15828;
wire            n15829;
wire            n15830;
wire            n15831;
wire            n15832;
wire            n15833;
wire            n15834;
wire            n15835;
wire            n15836;
wire            n15837;
wire            n15838;
wire            n15839;
wire            n15840;
wire            n15841;
wire            n15842;
wire            n15843;
wire            n15844;
wire            n15845;
wire            n15846;
wire            n15847;
wire            n15848;
wire            n15849;
wire            n15850;
wire            n15851;
wire            n15852;
wire            n15853;
wire            n15854;
wire            n15855;
wire            n15856;
wire            n15857;
wire            n15858;
wire            n15859;
wire            n15860;
wire            n15861;
wire            n15862;
wire            n15863;
wire            n15864;
wire            n15865;
wire            n15866;
wire            n15867;
wire            n15868;
wire            n15869;
wire            n15870;
wire            n15871;
wire            n15872;
wire            n15873;
wire            n15874;
wire            n15875;
wire            n15876;
wire            n15877;
wire            n15878;
wire            n15879;
wire            n15880;
wire            n15881;
wire            n15882;
wire            n15883;
wire            n15884;
wire            n15885;
wire            n15886;
wire            n15887;
wire            n15888;
wire            n15889;
wire            n15890;
wire            n15891;
wire            n15892;
wire            n15893;
wire            n15894;
wire            n15895;
wire            n15896;
wire            n15897;
wire            n15898;
wire            n15899;
wire            n15900;
wire            n15901;
wire            n15902;
wire            n15903;
wire            n15904;
wire            n15905;
wire            n15906;
wire            n15907;
wire            n15908;
wire            n15909;
wire            n15910;
wire            n15911;
wire            n15912;
wire            n15913;
wire            n15914;
wire            n15915;
wire            n15916;
wire            n15917;
wire            n15918;
wire            n15919;
wire            n15920;
wire            n15921;
wire            n15922;
wire            n15923;
wire            n15924;
wire            n15925;
wire            n15926;
wire            n15927;
wire            n15928;
wire            n15929;
wire            n15930;
wire            n15931;
wire            n15932;
wire            n15933;
wire            n15934;
wire            n15935;
wire            n15936;
wire            n15937;
wire            n15938;
wire            n15939;
wire            n15940;
wire            n15941;
wire            n15942;
wire            n15943;
wire            n15944;
wire            n15945;
wire            n15946;
wire            n15947;
wire            n15948;
wire            n15949;
wire            n15950;
wire            n15951;
wire            n15952;
wire            n15953;
wire            n15954;
wire            n15955;
wire            n15956;
wire            n15957;
wire            n15958;
wire            n15959;
wire            n15960;
wire            n15961;
wire            n15962;
wire            n15963;
wire            n15964;
wire            n15965;
wire            n15966;
wire            n15967;
wire            n15968;
wire            n15969;
wire            n15970;
wire            n15971;
wire            n15972;
wire            n15973;
wire            n15974;
wire            n15975;
wire            n15976;
wire            n15977;
wire            n15978;
wire            n15979;
wire            n15980;
wire            n15981;
wire            n15982;
wire            n15983;
wire            n15984;
wire            n15985;
wire            n15986;
wire            n15987;
wire            n15988;
wire            n15989;
wire            n15990;
wire            n15991;
wire            n15992;
wire            n15993;
wire            n15994;
wire            n15995;
wire            n15996;
wire            n15997;
wire            n15998;
wire            n15999;
wire            n16000;
wire            n16001;
wire            n16002;
wire            n16003;
wire            n16004;
wire            n16005;
wire            n16006;
wire            n16007;
wire            n16008;
wire            n16009;
wire            n16010;
wire            n16011;
wire            n16012;
wire            n16013;
wire            n16014;
wire            n16015;
wire            n16016;
wire            n16017;
wire            n16018;
wire            n16019;
wire            n16020;
wire            n16021;
wire            n16022;
wire            n16023;
wire            n16024;
wire            n16025;
wire            n16026;
wire            n16027;
wire            n16028;
wire            n16029;
wire            n16030;
wire            n16031;
wire            n16032;
wire            n16033;
wire            n16034;
wire            n16035;
wire            n16036;
wire            n16037;
wire            n16038;
wire            n16039;
wire            n16040;
wire            n16041;
wire            n16042;
wire            n16043;
wire            n16044;
wire            n16045;
wire            n16046;
wire            n16047;
wire            n16048;
wire            n16049;
wire            n16050;
wire            n16051;
wire            n16052;
wire            n16053;
wire            n16054;
wire            n16055;
wire            n16056;
wire            n16057;
wire            n16058;
wire            n16059;
wire            n16060;
wire            n16061;
wire            n16062;
wire            n16063;
wire            n16064;
wire            n16065;
wire            n16066;
wire            n16067;
wire            n16068;
wire            n16069;
wire            n16070;
wire            n16071;
wire            n16072;
wire            n16073;
wire            n16074;
wire            n16075;
wire            n16076;
wire            n16077;
wire            n16078;
wire            n16079;
wire            n16080;
wire            n16081;
wire            n16082;
wire            n16083;
wire            n16084;
wire            n16085;
wire            n16086;
wire            n16087;
wire            n16088;
wire            n16089;
wire            n16090;
wire            n16091;
wire            n16092;
wire            n16093;
wire            n16094;
wire            n16095;
wire            n16096;
wire            n16097;
wire            n16098;
wire            n16099;
wire            n16100;
wire            n16101;
wire            n16102;
wire            n16103;
wire            n16104;
wire            n16105;
wire            n16106;
wire            n16107;
wire            n16108;
wire            n16109;
wire            n16110;
wire            n16111;
wire            n16112;
wire            n16113;
wire            n16114;
wire            n16115;
wire            n16116;
wire            n16117;
wire            n16118;
wire            n16119;
wire            n16120;
wire            n16121;
wire            n16122;
wire            n16123;
wire            n16124;
wire            n16125;
wire            n16126;
wire            n16127;
wire            n16128;
wire            n16129;
wire            n16130;
wire            n16131;
wire            n16132;
wire            n16133;
wire            n16134;
wire            n16135;
wire            n16136;
wire            n16137;
wire            n16138;
wire            n16139;
wire            n16140;
wire            n16141;
wire            n16142;
wire            n16143;
wire            n16144;
wire            n16145;
wire            n16146;
wire            n16147;
wire            n16148;
wire            n16149;
wire            n16150;
wire            n16151;
wire            n16152;
wire            n16153;
wire            n16154;
wire            n16155;
wire            n16156;
wire            n16157;
wire            n16158;
wire            n16159;
wire            n16160;
wire            n16161;
wire            n16162;
wire            n16163;
wire            n16164;
wire            n16165;
wire            n16166;
wire            n16167;
wire            n16168;
wire            n16169;
wire            n16170;
wire            n16171;
wire            n16172;
wire            n16173;
wire            n16174;
wire            n16175;
wire            n16176;
wire            n16177;
wire            n16178;
wire            n16179;
wire            n16180;
wire            n16181;
wire            n16182;
wire            n16183;
wire            n16184;
wire            n16185;
wire            n16186;
wire            n16187;
wire            n16188;
wire            n16189;
wire            n16190;
wire            n16191;
wire            n16192;
wire            n16193;
wire            n16194;
wire            n16195;
wire            n16196;
wire            n16197;
wire            n16198;
wire            n16199;
wire            n16200;
wire            n16201;
wire            n16202;
wire            n16203;
wire            n16204;
wire            n16205;
wire            n16206;
wire            n16207;
wire            n16208;
wire            n16209;
wire            n16210;
wire            n16211;
wire            n16212;
wire            n16213;
wire            n16214;
wire            n16215;
wire            n16216;
wire            n16217;
wire            n16218;
wire            n16219;
wire            n16220;
wire            n16221;
wire            n16222;
wire            n16223;
wire            n16224;
wire            n16225;
wire            n16226;
wire            n16227;
wire            n16228;
wire            n16229;
wire            n16230;
wire            n16231;
wire            n16232;
wire            n16233;
wire            n16234;
wire            n16235;
wire            n16236;
wire            n16237;
wire            n16238;
wire            n16239;
wire            n16240;
wire            n16241;
wire            n16242;
wire            n16243;
wire            n16244;
wire            n16245;
wire            n16246;
wire            n16247;
wire            n16248;
wire            n16249;
wire            n16250;
wire            n16251;
wire            n16252;
wire            n16253;
wire            n16254;
wire            n16255;
wire            n16256;
wire            n16257;
wire            n16258;
wire            n16259;
wire            n16260;
wire            n16261;
wire            n16262;
wire            n16263;
wire            n16264;
wire            n16265;
wire            n16266;
wire            n16267;
wire            n16268;
wire            n16269;
wire            n16270;
wire            n16271;
wire            n16272;
wire            n16273;
wire            n16274;
wire            n16275;
wire            n16276;
wire            n16277;
wire            n16278;
wire            n16279;
wire            n16280;
wire            n16281;
wire            n16282;
wire            n16283;
wire            n16284;
wire            n16285;
wire            n16286;
wire            n16287;
wire            n16288;
wire            n16289;
wire            n16290;
wire            n16291;
wire            n16292;
wire            n16293;
wire            n16294;
wire            n16295;
wire            n16296;
wire            n16297;
wire            n16298;
wire            n16299;
wire            n16300;
wire            n16301;
wire            n16302;
wire            n16303;
wire            n16304;
wire            n16305;
wire            n16306;
wire            n16307;
wire            n16308;
wire            n16309;
wire            n16310;
wire     [31:0] n16311;
wire     [31:0] n16312;
wire     [31:0] n16313;
wire     [31:0] n16314;
wire     [31:0] n16315;
wire     [31:0] n16316;
wire     [31:0] n16317;
wire     [31:0] n16318;
wire     [31:0] n16319;
wire     [31:0] n16320;
wire     [31:0] n16321;
wire     [31:0] n16322;
wire     [31:0] n16323;
wire     [31:0] n16324;
wire     [31:0] n16325;
wire     [31:0] n16326;
wire     [31:0] n16327;
wire     [31:0] n16328;
wire     [31:0] n16329;
wire     [31:0] n16330;
wire     [31:0] n16331;
wire     [31:0] n16332;
wire     [31:0] n16333;
wire     [31:0] n16334;
wire     [31:0] n16335;
wire     [31:0] n16336;
wire     [31:0] n16337;
wire     [31:0] n16338;
wire     [31:0] n16339;
wire     [31:0] n16340;
wire     [31:0] n16341;
wire     [31:0] n16342;
wire     [31:0] n16343;
wire     [31:0] n16344;
wire     [31:0] n16345;
wire     [31:0] n16346;
wire     [31:0] n16347;
wire     [31:0] n16348;
wire     [31:0] n16349;
wire     [31:0] n16350;
wire     [31:0] n16351;
wire     [31:0] n16352;
wire     [31:0] n16353;
wire     [31:0] n16354;
wire     [31:0] n16355;
wire     [31:0] n16356;
wire     [31:0] n16357;
wire     [31:0] n16358;
wire     [31:0] n16359;
wire     [31:0] n16360;
wire     [31:0] n16361;
wire     [31:0] n16362;
wire     [31:0] n16363;
wire     [31:0] n16364;
wire     [31:0] n16365;
wire     [31:0] n16366;
wire     [31:0] n16367;
wire     [31:0] n16368;
wire     [31:0] n16369;
wire     [31:0] n16370;
wire     [31:0] n16371;
wire     [31:0] n16372;
wire     [31:0] n16373;
wire     [31:0] n16374;
wire     [31:0] n16375;
wire     [31:0] n16376;
wire     [31:0] n16377;
wire     [31:0] n16378;
wire     [31:0] n16379;
wire     [31:0] n16380;
wire     [31:0] n16381;
wire     [31:0] n16382;
wire     [31:0] n16383;
wire     [31:0] n16384;
wire     [31:0] n16385;
wire     [31:0] n16386;
wire     [31:0] n16387;
wire     [31:0] n16388;
wire     [31:0] n16389;
wire     [31:0] n16390;
wire     [31:0] n16391;
wire     [31:0] n16392;
wire     [31:0] n16393;
wire     [31:0] n16394;
wire     [31:0] n16395;
wire     [31:0] n16396;
wire     [31:0] n16397;
wire     [31:0] n16398;
wire     [31:0] n16399;
wire     [31:0] n16400;
wire     [31:0] n16401;
wire     [31:0] n16402;
wire     [31:0] n16403;
wire     [31:0] n16404;
wire     [31:0] n16405;
wire     [31:0] n16406;
wire     [31:0] n16407;
wire     [31:0] n16408;
wire     [31:0] n16409;
wire     [31:0] n16410;
wire     [31:0] n16411;
wire     [31:0] n16412;
wire     [31:0] n16413;
wire     [31:0] n16414;
wire     [31:0] n16415;
wire     [31:0] n16416;
wire     [31:0] n16417;
wire     [31:0] n16418;
wire     [31:0] n16419;
wire     [31:0] n16420;
wire     [31:0] n16421;
wire     [31:0] n16422;
wire     [31:0] n16423;
wire     [31:0] n16424;
wire     [31:0] n16425;
wire     [31:0] n16426;
wire     [31:0] n16427;
wire     [31:0] n16428;
wire     [31:0] n16429;
wire     [31:0] n16430;
wire     [31:0] n16431;
wire     [31:0] n16432;
wire     [31:0] n16433;
wire     [31:0] n16434;
wire     [31:0] n16435;
wire     [31:0] n16436;
wire     [31:0] n16437;
wire     [31:0] n16438;
wire     [31:0] n16439;
wire     [31:0] n16440;
wire     [31:0] n16441;
wire     [31:0] n16442;
wire     [31:0] n16443;
wire     [31:0] n16444;
wire     [31:0] n16445;
wire     [31:0] n16446;
wire     [31:0] n16447;
wire     [31:0] n16448;
wire     [31:0] n16449;
wire     [31:0] n16450;
wire     [31:0] n16451;
wire     [31:0] n16452;
wire     [31:0] n16453;
wire     [31:0] n16454;
wire     [31:0] n16455;
wire     [31:0] n16456;
wire     [31:0] n16457;
wire     [31:0] n16458;
wire     [31:0] n16459;
wire     [31:0] n16460;
wire     [31:0] n16461;
wire     [31:0] n16462;
wire     [31:0] n16463;
wire     [31:0] n16464;
wire     [31:0] n16465;
wire     [31:0] n16466;
wire     [31:0] n16467;
wire     [31:0] n16468;
wire     [31:0] n16469;
wire     [31:0] n16470;
wire     [31:0] n16471;
wire     [31:0] n16472;
wire     [31:0] n16473;
wire     [31:0] n16474;
wire     [31:0] n16475;
wire     [31:0] n16476;
wire     [31:0] n16477;
wire     [31:0] n16478;
wire     [31:0] n16479;
wire     [31:0] n16480;
wire     [31:0] n16481;
wire     [31:0] n16482;
wire     [31:0] n16483;
wire     [31:0] n16484;
wire     [31:0] n16485;
wire     [31:0] n16486;
wire     [31:0] n16487;
wire     [31:0] n16488;
wire     [31:0] n16489;
wire     [31:0] n16490;
wire     [31:0] n16491;
wire     [31:0] n16492;
wire     [31:0] n16493;
wire     [31:0] n16494;
wire     [31:0] n16495;
wire     [31:0] n16496;
wire     [31:0] n16497;
wire     [31:0] n16498;
wire     [31:0] n16499;
wire     [31:0] n16500;
wire     [31:0] n16501;
wire     [31:0] n16502;
wire     [31:0] n16503;
wire     [31:0] n16504;
wire     [31:0] n16505;
wire     [31:0] n16506;
wire     [31:0] n16507;
wire     [31:0] n16508;
wire     [31:0] n16509;
wire     [31:0] n16510;
wire     [31:0] n16511;
wire     [31:0] n16512;
wire     [31:0] n16513;
wire     [31:0] n16514;
wire     [31:0] n16515;
wire     [31:0] n16516;
wire     [31:0] n16517;
wire     [31:0] n16518;
wire     [31:0] n16519;
wire     [31:0] n16520;
wire     [31:0] n16521;
wire     [31:0] n16522;
wire     [31:0] n16523;
wire     [31:0] n16524;
wire     [31:0] n16525;
wire     [31:0] n16526;
wire     [31:0] n16527;
wire     [31:0] n16528;
wire     [31:0] n16529;
wire     [31:0] n16530;
wire     [31:0] n16531;
wire     [31:0] n16532;
wire     [31:0] n16533;
wire     [31:0] n16534;
wire     [31:0] n16535;
wire     [31:0] n16536;
wire     [31:0] n16537;
wire     [31:0] n16538;
wire     [31:0] n16539;
wire     [31:0] n16540;
wire     [31:0] n16541;
wire     [31:0] n16542;
wire     [31:0] n16543;
wire     [31:0] n16544;
wire     [31:0] n16545;
wire     [31:0] n16546;
wire     [31:0] n16547;
wire     [31:0] n16548;
wire     [31:0] n16549;
wire     [31:0] n16550;
wire     [31:0] n16551;
wire     [31:0] n16552;
wire     [31:0] n16553;
wire     [31:0] n16554;
wire     [31:0] n16555;
wire     [31:0] n16556;
wire     [31:0] n16557;
wire     [31:0] n16558;
wire     [31:0] n16559;
wire     [31:0] n16560;
wire     [31:0] n16561;
wire     [31:0] n16562;
wire     [31:0] n16563;
wire     [31:0] n16564;
wire     [31:0] n16565;
wire     [31:0] n16566;
wire     [31:0] n16567;
wire     [31:0] n16568;
wire     [31:0] n16569;
wire     [31:0] n16570;
wire     [31:0] n16571;
wire     [31:0] n16572;
wire     [31:0] n16573;
wire     [31:0] n16574;
wire     [31:0] n16575;
wire     [31:0] n16576;
wire     [31:0] n16577;
wire     [31:0] n16578;
wire     [31:0] n16579;
wire     [31:0] n16580;
wire     [31:0] n16581;
wire     [31:0] n16582;
wire     [31:0] n16583;
wire     [31:0] n16584;
wire     [31:0] n16585;
wire     [31:0] n16586;
wire     [31:0] n16587;
wire     [31:0] n16588;
wire     [31:0] n16589;
wire     [31:0] n16590;
wire     [31:0] n16591;
wire     [31:0] n16592;
wire     [31:0] n16593;
wire     [31:0] n16594;
wire     [31:0] n16595;
wire     [31:0] n16596;
wire     [31:0] n16597;
wire     [31:0] n16598;
wire     [31:0] n16599;
wire     [31:0] n16600;
wire     [31:0] n16601;
wire     [31:0] n16602;
wire     [31:0] n16603;
wire     [31:0] n16604;
wire     [31:0] n16605;
wire     [31:0] n16606;
wire     [31:0] n16607;
wire     [31:0] n16608;
wire     [31:0] n16609;
wire     [31:0] n16610;
wire     [31:0] n16611;
wire     [31:0] n16612;
wire     [31:0] n16613;
wire     [31:0] n16614;
wire     [31:0] n16615;
wire     [31:0] n16616;
wire     [31:0] n16617;
wire     [31:0] n16618;
wire     [31:0] n16619;
wire     [31:0] n16620;
wire     [31:0] n16621;
wire     [31:0] n16622;
wire     [31:0] n16623;
wire     [31:0] n16624;
wire     [31:0] n16625;
wire     [31:0] n16626;
wire     [31:0] n16627;
wire     [31:0] n16628;
wire     [31:0] n16629;
wire     [31:0] n16630;
wire     [31:0] n16631;
wire     [31:0] n16632;
wire     [31:0] n16633;
wire     [31:0] n16634;
wire     [31:0] n16635;
wire     [31:0] n16636;
wire     [31:0] n16637;
wire     [31:0] n16638;
wire     [31:0] n16639;
wire     [31:0] n16640;
wire     [31:0] n16641;
wire     [31:0] n16642;
wire     [31:0] n16643;
wire     [31:0] n16644;
wire     [31:0] n16645;
wire     [31:0] n16646;
wire     [31:0] n16647;
wire     [31:0] n16648;
wire     [31:0] n16649;
wire     [31:0] n16650;
wire     [31:0] n16651;
wire     [31:0] n16652;
wire     [31:0] n16653;
wire     [31:0] n16654;
wire     [31:0] n16655;
wire     [31:0] n16656;
wire     [31:0] n16657;
wire     [31:0] n16658;
wire     [31:0] n16659;
wire     [31:0] n16660;
wire     [31:0] n16661;
wire     [31:0] n16662;
wire     [31:0] n16663;
wire     [31:0] n16664;
wire     [31:0] n16665;
wire     [31:0] n16666;
wire     [31:0] n16667;
wire     [31:0] n16668;
wire     [31:0] n16669;
wire     [31:0] n16670;
wire     [31:0] n16671;
wire     [31:0] n16672;
wire     [31:0] n16673;
wire     [31:0] n16674;
wire     [31:0] n16675;
wire     [31:0] n16676;
wire     [31:0] n16677;
wire     [31:0] n16678;
wire     [31:0] n16679;
wire     [31:0] n16680;
wire     [31:0] n16681;
wire     [31:0] n16682;
wire     [31:0] n16683;
wire     [31:0] n16684;
wire     [31:0] n16685;
wire     [31:0] n16686;
wire     [31:0] n16687;
wire     [31:0] n16688;
wire     [31:0] n16689;
wire     [31:0] n16690;
wire     [31:0] n16691;
wire     [31:0] n16692;
wire     [31:0] n16693;
wire     [31:0] n16694;
wire     [31:0] n16695;
wire     [31:0] n16696;
wire     [31:0] n16697;
wire     [31:0] n16698;
wire     [31:0] n16699;
wire     [31:0] n16700;
wire     [31:0] n16701;
wire     [31:0] n16702;
wire     [31:0] n16703;
wire     [31:0] n16704;
wire     [31:0] n16705;
wire     [31:0] n16706;
wire     [31:0] n16707;
wire     [31:0] n16708;
wire     [31:0] n16709;
wire     [31:0] n16710;
wire     [31:0] n16711;
wire     [31:0] n16712;
wire     [31:0] n16713;
wire     [31:0] n16714;
wire     [31:0] n16715;
wire     [31:0] n16716;
wire     [31:0] n16717;
wire     [31:0] n16718;
wire     [31:0] n16719;
wire     [31:0] n16720;
wire     [31:0] n16721;
wire     [31:0] n16722;
wire     [31:0] n16723;
wire     [31:0] n16724;
wire     [31:0] n16725;
wire     [31:0] n16726;
wire     [31:0] n16727;
wire     [31:0] n16728;
wire     [31:0] n16729;
wire     [31:0] n16730;
wire     [31:0] n16731;
wire     [31:0] n16732;
wire     [31:0] n16733;
wire     [31:0] n16734;
wire     [31:0] n16735;
wire     [31:0] n16736;
wire     [31:0] n16737;
wire     [31:0] n16738;
wire     [31:0] n16739;
wire     [31:0] n16740;
wire     [31:0] n16741;
wire     [31:0] n16742;
wire     [31:0] n16743;
wire     [31:0] n16744;
wire     [31:0] n16745;
wire     [31:0] n16746;
wire     [31:0] n16747;
wire     [31:0] n16748;
wire     [31:0] n16749;
wire     [31:0] n16750;
wire     [31:0] n16751;
wire     [31:0] n16752;
wire     [31:0] n16753;
wire     [31:0] n16754;
wire     [31:0] n16755;
wire     [31:0] n16756;
wire     [31:0] n16757;
wire     [31:0] n16758;
wire     [31:0] n16759;
wire     [31:0] n16760;
wire     [31:0] n16761;
wire     [31:0] n16762;
wire     [31:0] n16763;
wire     [31:0] n16764;
wire     [31:0] n16765;
wire     [31:0] n16766;
wire     [31:0] n16767;
wire     [31:0] n16768;
wire     [31:0] n16769;
wire     [31:0] n16770;
wire     [31:0] n16771;
wire     [31:0] n16772;
wire     [31:0] n16773;
wire     [31:0] n16774;
wire     [31:0] n16775;
wire     [31:0] n16776;
wire     [31:0] n16777;
wire     [31:0] n16778;
wire     [31:0] n16779;
wire     [31:0] n16780;
wire     [31:0] n16781;
wire     [31:0] n16782;
wire     [31:0] n16783;
wire     [31:0] n16784;
wire     [31:0] n16785;
wire     [31:0] n16786;
wire     [31:0] n16787;
wire     [31:0] n16788;
wire     [31:0] n16789;
wire     [31:0] n16790;
wire     [31:0] n16791;
wire     [31:0] n16792;
wire     [31:0] n16793;
wire     [31:0] n16794;
wire     [31:0] n16795;
wire     [31:0] n16796;
wire     [31:0] n16797;
wire     [31:0] n16798;
wire     [31:0] n16799;
wire     [31:0] n16800;
wire     [31:0] n16801;
wire     [31:0] n16802;
wire     [31:0] n16803;
wire     [31:0] n16804;
wire     [31:0] n16805;
wire     [31:0] n16806;
wire     [31:0] n16807;
wire     [31:0] n16808;
wire     [31:0] n16809;
wire     [31:0] n16810;
wire     [31:0] n16811;
wire     [31:0] n16812;
wire     [31:0] n16813;
wire     [31:0] n16814;
wire     [31:0] n16815;
wire     [31:0] n16816;
wire     [31:0] n16817;
wire     [31:0] n16818;
wire     [31:0] n16819;
wire     [31:0] n16820;
wire     [31:0] n16821;
wire     [31:0] n16822;
wire     [31:0] n16823;
wire     [31:0] n16824;
wire     [31:0] n16825;
wire     [31:0] n16826;
wire     [31:0] n16827;
wire     [31:0] n16828;
wire     [31:0] n16829;
wire     [31:0] n16830;
wire     [31:0] n16831;
wire     [31:0] n16832;
wire            n16833;
wire            n16834;
wire            n16835;
wire            n16836;
wire            n16837;
wire            n16838;
wire            n16839;
wire            n16840;
wire            n16841;
wire            n16842;
wire            n16843;
wire            n16844;
wire            n16845;
wire            n16846;
wire            n16847;
wire            n16848;
wire            n16849;
wire            n16850;
wire            n16851;
wire            n16852;
wire            n16853;
wire            n16854;
wire            n16855;
wire            n16856;
wire            n16857;
wire            n16858;
wire            n16859;
wire            n16860;
wire            n16861;
wire            n16862;
wire            n16863;
wire            n16864;
wire            n16865;
wire            n16866;
wire            n16867;
wire            n16868;
wire            n16869;
wire            n16870;
wire            n16871;
wire            n16872;
wire            n16873;
wire            n16874;
wire            n16875;
wire            n16876;
wire            n16877;
wire            n16878;
wire            n16879;
wire            n16880;
wire            n16881;
wire            n16882;
wire            n16883;
wire            n16884;
wire            n16885;
wire            n16886;
wire            n16887;
wire            n16888;
wire            n16889;
wire            n16890;
wire            n16891;
wire            n16892;
wire            n16893;
wire            n16894;
wire            n16895;
wire            n16896;
wire            n16897;
wire            n16898;
wire            n16899;
wire            n16900;
wire            n16901;
wire            n16902;
wire            n16903;
wire            n16904;
wire            n16905;
wire            n16906;
wire            n16907;
wire            n16908;
wire            n16909;
wire            n16910;
wire            n16911;
wire            n16912;
wire            n16913;
wire            n16914;
wire            n16915;
wire            n16916;
wire            n16917;
wire            n16918;
wire            n16919;
wire            n16920;
wire            n16921;
wire            n16922;
wire            n16923;
wire            n16924;
wire            n16925;
wire            n16926;
wire            n16927;
wire            n16928;
wire            n16929;
wire            n16930;
wire            n16931;
wire            n16932;
wire            n16933;
wire            n16934;
wire            n16935;
wire            n16936;
wire            n16937;
wire            n16938;
wire            n16939;
wire            n16940;
wire            n16941;
wire            n16942;
wire            n16943;
wire            n16944;
wire            n16945;
wire            n16946;
wire            n16947;
wire            n16948;
wire            n16949;
wire            n16950;
wire            n16951;
wire            n16952;
wire            n16953;
wire            n16954;
wire            n16955;
wire            n16956;
wire            n16957;
wire            n16958;
wire            n16959;
wire            n16960;
wire            n16961;
wire            n16962;
wire            n16963;
wire            n16964;
wire            n16965;
wire            n16966;
wire            n16967;
wire            n16968;
wire            n16969;
wire            n16970;
wire            n16971;
wire            n16972;
wire            n16973;
wire            n16974;
wire            n16975;
wire            n16976;
wire            n16977;
wire            n16978;
wire            n16979;
wire            n16980;
wire            n16981;
wire            n16982;
wire            n16983;
wire            n16984;
wire            n16985;
wire            n16986;
wire            n16987;
wire            n16988;
wire            n16989;
wire            n16990;
wire            n16991;
wire            n16992;
wire            n16993;
wire            n16994;
wire            n16995;
wire            n16996;
wire            n16997;
wire            n16998;
wire            n16999;
wire            n17000;
wire            n17001;
wire            n17002;
wire            n17003;
wire            n17004;
wire            n17005;
wire            n17006;
wire            n17007;
wire            n17008;
wire            n17009;
wire            n17010;
wire            n17011;
wire            n17012;
wire            n17013;
wire            n17014;
wire            n17015;
wire            n17016;
wire            n17017;
wire            n17018;
wire            n17019;
wire            n17020;
wire            n17021;
wire            n17022;
wire            n17023;
wire            n17024;
wire            n17025;
wire            n17026;
wire            n17027;
wire            n17028;
wire            n17029;
wire            n17030;
wire            n17031;
wire            n17032;
wire            n17033;
wire            n17034;
wire            n17035;
wire            n17036;
wire            n17037;
wire            n17038;
wire            n17039;
wire            n17040;
wire            n17041;
wire            n17042;
wire            n17043;
wire            n17044;
wire            n17045;
wire            n17046;
wire            n17047;
wire            n17048;
wire            n17049;
wire            n17050;
wire            n17051;
wire            n17052;
wire            n17053;
wire            n17054;
wire            n17055;
wire            n17056;
wire            n17057;
wire            n17058;
wire            n17059;
wire            n17060;
wire            n17061;
wire            n17062;
wire            n17063;
wire            n17064;
wire            n17065;
wire            n17066;
wire            n17067;
wire            n17068;
wire            n17069;
wire            n17070;
wire            n17071;
wire            n17072;
wire            n17073;
wire            n17074;
wire            n17075;
wire            n17076;
wire            n17077;
wire            n17078;
wire            n17079;
wire            n17080;
wire            n17081;
wire            n17082;
wire            n17083;
wire            n17084;
wire            n17085;
wire            n17086;
wire            n17087;
wire            n17088;
wire            n17089;
wire            n17090;
wire            n17091;
wire            n17092;
wire            n17093;
wire            n17094;
wire            n17095;
wire            n17096;
wire            n17097;
wire            n17098;
wire            n17099;
wire            n17100;
wire            n17101;
wire            n17102;
wire            n17103;
wire            n17104;
wire            n17105;
wire            n17106;
wire            n17107;
wire            n17108;
wire            n17109;
wire            n17110;
wire            n17111;
wire            n17112;
wire            n17113;
wire            n17114;
wire            n17115;
wire            n17116;
wire            n17117;
wire            n17118;
wire            n17119;
wire            n17120;
wire            n17121;
wire            n17122;
wire            n17123;
wire            n17124;
wire            n17125;
wire            n17126;
wire            n17127;
wire            n17128;
wire            n17129;
wire            n17130;
wire            n17131;
wire            n17132;
wire            n17133;
wire            n17134;
wire            n17135;
wire            n17136;
wire            n17137;
wire            n17138;
wire            n17139;
wire            n17140;
wire            n17141;
wire            n17142;
wire            n17143;
wire            n17144;
wire            n17145;
wire            n17146;
wire            n17147;
wire            n17148;
wire            n17149;
wire            n17150;
wire            n17151;
wire            n17152;
wire            n17153;
wire            n17154;
wire            n17155;
wire            n17156;
wire            n17157;
wire            n17158;
wire            n17159;
wire            n17160;
wire            n17161;
wire            n17162;
wire            n17163;
wire            n17164;
wire            n17165;
wire            n17166;
wire            n17167;
wire            n17168;
wire            n17169;
wire            n17170;
wire            n17171;
wire            n17172;
wire            n17173;
wire            n17174;
wire            n17175;
wire            n17176;
wire            n17177;
wire            n17178;
wire            n17179;
wire            n17180;
wire            n17181;
wire            n17182;
wire            n17183;
wire            n17184;
wire            n17185;
wire            n17186;
wire            n17187;
wire            n17188;
wire            n17189;
wire            n17190;
wire            n17191;
wire            n17192;
wire            n17193;
wire            n17194;
wire            n17195;
wire            n17196;
wire            n17197;
wire            n17198;
wire            n17199;
wire            n17200;
wire            n17201;
wire            n17202;
wire            n17203;
wire            n17204;
wire            n17205;
wire            n17206;
wire            n17207;
wire            n17208;
wire            n17209;
wire            n17210;
wire            n17211;
wire            n17212;
wire            n17213;
wire            n17214;
wire            n17215;
wire            n17216;
wire            n17217;
wire            n17218;
wire            n17219;
wire            n17220;
wire            n17221;
wire            n17222;
wire            n17223;
wire            n17224;
wire            n17225;
wire            n17226;
wire            n17227;
wire            n17228;
wire            n17229;
wire            n17230;
wire            n17231;
wire            n17232;
wire            n17233;
wire            n17234;
wire            n17235;
wire            n17236;
wire            n17237;
wire            n17238;
wire            n17239;
wire            n17240;
wire            n17241;
wire            n17242;
wire            n17243;
wire            n17244;
wire            n17245;
wire            n17246;
wire            n17247;
wire            n17248;
wire            n17249;
wire            n17250;
wire            n17251;
wire            n17252;
wire            n17253;
wire            n17254;
wire            n17255;
wire            n17256;
wire            n17257;
wire            n17258;
wire            n17259;
wire            n17260;
wire            n17261;
wire            n17262;
wire            n17263;
wire            n17264;
wire            n17265;
wire            n17266;
wire            n17267;
wire            n17268;
wire            n17269;
wire            n17270;
wire            n17271;
wire            n17272;
wire            n17273;
wire            n17274;
wire            n17275;
wire            n17276;
wire            n17277;
wire            n17278;
wire            n17279;
wire            n17280;
wire            n17281;
wire            n17282;
wire            n17283;
wire            n17284;
wire            n17285;
wire            n17286;
wire            n17287;
wire            n17288;
wire            n17289;
wire            n17290;
wire            n17291;
wire            n17292;
wire            n17293;
wire            n17294;
wire            n17295;
wire            n17296;
wire            n17297;
wire            n17298;
wire            n17299;
wire            n17300;
wire            n17301;
wire            n17302;
wire            n17303;
wire            n17304;
wire            n17305;
wire            n17306;
wire            n17307;
wire            n17308;
wire            n17309;
wire            n17310;
wire            n17311;
wire            n17312;
wire            n17313;
wire            n17314;
wire            n17315;
wire            n17316;
wire            n17317;
wire            n17318;
wire            n17319;
wire            n17320;
wire            n17321;
wire            n17322;
wire            n17323;
wire            n17324;
wire            n17325;
wire            n17326;
wire            n17327;
wire            n17328;
wire            n17329;
wire            n17330;
wire            n17331;
wire            n17332;
wire            n17333;
wire            n17334;
wire            n17335;
wire            n17336;
wire            n17337;
wire            n17338;
wire            n17339;
wire            n17340;
wire            n17341;
wire            n17342;
wire            n17343;
wire            n17344;
wire     [31:0] n17345;
wire     [31:0] n17346;
wire     [31:0] n17347;
wire     [31:0] n17348;
wire     [31:0] n17349;
wire     [31:0] n17350;
wire     [31:0] n17351;
wire     [31:0] n17352;
wire     [31:0] n17353;
wire     [31:0] n17354;
wire     [31:0] n17355;
wire     [31:0] n17356;
wire     [31:0] n17357;
wire     [31:0] n17358;
wire     [31:0] n17359;
wire     [31:0] n17360;
wire     [31:0] n17361;
wire     [31:0] n17362;
wire     [31:0] n17363;
wire     [31:0] n17364;
wire     [31:0] n17365;
wire     [31:0] n17366;
wire     [31:0] n17367;
wire     [31:0] n17368;
wire     [31:0] n17369;
wire     [31:0] n17370;
wire     [31:0] n17371;
wire     [31:0] n17372;
wire     [31:0] n17373;
wire     [31:0] n17374;
wire     [31:0] n17375;
wire     [31:0] n17376;
wire     [31:0] n17377;
wire     [31:0] n17378;
wire     [31:0] n17379;
wire     [31:0] n17380;
wire     [31:0] n17381;
wire     [31:0] n17382;
wire     [31:0] n17383;
wire     [31:0] n17384;
wire     [31:0] n17385;
wire     [31:0] n17386;
wire     [31:0] n17387;
wire     [31:0] n17388;
wire     [31:0] n17389;
wire     [31:0] n17390;
wire     [31:0] n17391;
wire     [31:0] n17392;
wire     [31:0] n17393;
wire     [31:0] n17394;
wire     [31:0] n17395;
wire     [31:0] n17396;
wire     [31:0] n17397;
wire     [31:0] n17398;
wire     [31:0] n17399;
wire     [31:0] n17400;
wire     [31:0] n17401;
wire     [31:0] n17402;
wire     [31:0] n17403;
wire     [31:0] n17404;
wire     [31:0] n17405;
wire     [31:0] n17406;
wire     [31:0] n17407;
wire     [31:0] n17408;
wire     [31:0] n17409;
wire     [31:0] n17410;
wire     [31:0] n17411;
wire     [31:0] n17412;
wire     [31:0] n17413;
wire     [31:0] n17414;
wire     [31:0] n17415;
wire     [31:0] n17416;
wire     [31:0] n17417;
wire     [31:0] n17418;
wire     [31:0] n17419;
wire     [31:0] n17420;
wire     [31:0] n17421;
wire     [31:0] n17422;
wire     [31:0] n17423;
wire     [31:0] n17424;
wire     [31:0] n17425;
wire     [31:0] n17426;
wire     [31:0] n17427;
wire     [31:0] n17428;
wire     [31:0] n17429;
wire     [31:0] n17430;
wire     [31:0] n17431;
wire     [31:0] n17432;
wire     [31:0] n17433;
wire     [31:0] n17434;
wire     [31:0] n17435;
wire     [31:0] n17436;
wire     [31:0] n17437;
wire     [31:0] n17438;
wire     [31:0] n17439;
wire     [31:0] n17440;
wire     [31:0] n17441;
wire     [31:0] n17442;
wire     [31:0] n17443;
wire     [31:0] n17444;
wire     [31:0] n17445;
wire     [31:0] n17446;
wire     [31:0] n17447;
wire     [31:0] n17448;
wire     [31:0] n17449;
wire     [31:0] n17450;
wire     [31:0] n17451;
wire     [31:0] n17452;
wire     [31:0] n17453;
wire     [31:0] n17454;
wire     [31:0] n17455;
wire     [31:0] n17456;
wire     [31:0] n17457;
wire     [31:0] n17458;
wire     [31:0] n17459;
wire     [31:0] n17460;
wire     [31:0] n17461;
wire     [31:0] n17462;
wire     [31:0] n17463;
wire     [31:0] n17464;
wire     [31:0] n17465;
wire     [31:0] n17466;
wire     [31:0] n17467;
wire     [31:0] n17468;
wire     [31:0] n17469;
wire     [31:0] n17470;
wire     [31:0] n17471;
wire     [31:0] n17472;
wire     [31:0] n17473;
wire     [31:0] n17474;
wire     [31:0] n17475;
wire     [31:0] n17476;
wire     [31:0] n17477;
wire     [31:0] n17478;
wire     [31:0] n17479;
wire     [31:0] n17480;
wire     [31:0] n17481;
wire     [31:0] n17482;
wire     [31:0] n17483;
wire     [31:0] n17484;
wire     [31:0] n17485;
wire     [31:0] n17486;
wire     [31:0] n17487;
wire     [31:0] n17488;
wire     [31:0] n17489;
wire     [31:0] n17490;
wire     [31:0] n17491;
wire     [31:0] n17492;
wire     [31:0] n17493;
wire     [31:0] n17494;
wire     [31:0] n17495;
wire     [31:0] n17496;
wire     [31:0] n17497;
wire     [31:0] n17498;
wire     [31:0] n17499;
wire     [31:0] n17500;
wire     [31:0] n17501;
wire     [31:0] n17502;
wire     [31:0] n17503;
wire     [31:0] n17504;
wire     [31:0] n17505;
wire     [31:0] n17506;
wire     [31:0] n17507;
wire     [31:0] n17508;
wire     [31:0] n17509;
wire     [31:0] n17510;
wire     [31:0] n17511;
wire     [31:0] n17512;
wire     [31:0] n17513;
wire     [31:0] n17514;
wire     [31:0] n17515;
wire     [31:0] n17516;
wire     [31:0] n17517;
wire     [31:0] n17518;
wire     [31:0] n17519;
wire     [31:0] n17520;
wire     [31:0] n17521;
wire     [31:0] n17522;
wire     [31:0] n17523;
wire     [31:0] n17524;
wire     [31:0] n17525;
wire     [31:0] n17526;
wire     [31:0] n17527;
wire     [31:0] n17528;
wire     [31:0] n17529;
wire     [31:0] n17530;
wire     [31:0] n17531;
wire     [31:0] n17532;
wire     [31:0] n17533;
wire     [31:0] n17534;
wire     [31:0] n17535;
wire     [31:0] n17536;
wire     [31:0] n17537;
wire     [31:0] n17538;
wire     [31:0] n17539;
wire     [31:0] n17540;
wire     [31:0] n17541;
wire     [31:0] n17542;
wire     [31:0] n17543;
wire     [31:0] n17544;
wire     [31:0] n17545;
wire     [31:0] n17546;
wire     [31:0] n17547;
wire     [31:0] n17548;
wire     [31:0] n17549;
wire     [31:0] n17550;
wire     [31:0] n17551;
wire     [31:0] n17552;
wire     [31:0] n17553;
wire     [31:0] n17554;
wire     [31:0] n17555;
wire     [31:0] n17556;
wire     [31:0] n17557;
wire     [31:0] n17558;
wire     [31:0] n17559;
wire     [31:0] n17560;
wire     [31:0] n17561;
wire     [31:0] n17562;
wire     [31:0] n17563;
wire     [31:0] n17564;
wire     [31:0] n17565;
wire     [31:0] n17566;
wire     [31:0] n17567;
wire     [31:0] n17568;
wire     [31:0] n17569;
wire     [31:0] n17570;
wire     [31:0] n17571;
wire     [31:0] n17572;
wire     [31:0] n17573;
wire     [31:0] n17574;
wire     [31:0] n17575;
wire     [31:0] n17576;
wire     [31:0] n17577;
wire     [31:0] n17578;
wire     [31:0] n17579;
wire     [31:0] n17580;
wire     [31:0] n17581;
wire     [31:0] n17582;
wire     [31:0] n17583;
wire     [31:0] n17584;
wire     [31:0] n17585;
wire     [31:0] n17586;
wire     [31:0] n17587;
wire     [31:0] n17588;
wire     [31:0] n17589;
wire     [31:0] n17590;
wire     [31:0] n17591;
wire     [31:0] n17592;
wire     [31:0] n17593;
wire     [31:0] n17594;
wire     [31:0] n17595;
wire     [31:0] n17596;
wire     [31:0] n17597;
wire     [31:0] n17598;
wire     [31:0] n17599;
wire     [31:0] n17600;
wire     [31:0] n17601;
wire     [31:0] n17602;
wire     [31:0] n17603;
wire     [31:0] n17604;
wire     [31:0] n17605;
wire     [31:0] n17606;
wire     [31:0] n17607;
wire     [31:0] n17608;
wire     [31:0] n17609;
wire     [31:0] n17610;
wire     [31:0] n17611;
wire     [31:0] n17612;
wire     [31:0] n17613;
wire     [31:0] n17614;
wire     [31:0] n17615;
wire     [31:0] n17616;
wire     [31:0] n17617;
wire     [31:0] n17618;
wire     [31:0] n17619;
wire     [31:0] n17620;
wire     [31:0] n17621;
wire     [31:0] n17622;
wire     [31:0] n17623;
wire     [31:0] n17624;
wire     [31:0] n17625;
wire     [31:0] n17626;
wire     [31:0] n17627;
wire     [31:0] n17628;
wire     [31:0] n17629;
wire     [31:0] n17630;
wire     [31:0] n17631;
wire     [31:0] n17632;
wire     [31:0] n17633;
wire     [31:0] n17634;
wire     [31:0] n17635;
wire     [31:0] n17636;
wire     [31:0] n17637;
wire     [31:0] n17638;
wire     [31:0] n17639;
wire     [31:0] n17640;
wire     [31:0] n17641;
wire     [31:0] n17642;
wire     [31:0] n17643;
wire     [31:0] n17644;
wire     [31:0] n17645;
wire     [31:0] n17646;
wire     [31:0] n17647;
wire     [31:0] n17648;
wire     [31:0] n17649;
wire     [31:0] n17650;
wire     [31:0] n17651;
wire     [31:0] n17652;
wire     [31:0] n17653;
wire     [31:0] n17654;
wire     [31:0] n17655;
wire     [31:0] n17656;
wire     [31:0] n17657;
wire     [31:0] n17658;
wire     [31:0] n17659;
wire     [31:0] n17660;
wire     [31:0] n17661;
wire     [31:0] n17662;
wire     [31:0] n17663;
wire     [31:0] n17664;
wire     [31:0] n17665;
wire     [31:0] n17666;
wire     [31:0] n17667;
wire     [31:0] n17668;
wire     [31:0] n17669;
wire     [31:0] n17670;
wire     [31:0] n17671;
wire     [31:0] n17672;
wire     [31:0] n17673;
wire     [31:0] n17674;
wire     [31:0] n17675;
wire     [31:0] n17676;
wire     [31:0] n17677;
wire     [31:0] n17678;
wire     [31:0] n17679;
wire     [31:0] n17680;
wire     [31:0] n17681;
wire     [31:0] n17682;
wire     [31:0] n17683;
wire     [31:0] n17684;
wire     [31:0] n17685;
wire     [31:0] n17686;
wire     [31:0] n17687;
wire     [31:0] n17688;
wire     [31:0] n17689;
wire     [31:0] n17690;
wire     [31:0] n17691;
wire     [31:0] n17692;
wire     [31:0] n17693;
wire     [31:0] n17694;
wire     [31:0] n17695;
wire     [31:0] n17696;
wire     [31:0] n17697;
wire     [31:0] n17698;
wire     [31:0] n17699;
wire     [31:0] n17700;
wire     [31:0] n17701;
wire     [31:0] n17702;
wire     [31:0] n17703;
wire     [31:0] n17704;
wire     [31:0] n17705;
wire     [31:0] n17706;
wire     [31:0] n17707;
wire     [31:0] n17708;
wire     [31:0] n17709;
wire     [31:0] n17710;
wire     [31:0] n17711;
wire     [31:0] n17712;
wire     [31:0] n17713;
wire     [31:0] n17714;
wire     [31:0] n17715;
wire     [31:0] n17716;
wire     [31:0] n17717;
wire     [31:0] n17718;
wire     [31:0] n17719;
wire     [31:0] n17720;
wire     [31:0] n17721;
wire     [31:0] n17722;
wire     [31:0] n17723;
wire     [31:0] n17724;
wire     [31:0] n17725;
wire     [31:0] n17726;
wire     [31:0] n17727;
wire     [31:0] n17728;
wire     [31:0] n17729;
wire     [31:0] n17730;
wire     [31:0] n17731;
wire     [31:0] n17732;
wire     [31:0] n17733;
wire     [31:0] n17734;
wire     [31:0] n17735;
wire     [31:0] n17736;
wire     [31:0] n17737;
wire     [31:0] n17738;
wire     [31:0] n17739;
wire     [31:0] n17740;
wire     [31:0] n17741;
wire     [31:0] n17742;
wire     [31:0] n17743;
wire     [31:0] n17744;
wire     [31:0] n17745;
wire     [31:0] n17746;
wire     [31:0] n17747;
wire     [31:0] n17748;
wire     [31:0] n17749;
wire     [31:0] n17750;
wire     [31:0] n17751;
wire     [31:0] n17752;
wire     [31:0] n17753;
wire     [31:0] n17754;
wire     [31:0] n17755;
wire     [31:0] n17756;
wire     [31:0] n17757;
wire     [31:0] n17758;
wire     [31:0] n17759;
wire     [31:0] n17760;
wire     [31:0] n17761;
wire     [31:0] n17762;
wire     [31:0] n17763;
wire     [31:0] n17764;
wire     [31:0] n17765;
wire     [31:0] n17766;
wire     [31:0] n17767;
wire     [31:0] n17768;
wire     [31:0] n17769;
wire     [31:0] n17770;
wire     [31:0] n17771;
wire     [31:0] n17772;
wire     [31:0] n17773;
wire     [31:0] n17774;
wire     [31:0] n17775;
wire     [31:0] n17776;
wire     [31:0] n17777;
wire     [31:0] n17778;
wire     [31:0] n17779;
wire     [31:0] n17780;
wire     [31:0] n17781;
wire     [31:0] n17782;
wire     [31:0] n17783;
wire     [31:0] n17784;
wire     [31:0] n17785;
wire     [31:0] n17786;
wire     [31:0] n17787;
wire     [31:0] n17788;
wire     [31:0] n17789;
wire     [31:0] n17790;
wire     [31:0] n17791;
wire     [31:0] n17792;
wire     [31:0] n17793;
wire     [31:0] n17794;
wire     [31:0] n17795;
wire     [31:0] n17796;
wire     [31:0] n17797;
wire     [31:0] n17798;
wire     [31:0] n17799;
wire     [31:0] n17800;
wire     [31:0] n17801;
wire     [31:0] n17802;
wire     [31:0] n17803;
wire     [31:0] n17804;
wire     [31:0] n17805;
wire     [31:0] n17806;
wire     [31:0] n17807;
wire     [31:0] n17808;
wire     [31:0] n17809;
wire     [31:0] n17810;
wire     [31:0] n17811;
wire     [31:0] n17812;
wire     [31:0] n17813;
wire     [31:0] n17814;
wire     [31:0] n17815;
wire     [31:0] n17816;
wire     [31:0] n17817;
wire     [31:0] n17818;
wire     [31:0] n17819;
wire     [31:0] n17820;
wire     [31:0] n17821;
wire     [31:0] n17822;
wire     [31:0] n17823;
wire     [31:0] n17824;
wire     [31:0] n17825;
wire     [31:0] n17826;
wire     [31:0] n17827;
wire     [31:0] n17828;
wire     [31:0] n17829;
wire     [31:0] n17830;
wire     [31:0] n17831;
wire     [31:0] n17832;
wire     [31:0] n17833;
wire     [31:0] n17834;
wire     [31:0] n17835;
wire     [31:0] n17836;
wire     [31:0] n17837;
wire     [31:0] n17838;
wire     [31:0] n17839;
wire     [31:0] n17840;
wire     [31:0] n17841;
wire     [31:0] n17842;
wire     [31:0] n17843;
wire     [31:0] n17844;
wire     [31:0] n17845;
wire     [31:0] n17846;
wire     [31:0] n17847;
wire     [31:0] n17848;
wire     [31:0] n17849;
wire     [31:0] n17850;
wire     [31:0] n17851;
wire     [31:0] n17852;
wire     [31:0] n17853;
wire     [31:0] n17854;
wire     [31:0] n17855;
wire     [31:0] n17856;
wire     [31:0] n17857;
wire     [31:0] n17858;
wire     [31:0] n17859;
wire     [31:0] n17860;
wire     [31:0] n17861;
wire     [31:0] n17862;
wire     [31:0] n17863;
wire     [31:0] n17864;
wire     [31:0] n17865;
wire     [31:0] n17866;
wire            n17867;
wire            n17868;
wire     [31:0] n17869;
wire     [31:0] n17870;
wire     [31:0] n17871;
wire     [31:0] n17872;
wire     [31:0] n17873;
wire     [31:0] n17874;
wire     [31:0] n17875;
wire     [31:0] n17876;
wire     [31:0] n17877;
wire     [31:0] n17878;
wire     [31:0] n17879;
wire     [31:0] n17880;
wire     [31:0] n17881;
wire     [31:0] n17882;
wire     [31:0] n17883;
wire     [31:0] n17884;
wire     [31:0] n17885;
wire     [31:0] n17886;
wire     [31:0] n17887;
wire     [31:0] n17888;
wire     [31:0] n17889;
wire     [31:0] n17890;
wire     [31:0] n17891;
wire     [31:0] n17892;
wire     [31:0] n17893;
wire     [31:0] n17894;
wire     [31:0] n17895;
wire     [31:0] n17896;
wire     [31:0] n17897;
wire     [31:0] n17898;
wire     [31:0] n17899;
wire     [31:0] n17900;
wire     [31:0] n17901;
wire            n17902;
wire            n17903;
wire            n17904;
wire            n17905;
wire            n17906;
wire            n17907;
wire            n17908;
wire            n17909;
wire            n17910;
wire            n17911;
wire            n17912;
wire            n17913;
wire            n17914;
wire            n17915;
wire            n17916;
wire            n17917;
wire            n17918;
wire            n17919;
wire            n17920;
wire            n17921;
wire            n17922;
wire            n17923;
wire            n17924;
wire            n17925;
wire            n17926;
wire            n17927;
wire            n17928;
wire            n17929;
wire            n17930;
wire            n17931;
wire            n17932;
wire            n17933;
wire            n17934;
wire            n17935;
wire            n17936;
wire            n17937;
wire            n17938;
wire            n17939;
wire            n17940;
wire            n17941;
wire            n17942;
wire            n17943;
wire            n17944;
wire            n17945;
wire            n17946;
wire            n17947;
wire            n17948;
wire            n17949;
wire            n17950;
wire            n17951;
wire            n17952;
wire            n17953;
wire            n17954;
wire            n17955;
wire            n17956;
wire            n17957;
wire            n17958;
wire            n17959;
wire            n17960;
wire            n17961;
wire            n17962;
wire            n17963;
wire            n17964;
wire            n17965;
wire            n17966;
wire            n17967;
wire            n17968;
wire            n17969;
wire            n17970;
wire            n17971;
wire            n17972;
wire            n17973;
wire            n17974;
wire            n17975;
wire            n17976;
wire            n17977;
wire            n17978;
wire            n17979;
wire            n17980;
wire            n17981;
wire            n17982;
wire            n17983;
wire            n17984;
wire            n17985;
wire            n17986;
wire            n17987;
wire            n17988;
wire            n17989;
wire            n17990;
wire            n17991;
wire            n17992;
wire            n17993;
wire            n17994;
wire            n17995;
wire            n17996;
wire            n17997;
wire            n17998;
wire            n17999;
wire            n18000;
wire            n18001;
wire            n18002;
wire            n18003;
wire            n18004;
wire            n18005;
wire            n18006;
wire            n18007;
wire            n18008;
wire            n18009;
wire            n18010;
wire            n18011;
wire            n18012;
wire            n18013;
wire            n18014;
wire            n18015;
wire            n18016;
wire            n18017;
wire            n18018;
wire            n18019;
wire            n18020;
wire            n18021;
wire            n18022;
wire            n18023;
wire            n18024;
wire            n18025;
wire            n18026;
wire            n18027;
wire            n18028;
wire            n18029;
wire            n18030;
wire            n18031;
wire            n18032;
wire            n18033;
wire            n18034;
wire            n18035;
wire            n18036;
wire            n18037;
wire            n18038;
wire            n18039;
wire            n18040;
wire            n18041;
wire            n18042;
wire            n18043;
wire            n18044;
wire            n18045;
wire            n18046;
wire            n18047;
wire            n18048;
wire            n18049;
wire            n18050;
wire            n18051;
wire            n18052;
wire            n18053;
wire            n18054;
wire            n18055;
wire            n18056;
wire            n18057;
wire            n18058;
wire            n18059;
wire            n18060;
wire            n18061;
wire            n18062;
wire            n18063;
wire            n18064;
wire            n18065;
wire            n18066;
wire            n18067;
wire            n18068;
wire            n18069;
wire            n18070;
wire            n18071;
wire            n18072;
wire            n18073;
wire            n18074;
wire            n18075;
wire            n18076;
wire            n18077;
wire            n18078;
wire            n18079;
wire            n18080;
wire            n18081;
wire            n18082;
wire            n18083;
wire            n18084;
wire            n18085;
wire            n18086;
wire            n18087;
wire            n18088;
wire            n18089;
wire            n18090;
wire            n18091;
wire            n18092;
wire            n18093;
wire            n18094;
wire            n18095;
wire            n18096;
wire            n18097;
wire            n18098;
wire            n18099;
wire            n18100;
wire            n18101;
wire            n18102;
wire            n18103;
wire            n18104;
wire            n18105;
wire            n18106;
wire            n18107;
wire            n18108;
wire            n18109;
wire            n18110;
wire            n18111;
wire            n18112;
wire            n18113;
wire            n18114;
wire            n18115;
wire            n18116;
wire            n18117;
wire            n18118;
wire            n18119;
wire            n18120;
wire            n18121;
wire            n18122;
wire            n18123;
wire            n18124;
wire            n18125;
wire            n18126;
wire            n18127;
wire            n18128;
wire            n18129;
wire            n18130;
wire            n18131;
wire            n18132;
wire            n18133;
wire            n18134;
wire            n18135;
wire            n18136;
wire            n18137;
wire            n18138;
wire            n18139;
wire            n18140;
wire            n18141;
wire            n18142;
wire            n18143;
wire            n18144;
wire            n18145;
wire            n18146;
wire            n18147;
wire            n18148;
wire            n18149;
wire            n18150;
wire            n18151;
wire            n18152;
wire            n18153;
wire            n18154;
wire            n18155;
wire            n18156;
wire            n18157;
wire            n18158;
wire            n18159;
wire            n18160;
wire            n18161;
wire            n18162;
wire            n18163;
wire            n18164;
wire            n18165;
wire            n18166;
wire            n18167;
wire            n18168;
wire            n18169;
wire            n18170;
wire            n18171;
wire            n18172;
wire            n18173;
wire            n18174;
wire            n18175;
wire            n18176;
wire            n18177;
wire            n18178;
wire            n18179;
wire            n18180;
wire            n18181;
wire            n18182;
wire            n18183;
wire            n18184;
wire            n18185;
wire            n18186;
wire            n18187;
wire            n18188;
wire            n18189;
wire            n18190;
wire            n18191;
wire            n18192;
wire            n18193;
wire            n18194;
wire            n18195;
wire            n18196;
wire            n18197;
wire            n18198;
wire            n18199;
wire            n18200;
wire            n18201;
wire            n18202;
wire            n18203;
wire            n18204;
wire            n18205;
wire            n18206;
wire            n18207;
wire            n18208;
wire            n18209;
wire            n18210;
wire            n18211;
wire            n18212;
wire            n18213;
wire            n18214;
wire            n18215;
wire            n18216;
wire            n18217;
wire            n18218;
wire            n18219;
wire            n18220;
wire            n18221;
wire            n18222;
wire            n18223;
wire            n18224;
wire            n18225;
wire            n18226;
wire            n18227;
wire            n18228;
wire            n18229;
wire            n18230;
wire            n18231;
wire            n18232;
wire            n18233;
wire            n18234;
wire            n18235;
wire            n18236;
wire            n18237;
wire            n18238;
wire            n18239;
wire            n18240;
wire            n18241;
wire            n18242;
wire            n18243;
wire            n18244;
wire            n18245;
wire            n18246;
wire            n18247;
wire            n18248;
wire            n18249;
wire            n18250;
wire            n18251;
wire            n18252;
wire            n18253;
wire            n18254;
wire            n18255;
wire            n18256;
wire            n18257;
wire            n18258;
wire            n18259;
wire            n18260;
wire            n18261;
wire            n18262;
wire            n18263;
wire            n18264;
wire            n18265;
wire            n18266;
wire            n18267;
wire            n18268;
wire            n18269;
wire            n18270;
wire            n18271;
wire            n18272;
wire            n18273;
wire            n18274;
wire            n18275;
wire            n18276;
wire            n18277;
wire            n18278;
wire            n18279;
wire            n18280;
wire            n18281;
wire            n18282;
wire            n18283;
wire            n18284;
wire            n18285;
wire            n18286;
wire            n18287;
wire            n18288;
wire            n18289;
wire            n18290;
wire            n18291;
wire            n18292;
wire            n18293;
wire            n18294;
wire            n18295;
wire            n18296;
wire            n18297;
wire            n18298;
wire            n18299;
wire            n18300;
wire            n18301;
wire            n18302;
wire            n18303;
wire            n18304;
wire            n18305;
wire            n18306;
wire            n18307;
wire            n18308;
wire            n18309;
wire            n18310;
wire            n18311;
wire            n18312;
wire            n18313;
wire            n18314;
wire            n18315;
wire            n18316;
wire            n18317;
wire            n18318;
wire            n18319;
wire            n18320;
wire            n18321;
wire            n18322;
wire            n18323;
wire            n18324;
wire            n18325;
wire            n18326;
wire            n18327;
wire            n18328;
wire            n18329;
wire            n18330;
wire            n18331;
wire            n18332;
wire            n18333;
wire            n18334;
wire            n18335;
wire            n18336;
wire            n18337;
wire            n18338;
wire            n18339;
wire            n18340;
wire            n18341;
wire            n18342;
wire            n18343;
wire            n18344;
wire            n18345;
wire            n18346;
wire            n18347;
wire            n18348;
wire            n18349;
wire            n18350;
wire            n18351;
wire            n18352;
wire            n18353;
wire            n18354;
wire            n18355;
wire            n18356;
wire            n18357;
wire            n18358;
wire            n18359;
wire            n18360;
wire            n18361;
wire            n18362;
wire            n18363;
wire            n18364;
wire            n18365;
wire            n18366;
wire            n18367;
wire            n18368;
wire            n18369;
wire            n18370;
wire            n18371;
wire            n18372;
wire            n18373;
wire            n18374;
wire            n18375;
wire            n18376;
wire            n18377;
wire            n18378;
wire            n18379;
wire            n18380;
wire            n18381;
wire            n18382;
wire            n18383;
wire            n18384;
wire            n18385;
wire            n18386;
wire            n18387;
wire            n18388;
wire            n18389;
wire            n18390;
wire            n18391;
wire            n18392;
wire            n18393;
wire            n18394;
wire            n18395;
wire            n18396;
wire            n18397;
wire            n18398;
wire            n18399;
wire            n18400;
wire            n18401;
wire            n18402;
wire            n18403;
wire            n18404;
wire            n18405;
wire            n18406;
wire            n18407;
wire            n18408;
wire            n18409;
wire            n18410;
wire            n18411;
wire            n18412;
wire            n18413;
wire            n18414;
wire            n18415;
wire            n18416;
wire            n18417;
wire            n18418;
wire            n18419;
wire            n18420;
wire            n18421;
wire            n18422;
wire            n18423;
wire            n18424;
wire            n18425;
wire            n18426;
wire            n18427;
wire            n18428;
wire            n18429;
wire     [31:0] n18430;
wire     [31:0] n18431;
wire     [31:0] n18432;
wire     [31:0] n18433;
wire     [31:0] n18434;
wire     [31:0] n18435;
wire     [31:0] n18436;
wire     [31:0] n18437;
wire     [31:0] n18438;
wire     [31:0] n18439;
wire     [31:0] n18440;
wire     [31:0] n18441;
wire     [31:0] n18442;
wire     [31:0] n18443;
wire     [31:0] n18444;
wire     [31:0] n18445;
wire     [31:0] n18446;
wire     [31:0] n18447;
wire     [31:0] n18448;
wire     [31:0] n18449;
wire     [31:0] n18450;
wire     [31:0] n18451;
wire     [31:0] n18452;
wire     [31:0] n18453;
wire     [31:0] n18454;
wire     [31:0] n18455;
wire     [31:0] n18456;
wire     [31:0] n18457;
wire     [31:0] n18458;
wire     [31:0] n18459;
wire     [31:0] n18460;
wire     [31:0] n18461;
wire     [31:0] n18462;
wire     [31:0] n18463;
wire     [31:0] n18464;
wire     [31:0] n18465;
wire     [31:0] n18466;
wire     [31:0] n18467;
wire     [31:0] n18468;
wire     [31:0] n18469;
wire     [31:0] n18470;
wire     [31:0] n18471;
wire     [31:0] n18472;
wire     [31:0] n18473;
wire     [31:0] n18474;
wire     [31:0] n18475;
wire     [31:0] n18476;
wire     [31:0] n18477;
wire     [31:0] n18478;
wire     [31:0] n18479;
wire     [31:0] n18480;
wire     [31:0] n18481;
wire     [31:0] n18482;
wire     [31:0] n18483;
wire     [31:0] n18484;
wire     [31:0] n18485;
wire     [31:0] n18486;
wire     [31:0] n18487;
wire     [31:0] n18488;
wire     [31:0] n18489;
wire     [31:0] n18490;
wire     [31:0] n18491;
wire     [31:0] n18492;
wire     [31:0] n18493;
wire     [31:0] n18494;
wire     [31:0] n18495;
wire     [31:0] n18496;
wire     [31:0] n18497;
wire     [31:0] n18498;
wire     [31:0] n18499;
wire     [31:0] n18500;
wire     [31:0] n18501;
wire     [31:0] n18502;
wire     [31:0] n18503;
wire     [31:0] n18504;
wire     [31:0] n18505;
wire     [31:0] n18506;
wire     [31:0] n18507;
wire     [31:0] n18508;
wire     [31:0] n18509;
wire     [31:0] n18510;
wire     [31:0] n18511;
wire     [31:0] n18512;
wire     [31:0] n18513;
wire     [31:0] n18514;
wire     [31:0] n18515;
wire     [31:0] n18516;
wire     [31:0] n18517;
wire     [31:0] n18518;
wire     [31:0] n18519;
wire     [31:0] n18520;
wire     [31:0] n18521;
wire     [31:0] n18522;
wire     [31:0] n18523;
wire     [31:0] n18524;
wire     [31:0] n18525;
wire     [31:0] n18526;
wire     [31:0] n18527;
wire     [31:0] n18528;
wire     [31:0] n18529;
wire     [31:0] n18530;
wire     [31:0] n18531;
wire     [31:0] n18532;
wire     [31:0] n18533;
wire     [31:0] n18534;
wire     [31:0] n18535;
wire     [31:0] n18536;
wire     [31:0] n18537;
wire     [31:0] n18538;
wire     [31:0] n18539;
wire     [31:0] n18540;
wire     [31:0] n18541;
wire     [31:0] n18542;
wire     [31:0] n18543;
wire     [31:0] n18544;
wire     [31:0] n18545;
wire     [31:0] n18546;
wire     [31:0] n18547;
wire     [31:0] n18548;
wire     [31:0] n18549;
wire     [31:0] n18550;
wire     [31:0] n18551;
wire     [31:0] n18552;
wire     [31:0] n18553;
wire     [31:0] n18554;
wire     [31:0] n18555;
wire     [31:0] n18556;
wire     [31:0] n18557;
wire     [31:0] n18558;
wire     [31:0] n18559;
wire     [31:0] n18560;
wire     [31:0] n18561;
wire     [31:0] n18562;
wire     [31:0] n18563;
wire     [31:0] n18564;
wire     [31:0] n18565;
wire     [31:0] n18566;
wire     [31:0] n18567;
wire     [31:0] n18568;
wire     [31:0] n18569;
wire     [31:0] n18570;
wire     [31:0] n18571;
wire     [31:0] n18572;
wire     [31:0] n18573;
wire     [31:0] n18574;
wire     [31:0] n18575;
wire     [31:0] n18576;
wire     [31:0] n18577;
wire     [31:0] n18578;
wire     [31:0] n18579;
wire     [31:0] n18580;
wire     [31:0] n18581;
wire     [31:0] n18582;
wire     [31:0] n18583;
wire     [31:0] n18584;
wire     [31:0] n18585;
wire     [31:0] n18586;
wire     [31:0] n18587;
wire     [31:0] n18588;
wire     [31:0] n18589;
wire     [31:0] n18590;
wire     [31:0] n18591;
wire     [31:0] n18592;
wire     [31:0] n18593;
wire     [31:0] n18594;
wire     [31:0] n18595;
wire     [31:0] n18596;
wire     [31:0] n18597;
wire     [31:0] n18598;
wire     [31:0] n18599;
wire     [31:0] n18600;
wire     [31:0] n18601;
wire     [31:0] n18602;
wire     [31:0] n18603;
wire     [31:0] n18604;
wire     [31:0] n18605;
wire     [31:0] n18606;
wire     [31:0] n18607;
wire     [31:0] n18608;
wire     [31:0] n18609;
wire     [31:0] n18610;
wire     [31:0] n18611;
wire     [31:0] n18612;
wire     [31:0] n18613;
wire     [31:0] n18614;
wire     [31:0] n18615;
wire     [31:0] n18616;
wire     [31:0] n18617;
wire     [31:0] n18618;
wire     [31:0] n18619;
wire     [31:0] n18620;
wire     [31:0] n18621;
wire     [31:0] n18622;
wire     [31:0] n18623;
wire     [31:0] n18624;
wire     [31:0] n18625;
wire     [31:0] n18626;
wire     [31:0] n18627;
wire     [31:0] n18628;
wire     [31:0] n18629;
wire     [31:0] n18630;
wire     [31:0] n18631;
wire     [31:0] n18632;
wire     [31:0] n18633;
wire     [31:0] n18634;
wire     [31:0] n18635;
wire     [31:0] n18636;
wire     [31:0] n18637;
wire     [31:0] n18638;
wire     [31:0] n18639;
wire     [31:0] n18640;
wire     [31:0] n18641;
wire     [31:0] n18642;
wire     [31:0] n18643;
wire     [31:0] n18644;
wire     [31:0] n18645;
wire     [31:0] n18646;
wire     [31:0] n18647;
wire     [31:0] n18648;
wire     [31:0] n18649;
wire     [31:0] n18650;
wire     [31:0] n18651;
wire     [31:0] n18652;
wire     [31:0] n18653;
wire     [31:0] n18654;
wire     [31:0] n18655;
wire     [31:0] n18656;
wire     [31:0] n18657;
wire     [31:0] n18658;
wire     [31:0] n18659;
wire     [31:0] n18660;
wire     [31:0] n18661;
wire     [31:0] n18662;
wire     [31:0] n18663;
wire     [31:0] n18664;
wire     [31:0] n18665;
wire     [31:0] n18666;
wire     [31:0] n18667;
wire     [31:0] n18668;
wire     [31:0] n18669;
wire     [31:0] n18670;
wire     [31:0] n18671;
wire     [31:0] n18672;
wire     [31:0] n18673;
wire     [31:0] n18674;
wire     [31:0] n18675;
wire     [31:0] n18676;
wire     [31:0] n18677;
wire     [31:0] n18678;
wire     [31:0] n18679;
wire     [31:0] n18680;
wire     [31:0] n18681;
wire     [31:0] n18682;
wire     [31:0] n18683;
wire     [31:0] n18684;
wire     [31:0] n18685;
wire     [31:0] n18686;
wire     [31:0] n18687;
wire     [31:0] n18688;
wire     [31:0] n18689;
wire     [31:0] n18690;
wire     [31:0] n18691;
wire     [31:0] n18692;
wire     [31:0] n18693;
wire     [31:0] n18694;
wire     [31:0] n18695;
wire     [31:0] n18696;
wire     [31:0] n18697;
wire     [31:0] n18698;
wire     [31:0] n18699;
wire     [31:0] n18700;
wire     [31:0] n18701;
wire     [31:0] n18702;
wire     [31:0] n18703;
wire     [31:0] n18704;
wire     [31:0] n18705;
wire     [31:0] n18706;
wire     [31:0] n18707;
wire     [31:0] n18708;
wire     [31:0] n18709;
wire     [31:0] n18710;
wire     [31:0] n18711;
wire     [31:0] n18712;
wire     [31:0] n18713;
wire     [31:0] n18714;
wire     [31:0] n18715;
wire     [31:0] n18716;
wire     [31:0] n18717;
wire     [31:0] n18718;
wire     [31:0] n18719;
wire     [31:0] n18720;
wire     [31:0] n18721;
wire     [31:0] n18722;
wire     [31:0] n18723;
wire     [31:0] n18724;
wire     [31:0] n18725;
wire     [31:0] n18726;
wire     [31:0] n18727;
wire     [31:0] n18728;
wire     [31:0] n18729;
wire     [31:0] n18730;
wire     [31:0] n18731;
wire     [31:0] n18732;
wire     [31:0] n18733;
wire     [31:0] n18734;
wire     [31:0] n18735;
wire     [31:0] n18736;
wire     [31:0] n18737;
wire     [31:0] n18738;
wire     [31:0] n18739;
wire     [31:0] n18740;
wire     [31:0] n18741;
wire     [31:0] n18742;
wire     [31:0] n18743;
wire     [31:0] n18744;
wire     [31:0] n18745;
wire     [31:0] n18746;
wire     [31:0] n18747;
wire     [31:0] n18748;
wire     [31:0] n18749;
wire     [31:0] n18750;
wire     [31:0] n18751;
wire     [31:0] n18752;
wire     [31:0] n18753;
wire     [31:0] n18754;
wire     [31:0] n18755;
wire     [31:0] n18756;
wire     [31:0] n18757;
wire     [31:0] n18758;
wire     [31:0] n18759;
wire     [31:0] n18760;
wire     [31:0] n18761;
wire     [31:0] n18762;
wire     [31:0] n18763;
wire     [31:0] n18764;
wire     [31:0] n18765;
wire     [31:0] n18766;
wire     [31:0] n18767;
wire     [31:0] n18768;
wire     [31:0] n18769;
wire     [31:0] n18770;
wire     [31:0] n18771;
wire     [31:0] n18772;
wire     [31:0] n18773;
wire     [31:0] n18774;
wire     [31:0] n18775;
wire     [31:0] n18776;
wire     [31:0] n18777;
wire     [31:0] n18778;
wire     [31:0] n18779;
wire     [31:0] n18780;
wire     [31:0] n18781;
wire     [31:0] n18782;
wire     [31:0] n18783;
wire     [31:0] n18784;
wire     [31:0] n18785;
wire     [31:0] n18786;
wire     [31:0] n18787;
wire     [31:0] n18788;
wire     [31:0] n18789;
wire     [31:0] n18790;
wire     [31:0] n18791;
wire     [31:0] n18792;
wire     [31:0] n18793;
wire     [31:0] n18794;
wire     [31:0] n18795;
wire     [31:0] n18796;
wire     [31:0] n18797;
wire     [31:0] n18798;
wire     [31:0] n18799;
wire     [31:0] n18800;
wire     [31:0] n18801;
wire     [31:0] n18802;
wire     [31:0] n18803;
wire     [31:0] n18804;
wire     [31:0] n18805;
wire     [31:0] n18806;
wire     [31:0] n18807;
wire     [31:0] n18808;
wire     [31:0] n18809;
wire     [31:0] n18810;
wire     [31:0] n18811;
wire     [31:0] n18812;
wire     [31:0] n18813;
wire     [31:0] n18814;
wire     [31:0] n18815;
wire     [31:0] n18816;
wire     [31:0] n18817;
wire     [31:0] n18818;
wire     [31:0] n18819;
wire     [31:0] n18820;
wire     [31:0] n18821;
wire     [31:0] n18822;
wire     [31:0] n18823;
wire     [31:0] n18824;
wire     [31:0] n18825;
wire     [31:0] n18826;
wire     [31:0] n18827;
wire     [31:0] n18828;
wire     [31:0] n18829;
wire     [31:0] n18830;
wire     [31:0] n18831;
wire     [31:0] n18832;
wire     [31:0] n18833;
wire     [31:0] n18834;
wire     [31:0] n18835;
wire     [31:0] n18836;
wire     [31:0] n18837;
wire     [31:0] n18838;
wire     [31:0] n18839;
wire     [31:0] n18840;
wire     [31:0] n18841;
wire     [31:0] n18842;
wire     [31:0] n18843;
wire     [31:0] n18844;
wire     [31:0] n18845;
wire     [31:0] n18846;
wire     [31:0] n18847;
wire     [31:0] n18848;
wire     [31:0] n18849;
wire     [31:0] n18850;
wire     [31:0] n18851;
wire     [31:0] n18852;
wire     [31:0] n18853;
wire     [31:0] n18854;
wire     [31:0] n18855;
wire     [31:0] n18856;
wire     [31:0] n18857;
wire     [31:0] n18858;
wire     [31:0] n18859;
wire     [31:0] n18860;
wire     [31:0] n18861;
wire     [31:0] n18862;
wire     [31:0] n18863;
wire     [31:0] n18864;
wire     [31:0] n18865;
wire     [31:0] n18866;
wire     [31:0] n18867;
wire     [31:0] n18868;
wire     [31:0] n18869;
wire     [31:0] n18870;
wire     [31:0] n18871;
wire     [31:0] n18872;
wire     [31:0] n18873;
wire     [31:0] n18874;
wire     [31:0] n18875;
wire     [31:0] n18876;
wire     [31:0] n18877;
wire     [31:0] n18878;
wire     [31:0] n18879;
wire     [31:0] n18880;
wire     [31:0] n18881;
wire     [31:0] n18882;
wire     [31:0] n18883;
wire     [31:0] n18884;
wire     [31:0] n18885;
wire     [31:0] n18886;
wire     [31:0] n18887;
wire     [31:0] n18888;
wire     [31:0] n18889;
wire     [31:0] n18890;
wire     [31:0] n18891;
wire     [31:0] n18892;
wire     [31:0] n18893;
wire     [31:0] n18894;
wire     [31:0] n18895;
wire     [31:0] n18896;
wire     [31:0] n18897;
wire     [31:0] n18898;
wire     [31:0] n18899;
wire     [31:0] n18900;
wire     [31:0] n18901;
wire     [31:0] n18902;
wire     [31:0] n18903;
wire     [31:0] n18904;
wire     [31:0] n18905;
wire     [31:0] n18906;
wire     [31:0] n18907;
wire     [31:0] n18908;
wire     [31:0] n18909;
wire     [31:0] n18910;
wire     [31:0] n18911;
wire     [31:0] n18912;
wire     [31:0] n18913;
wire     [31:0] n18914;
wire     [31:0] n18915;
wire     [31:0] n18916;
wire     [31:0] n18917;
wire     [31:0] n18918;
wire     [31:0] n18919;
wire     [31:0] n18920;
wire     [31:0] n18921;
wire     [31:0] n18922;
wire     [31:0] n18923;
wire     [31:0] n18924;
wire     [31:0] n18925;
wire     [31:0] n18926;
wire     [31:0] n18927;
wire     [31:0] n18928;
wire     [31:0] n18929;
wire     [31:0] n18930;
wire     [31:0] n18931;
wire     [31:0] n18932;
wire     [31:0] n18933;
wire     [31:0] n18934;
wire     [31:0] n18935;
wire     [31:0] n18936;
wire     [31:0] n18937;
wire     [31:0] n18938;
wire     [31:0] n18939;
wire     [31:0] n18940;
wire     [31:0] n18941;
wire     [31:0] n18942;
wire     [31:0] n18943;
wire     [31:0] n18944;
wire     [31:0] n18945;
wire     [31:0] n18946;
wire     [31:0] n18947;
wire     [31:0] n18948;
wire     [31:0] n18949;
wire     [31:0] n18950;
wire     [31:0] n18951;
wire            n18952;
wire            n18953;
wire            n18954;
wire            n18955;
wire            n18956;
wire            n18957;
wire            n18958;
wire            n18959;
wire            n18960;
wire            n18961;
wire            n18962;
wire            n18963;
wire            n18964;
wire            n18965;
wire            n18966;
wire            n18967;
wire            n18968;
wire            n18969;
wire            n18970;
wire            n18971;
wire            n18972;
wire            n18973;
wire            n18974;
wire            n18975;
wire            n18976;
wire            n18977;
wire            n18978;
wire            n18979;
wire            n18980;
wire            n18981;
wire            n18982;
wire            n18983;
wire            n18984;
wire            n18985;
wire            n18986;
wire            n18987;
wire            n18988;
wire            n18989;
wire            n18990;
wire            n18991;
wire            n18992;
wire            n18993;
wire            n18994;
wire            n18995;
wire            n18996;
wire            n18997;
wire            n18998;
wire            n18999;
wire            n19000;
wire            n19001;
wire            n19002;
wire            n19003;
wire            n19004;
wire            n19005;
wire            n19006;
wire            n19007;
wire            n19008;
wire            n19009;
wire            n19010;
wire            n19011;
wire            n19012;
wire            n19013;
wire            n19014;
wire            n19015;
wire            n19016;
wire            n19017;
wire            n19018;
wire            n19019;
wire            n19020;
wire            n19021;
wire            n19022;
wire            n19023;
wire            n19024;
wire            n19025;
wire            n19026;
wire            n19027;
wire            n19028;
wire            n19029;
wire            n19030;
wire            n19031;
wire            n19032;
wire            n19033;
wire            n19034;
wire            n19035;
wire            n19036;
wire            n19037;
wire            n19038;
wire            n19039;
wire            n19040;
wire            n19041;
wire            n19042;
wire            n19043;
wire            n19044;
wire            n19045;
wire            n19046;
wire            n19047;
wire            n19048;
wire            n19049;
wire            n19050;
wire            n19051;
wire            n19052;
wire            n19053;
wire            n19054;
wire            n19055;
wire            n19056;
wire            n19057;
wire            n19058;
wire            n19059;
wire            n19060;
wire            n19061;
wire            n19062;
wire            n19063;
wire            n19064;
wire            n19065;
wire            n19066;
wire            n19067;
wire            n19068;
wire            n19069;
wire            n19070;
wire            n19071;
wire            n19072;
wire            n19073;
wire            n19074;
wire            n19075;
wire            n19076;
wire            n19077;
wire            n19078;
wire            n19079;
wire            n19080;
wire            n19081;
wire            n19082;
wire            n19083;
wire            n19084;
wire            n19085;
wire            n19086;
wire            n19087;
wire            n19088;
wire            n19089;
wire            n19090;
wire            n19091;
wire            n19092;
wire            n19093;
wire            n19094;
wire            n19095;
wire            n19096;
wire            n19097;
wire            n19098;
wire            n19099;
wire            n19100;
wire            n19101;
wire            n19102;
wire            n19103;
wire            n19104;
wire            n19105;
wire            n19106;
wire            n19107;
wire            n19108;
wire            n19109;
wire            n19110;
wire            n19111;
wire            n19112;
wire            n19113;
wire            n19114;
wire            n19115;
wire            n19116;
wire            n19117;
wire            n19118;
wire            n19119;
wire            n19120;
wire            n19121;
wire            n19122;
wire            n19123;
wire            n19124;
wire            n19125;
wire            n19126;
wire            n19127;
wire            n19128;
wire            n19129;
wire            n19130;
wire            n19131;
wire            n19132;
wire            n19133;
wire            n19134;
wire            n19135;
wire            n19136;
wire            n19137;
wire            n19138;
wire            n19139;
wire            n19140;
wire            n19141;
wire            n19142;
wire            n19143;
wire            n19144;
wire            n19145;
wire            n19146;
wire            n19147;
wire            n19148;
wire            n19149;
wire            n19150;
wire            n19151;
wire            n19152;
wire            n19153;
wire            n19154;
wire            n19155;
wire            n19156;
wire            n19157;
wire            n19158;
wire            n19159;
wire            n19160;
wire            n19161;
wire            n19162;
wire            n19163;
wire            n19164;
wire            n19165;
wire            n19166;
wire            n19167;
wire            n19168;
wire            n19169;
wire            n19170;
wire            n19171;
wire            n19172;
wire            n19173;
wire            n19174;
wire            n19175;
wire            n19176;
wire            n19177;
wire            n19178;
wire            n19179;
wire            n19180;
wire            n19181;
wire            n19182;
wire            n19183;
wire            n19184;
wire            n19185;
wire            n19186;
wire            n19187;
wire            n19188;
wire            n19189;
wire            n19190;
wire            n19191;
wire            n19192;
wire            n19193;
wire            n19194;
wire            n19195;
wire            n19196;
wire            n19197;
wire            n19198;
wire            n19199;
wire            n19200;
wire            n19201;
wire            n19202;
wire            n19203;
wire            n19204;
wire            n19205;
wire            n19206;
wire            n19207;
wire            n19208;
wire            n19209;
wire            n19210;
wire            n19211;
wire            n19212;
wire            n19213;
wire            n19214;
wire            n19215;
wire            n19216;
wire            n19217;
wire            n19218;
wire            n19219;
wire            n19220;
wire            n19221;
wire            n19222;
wire            n19223;
wire            n19224;
wire            n19225;
wire            n19226;
wire            n19227;
wire            n19228;
wire            n19229;
wire            n19230;
wire            n19231;
wire            n19232;
wire            n19233;
wire            n19234;
wire            n19235;
wire            n19236;
wire            n19237;
wire            n19238;
wire            n19239;
wire            n19240;
wire            n19241;
wire            n19242;
wire            n19243;
wire            n19244;
wire            n19245;
wire            n19246;
wire            n19247;
wire            n19248;
wire            n19249;
wire            n19250;
wire            n19251;
wire            n19252;
wire            n19253;
wire            n19254;
wire            n19255;
wire            n19256;
wire            n19257;
wire            n19258;
wire            n19259;
wire            n19260;
wire            n19261;
wire            n19262;
wire            n19263;
wire            n19264;
wire            n19265;
wire            n19266;
wire            n19267;
wire            n19268;
wire            n19269;
wire            n19270;
wire            n19271;
wire            n19272;
wire            n19273;
wire            n19274;
wire            n19275;
wire            n19276;
wire            n19277;
wire            n19278;
wire            n19279;
wire            n19280;
wire            n19281;
wire            n19282;
wire            n19283;
wire            n19284;
wire            n19285;
wire            n19286;
wire            n19287;
wire            n19288;
wire            n19289;
wire            n19290;
wire            n19291;
wire            n19292;
wire            n19293;
wire            n19294;
wire            n19295;
wire            n19296;
wire            n19297;
wire            n19298;
wire            n19299;
wire            n19300;
wire            n19301;
wire            n19302;
wire            n19303;
wire            n19304;
wire            n19305;
wire            n19306;
wire            n19307;
wire            n19308;
wire            n19309;
wire            n19310;
wire            n19311;
wire            n19312;
wire            n19313;
wire            n19314;
wire            n19315;
wire            n19316;
wire            n19317;
wire            n19318;
wire            n19319;
wire            n19320;
wire            n19321;
wire            n19322;
wire            n19323;
wire            n19324;
wire            n19325;
wire            n19326;
wire            n19327;
wire            n19328;
wire            n19329;
wire            n19330;
wire            n19331;
wire            n19332;
wire            n19333;
wire            n19334;
wire            n19335;
wire            n19336;
wire            n19337;
wire            n19338;
wire            n19339;
wire            n19340;
wire            n19341;
wire            n19342;
wire            n19343;
wire            n19344;
wire            n19345;
wire            n19346;
wire            n19347;
wire            n19348;
wire            n19349;
wire            n19350;
wire            n19351;
wire            n19352;
wire            n19353;
wire            n19354;
wire            n19355;
wire            n19356;
wire            n19357;
wire            n19358;
wire            n19359;
wire            n19360;
wire            n19361;
wire            n19362;
wire            n19363;
wire            n19364;
wire            n19365;
wire            n19366;
wire            n19367;
wire            n19368;
wire            n19369;
wire            n19370;
wire            n19371;
wire            n19372;
wire            n19373;
wire            n19374;
wire            n19375;
wire            n19376;
wire            n19377;
wire            n19378;
wire            n19379;
wire            n19380;
wire            n19381;
wire            n19382;
wire            n19383;
wire            n19384;
wire            n19385;
wire            n19386;
wire            n19387;
wire            n19388;
wire            n19389;
wire            n19390;
wire            n19391;
wire            n19392;
wire            n19393;
wire            n19394;
wire            n19395;
wire            n19396;
wire            n19397;
wire            n19398;
wire            n19399;
wire            n19400;
wire            n19401;
wire            n19402;
wire            n19403;
wire            n19404;
wire            n19405;
wire            n19406;
wire            n19407;
wire            n19408;
wire            n19409;
wire            n19410;
wire            n19411;
wire            n19412;
wire            n19413;
wire            n19414;
wire            n19415;
wire            n19416;
wire            n19417;
wire            n19418;
wire            n19419;
wire            n19420;
wire            n19421;
wire            n19422;
wire            n19423;
wire            n19424;
wire            n19425;
wire            n19426;
wire            n19427;
wire            n19428;
wire            n19429;
wire            n19430;
wire            n19431;
wire            n19432;
wire            n19433;
wire            n19434;
wire            n19435;
wire            n19436;
wire            n19437;
wire            n19438;
wire            n19439;
wire            n19440;
wire            n19441;
wire            n19442;
wire            n19443;
wire            n19444;
wire            n19445;
wire            n19446;
wire            n19447;
wire            n19448;
wire            n19449;
wire            n19450;
wire            n19451;
wire            n19452;
wire            n19453;
wire            n19454;
wire            n19455;
wire            n19456;
wire            n19457;
wire            n19458;
wire            n19459;
wire            n19460;
wire            n19461;
wire            n19462;
wire            n19463;
wire     [31:0] n19464;
wire     [31:0] n19465;
wire     [31:0] n19466;
wire     [31:0] n19467;
wire     [31:0] n19468;
wire     [31:0] n19469;
wire     [31:0] n19470;
wire     [31:0] n19471;
wire     [31:0] n19472;
wire     [31:0] n19473;
wire     [31:0] n19474;
wire     [31:0] n19475;
wire     [31:0] n19476;
wire     [31:0] n19477;
wire     [31:0] n19478;
wire     [31:0] n19479;
wire     [31:0] n19480;
wire     [31:0] n19481;
wire     [31:0] n19482;
wire     [31:0] n19483;
wire     [31:0] n19484;
wire     [31:0] n19485;
wire     [31:0] n19486;
wire     [31:0] n19487;
wire     [31:0] n19488;
wire     [31:0] n19489;
wire     [31:0] n19490;
wire     [31:0] n19491;
wire     [31:0] n19492;
wire     [31:0] n19493;
wire     [31:0] n19494;
wire     [31:0] n19495;
wire     [31:0] n19496;
wire     [31:0] n19497;
wire     [31:0] n19498;
wire     [31:0] n19499;
wire     [31:0] n19500;
wire     [31:0] n19501;
wire     [31:0] n19502;
wire     [31:0] n19503;
wire     [31:0] n19504;
wire     [31:0] n19505;
wire     [31:0] n19506;
wire     [31:0] n19507;
wire     [31:0] n19508;
wire     [31:0] n19509;
wire     [31:0] n19510;
wire     [31:0] n19511;
wire     [31:0] n19512;
wire     [31:0] n19513;
wire     [31:0] n19514;
wire     [31:0] n19515;
wire     [31:0] n19516;
wire     [31:0] n19517;
wire     [31:0] n19518;
wire     [31:0] n19519;
wire     [31:0] n19520;
wire     [31:0] n19521;
wire     [31:0] n19522;
wire     [31:0] n19523;
wire     [31:0] n19524;
wire     [31:0] n19525;
wire     [31:0] n19526;
wire     [31:0] n19527;
wire     [31:0] n19528;
wire     [31:0] n19529;
wire     [31:0] n19530;
wire     [31:0] n19531;
wire     [31:0] n19532;
wire     [31:0] n19533;
wire     [31:0] n19534;
wire     [31:0] n19535;
wire     [31:0] n19536;
wire     [31:0] n19537;
wire     [31:0] n19538;
wire     [31:0] n19539;
wire     [31:0] n19540;
wire     [31:0] n19541;
wire     [31:0] n19542;
wire     [31:0] n19543;
wire     [31:0] n19544;
wire     [31:0] n19545;
wire     [31:0] n19546;
wire     [31:0] n19547;
wire     [31:0] n19548;
wire     [31:0] n19549;
wire     [31:0] n19550;
wire     [31:0] n19551;
wire     [31:0] n19552;
wire     [31:0] n19553;
wire     [31:0] n19554;
wire     [31:0] n19555;
wire     [31:0] n19556;
wire     [31:0] n19557;
wire     [31:0] n19558;
wire     [31:0] n19559;
wire     [31:0] n19560;
wire     [31:0] n19561;
wire     [31:0] n19562;
wire     [31:0] n19563;
wire     [31:0] n19564;
wire     [31:0] n19565;
wire     [31:0] n19566;
wire     [31:0] n19567;
wire     [31:0] n19568;
wire     [31:0] n19569;
wire     [31:0] n19570;
wire     [31:0] n19571;
wire     [31:0] n19572;
wire     [31:0] n19573;
wire     [31:0] n19574;
wire     [31:0] n19575;
wire     [31:0] n19576;
wire     [31:0] n19577;
wire     [31:0] n19578;
wire     [31:0] n19579;
wire     [31:0] n19580;
wire     [31:0] n19581;
wire     [31:0] n19582;
wire     [31:0] n19583;
wire     [31:0] n19584;
wire     [31:0] n19585;
wire     [31:0] n19586;
wire     [31:0] n19587;
wire     [31:0] n19588;
wire     [31:0] n19589;
wire     [31:0] n19590;
wire     [31:0] n19591;
wire     [31:0] n19592;
wire     [31:0] n19593;
wire     [31:0] n19594;
wire     [31:0] n19595;
wire     [31:0] n19596;
wire     [31:0] n19597;
wire     [31:0] n19598;
wire     [31:0] n19599;
wire     [31:0] n19600;
wire     [31:0] n19601;
wire     [31:0] n19602;
wire     [31:0] n19603;
wire     [31:0] n19604;
wire     [31:0] n19605;
wire     [31:0] n19606;
wire     [31:0] n19607;
wire     [31:0] n19608;
wire     [31:0] n19609;
wire     [31:0] n19610;
wire     [31:0] n19611;
wire     [31:0] n19612;
wire     [31:0] n19613;
wire     [31:0] n19614;
wire     [31:0] n19615;
wire     [31:0] n19616;
wire     [31:0] n19617;
wire     [31:0] n19618;
wire     [31:0] n19619;
wire     [31:0] n19620;
wire     [31:0] n19621;
wire     [31:0] n19622;
wire     [31:0] n19623;
wire     [31:0] n19624;
wire     [31:0] n19625;
wire     [31:0] n19626;
wire     [31:0] n19627;
wire     [31:0] n19628;
wire     [31:0] n19629;
wire     [31:0] n19630;
wire     [31:0] n19631;
wire     [31:0] n19632;
wire     [31:0] n19633;
wire     [31:0] n19634;
wire     [31:0] n19635;
wire     [31:0] n19636;
wire     [31:0] n19637;
wire     [31:0] n19638;
wire     [31:0] n19639;
wire     [31:0] n19640;
wire     [31:0] n19641;
wire     [31:0] n19642;
wire     [31:0] n19643;
wire     [31:0] n19644;
wire     [31:0] n19645;
wire     [31:0] n19646;
wire     [31:0] n19647;
wire     [31:0] n19648;
wire     [31:0] n19649;
wire     [31:0] n19650;
wire     [31:0] n19651;
wire     [31:0] n19652;
wire     [31:0] n19653;
wire     [31:0] n19654;
wire     [31:0] n19655;
wire     [31:0] n19656;
wire     [31:0] n19657;
wire     [31:0] n19658;
wire     [31:0] n19659;
wire     [31:0] n19660;
wire     [31:0] n19661;
wire     [31:0] n19662;
wire     [31:0] n19663;
wire     [31:0] n19664;
wire     [31:0] n19665;
wire     [31:0] n19666;
wire     [31:0] n19667;
wire     [31:0] n19668;
wire     [31:0] n19669;
wire     [31:0] n19670;
wire     [31:0] n19671;
wire     [31:0] n19672;
wire     [31:0] n19673;
wire     [31:0] n19674;
wire     [31:0] n19675;
wire     [31:0] n19676;
wire     [31:0] n19677;
wire     [31:0] n19678;
wire     [31:0] n19679;
wire     [31:0] n19680;
wire     [31:0] n19681;
wire     [31:0] n19682;
wire     [31:0] n19683;
wire     [31:0] n19684;
wire     [31:0] n19685;
wire     [31:0] n19686;
wire     [31:0] n19687;
wire     [31:0] n19688;
wire     [31:0] n19689;
wire     [31:0] n19690;
wire     [31:0] n19691;
wire     [31:0] n19692;
wire     [31:0] n19693;
wire     [31:0] n19694;
wire     [31:0] n19695;
wire     [31:0] n19696;
wire     [31:0] n19697;
wire     [31:0] n19698;
wire     [31:0] n19699;
wire     [31:0] n19700;
wire     [31:0] n19701;
wire     [31:0] n19702;
wire     [31:0] n19703;
wire     [31:0] n19704;
wire     [31:0] n19705;
wire     [31:0] n19706;
wire     [31:0] n19707;
wire     [31:0] n19708;
wire     [31:0] n19709;
wire     [31:0] n19710;
wire     [31:0] n19711;
wire     [31:0] n19712;
wire     [31:0] n19713;
wire     [31:0] n19714;
wire     [31:0] n19715;
wire     [31:0] n19716;
wire     [31:0] n19717;
wire     [31:0] n19718;
wire     [31:0] n19719;
wire     [31:0] n19720;
wire     [31:0] n19721;
wire     [31:0] n19722;
wire     [31:0] n19723;
wire     [31:0] n19724;
wire     [31:0] n19725;
wire     [31:0] n19726;
wire     [31:0] n19727;
wire     [31:0] n19728;
wire     [31:0] n19729;
wire     [31:0] n19730;
wire     [31:0] n19731;
wire     [31:0] n19732;
wire     [31:0] n19733;
wire     [31:0] n19734;
wire     [31:0] n19735;
wire     [31:0] n19736;
wire     [31:0] n19737;
wire     [31:0] n19738;
wire     [31:0] n19739;
wire     [31:0] n19740;
wire     [31:0] n19741;
wire     [31:0] n19742;
wire     [31:0] n19743;
wire     [31:0] n19744;
wire     [31:0] n19745;
wire     [31:0] n19746;
wire     [31:0] n19747;
wire     [31:0] n19748;
wire     [31:0] n19749;
wire     [31:0] n19750;
wire     [31:0] n19751;
wire     [31:0] n19752;
wire     [31:0] n19753;
wire     [31:0] n19754;
wire     [31:0] n19755;
wire     [31:0] n19756;
wire     [31:0] n19757;
wire     [31:0] n19758;
wire     [31:0] n19759;
wire     [31:0] n19760;
wire     [31:0] n19761;
wire     [31:0] n19762;
wire     [31:0] n19763;
wire     [31:0] n19764;
wire     [31:0] n19765;
wire     [31:0] n19766;
wire     [31:0] n19767;
wire     [31:0] n19768;
wire     [31:0] n19769;
wire     [31:0] n19770;
wire     [31:0] n19771;
wire     [31:0] n19772;
wire     [31:0] n19773;
wire     [31:0] n19774;
wire     [31:0] n19775;
wire     [31:0] n19776;
wire     [31:0] n19777;
wire     [31:0] n19778;
wire     [31:0] n19779;
wire     [31:0] n19780;
wire     [31:0] n19781;
wire     [31:0] n19782;
wire     [31:0] n19783;
wire     [31:0] n19784;
wire     [31:0] n19785;
wire     [31:0] n19786;
wire     [31:0] n19787;
wire     [31:0] n19788;
wire     [31:0] n19789;
wire     [31:0] n19790;
wire     [31:0] n19791;
wire     [31:0] n19792;
wire     [31:0] n19793;
wire     [31:0] n19794;
wire     [31:0] n19795;
wire     [31:0] n19796;
wire     [31:0] n19797;
wire     [31:0] n19798;
wire     [31:0] n19799;
wire     [31:0] n19800;
wire     [31:0] n19801;
wire     [31:0] n19802;
wire     [31:0] n19803;
wire     [31:0] n19804;
wire     [31:0] n19805;
wire     [31:0] n19806;
wire     [31:0] n19807;
wire     [31:0] n19808;
wire     [31:0] n19809;
wire     [31:0] n19810;
wire     [31:0] n19811;
wire     [31:0] n19812;
wire     [31:0] n19813;
wire     [31:0] n19814;
wire     [31:0] n19815;
wire     [31:0] n19816;
wire     [31:0] n19817;
wire     [31:0] n19818;
wire     [31:0] n19819;
wire     [31:0] n19820;
wire     [31:0] n19821;
wire     [31:0] n19822;
wire     [31:0] n19823;
wire     [31:0] n19824;
wire     [31:0] n19825;
wire     [31:0] n19826;
wire     [31:0] n19827;
wire     [31:0] n19828;
wire     [31:0] n19829;
wire     [31:0] n19830;
wire     [31:0] n19831;
wire     [31:0] n19832;
wire     [31:0] n19833;
wire     [31:0] n19834;
wire     [31:0] n19835;
wire     [31:0] n19836;
wire     [31:0] n19837;
wire     [31:0] n19838;
wire     [31:0] n19839;
wire     [31:0] n19840;
wire     [31:0] n19841;
wire     [31:0] n19842;
wire     [31:0] n19843;
wire     [31:0] n19844;
wire     [31:0] n19845;
wire     [31:0] n19846;
wire     [31:0] n19847;
wire     [31:0] n19848;
wire     [31:0] n19849;
wire     [31:0] n19850;
wire     [31:0] n19851;
wire     [31:0] n19852;
wire     [31:0] n19853;
wire     [31:0] n19854;
wire     [31:0] n19855;
wire     [31:0] n19856;
wire     [31:0] n19857;
wire     [31:0] n19858;
wire     [31:0] n19859;
wire     [31:0] n19860;
wire     [31:0] n19861;
wire     [31:0] n19862;
wire     [31:0] n19863;
wire     [31:0] n19864;
wire     [31:0] n19865;
wire     [31:0] n19866;
wire     [31:0] n19867;
wire     [31:0] n19868;
wire     [31:0] n19869;
wire     [31:0] n19870;
wire     [31:0] n19871;
wire     [31:0] n19872;
wire     [31:0] n19873;
wire     [31:0] n19874;
wire     [31:0] n19875;
wire     [31:0] n19876;
wire     [31:0] n19877;
wire     [31:0] n19878;
wire     [31:0] n19879;
wire     [31:0] n19880;
wire     [31:0] n19881;
wire     [31:0] n19882;
wire     [31:0] n19883;
wire     [31:0] n19884;
wire     [31:0] n19885;
wire     [31:0] n19886;
wire     [31:0] n19887;
wire     [31:0] n19888;
wire     [31:0] n19889;
wire     [31:0] n19890;
wire     [31:0] n19891;
wire     [31:0] n19892;
wire     [31:0] n19893;
wire     [31:0] n19894;
wire     [31:0] n19895;
wire     [31:0] n19896;
wire     [31:0] n19897;
wire     [31:0] n19898;
wire     [31:0] n19899;
wire     [31:0] n19900;
wire     [31:0] n19901;
wire     [31:0] n19902;
wire     [31:0] n19903;
wire     [31:0] n19904;
wire     [31:0] n19905;
wire     [31:0] n19906;
wire     [31:0] n19907;
wire     [31:0] n19908;
wire     [31:0] n19909;
wire     [31:0] n19910;
wire     [31:0] n19911;
wire     [31:0] n19912;
wire     [31:0] n19913;
wire     [31:0] n19914;
wire     [31:0] n19915;
wire     [31:0] n19916;
wire     [31:0] n19917;
wire     [31:0] n19918;
wire     [31:0] n19919;
wire     [31:0] n19920;
wire     [31:0] n19921;
wire     [31:0] n19922;
wire     [31:0] n19923;
wire     [31:0] n19924;
wire     [31:0] n19925;
wire     [31:0] n19926;
wire     [31:0] n19927;
wire     [31:0] n19928;
wire     [31:0] n19929;
wire     [31:0] n19930;
wire     [31:0] n19931;
wire     [31:0] n19932;
wire     [31:0] n19933;
wire     [31:0] n19934;
wire     [31:0] n19935;
wire     [31:0] n19936;
wire     [31:0] n19937;
wire     [31:0] n19938;
wire     [31:0] n19939;
wire     [31:0] n19940;
wire     [31:0] n19941;
wire     [31:0] n19942;
wire     [31:0] n19943;
wire     [31:0] n19944;
wire     [31:0] n19945;
wire     [31:0] n19946;
wire     [31:0] n19947;
wire     [31:0] n19948;
wire     [31:0] n19949;
wire     [31:0] n19950;
wire     [31:0] n19951;
wire     [31:0] n19952;
wire     [31:0] n19953;
wire     [31:0] n19954;
wire     [31:0] n19955;
wire     [31:0] n19956;
wire     [31:0] n19957;
wire     [31:0] n19958;
wire     [31:0] n19959;
wire     [31:0] n19960;
wire     [31:0] n19961;
wire     [31:0] n19962;
wire     [31:0] n19963;
wire     [31:0] n19964;
wire     [31:0] n19965;
wire     [31:0] n19966;
wire     [31:0] n19967;
wire     [31:0] n19968;
wire     [31:0] n19969;
wire     [31:0] n19970;
wire     [31:0] n19971;
wire     [31:0] n19972;
wire     [31:0] n19973;
wire     [31:0] n19974;
wire     [31:0] n19975;
wire     [31:0] n19976;
wire     [31:0] n19977;
wire     [31:0] n19978;
wire     [31:0] n19979;
wire     [31:0] n19980;
wire     [31:0] n19981;
wire     [31:0] n19982;
wire     [31:0] n19983;
wire     [31:0] n19984;
wire     [31:0] n19985;
wire            n19986;
wire            n19987;
wire     [31:0] n19988;
wire     [31:0] n19989;
wire     [31:0] n19990;
wire     [31:0] n19991;
wire     [31:0] n19992;
wire     [31:0] n19993;
wire     [31:0] n19994;
wire     [31:0] n19995;
wire     [31:0] n19996;
wire     [31:0] n19997;
wire     [31:0] n19998;
wire     [31:0] n19999;
wire     [31:0] n20000;
wire     [31:0] n20001;
wire     [31:0] n20002;
wire     [31:0] n20003;
wire     [31:0] n20004;
wire     [31:0] n20005;
wire     [31:0] n20006;
wire     [31:0] n20007;
wire     [31:0] n20008;
wire     [31:0] n20009;
wire     [31:0] n20010;
wire     [31:0] n20011;
wire     [31:0] n20012;
wire     [31:0] n20013;
wire     [31:0] n20014;
wire     [31:0] n20015;
wire     [31:0] n20016;
wire     [31:0] n20017;
wire     [31:0] n20018;
wire     [31:0] n20019;
wire     [31:0] n20020;
wire            n20021;
wire            n20022;
wire            n20023;
wire            n20024;
wire            n20025;
wire            n20026;
wire            n20027;
wire            n20028;
wire            n20029;
wire            n20030;
wire            n20031;
wire            n20032;
wire            n20033;
wire            n20034;
wire            n20035;
wire            n20036;
wire            n20037;
wire            n20038;
wire            n20039;
wire            n20040;
wire            n20041;
wire            n20042;
wire            n20043;
wire            n20044;
wire            n20045;
wire            n20046;
wire            n20047;
wire            n20048;
wire            n20049;
wire            n20050;
wire            n20051;
wire            n20052;
wire            n20053;
wire            n20054;
wire            n20055;
wire            n20056;
wire            n20057;
wire            n20058;
wire            n20059;
wire            n20060;
wire            n20061;
wire            n20062;
wire            n20063;
wire            n20064;
wire            n20065;
wire            n20066;
wire            n20067;
wire            n20068;
wire            n20069;
wire            n20070;
wire            n20071;
wire            n20072;
wire            n20073;
wire            n20074;
wire            n20075;
wire            n20076;
wire            n20077;
wire            n20078;
wire            n20079;
wire            n20080;
wire            n20081;
wire            n20082;
wire            n20083;
wire            n20084;
wire            n20085;
wire            n20086;
wire            n20087;
wire            n20088;
wire            n20089;
wire            n20090;
wire            n20091;
wire            n20092;
wire            n20093;
wire            n20094;
wire            n20095;
wire            n20096;
wire            n20097;
wire            n20098;
wire            n20099;
wire            n20100;
wire            n20101;
wire            n20102;
wire            n20103;
wire            n20104;
wire            n20105;
wire            n20106;
wire            n20107;
wire            n20108;
wire            n20109;
wire            n20110;
wire            n20111;
wire            n20112;
wire            n20113;
wire            n20114;
wire            n20115;
wire            n20116;
wire            n20117;
wire            n20118;
wire            n20119;
wire            n20120;
wire            n20121;
wire            n20122;
wire            n20123;
wire            n20124;
wire            n20125;
wire            n20126;
wire            n20127;
wire            n20128;
wire            n20129;
wire            n20130;
wire            n20131;
wire            n20132;
wire            n20133;
wire            n20134;
wire            n20135;
wire            n20136;
wire            n20137;
wire            n20138;
wire            n20139;
wire            n20140;
wire            n20141;
wire            n20142;
wire            n20143;
wire            n20144;
wire            n20145;
wire            n20146;
wire            n20147;
wire            n20148;
wire            n20149;
wire            n20150;
wire            n20151;
wire            n20152;
wire            n20153;
wire            n20154;
wire            n20155;
wire            n20156;
wire            n20157;
wire            n20158;
wire            n20159;
wire            n20160;
wire            n20161;
wire            n20162;
wire            n20163;
wire            n20164;
wire            n20165;
wire            n20166;
wire            n20167;
wire            n20168;
wire            n20169;
wire            n20170;
wire            n20171;
wire            n20172;
wire            n20173;
wire            n20174;
wire            n20175;
wire            n20176;
wire            n20177;
wire            n20178;
wire            n20179;
wire            n20180;
wire            n20181;
wire            n20182;
wire            n20183;
wire            n20184;
wire            n20185;
wire            n20186;
wire            n20187;
wire            n20188;
wire            n20189;
wire            n20190;
wire            n20191;
wire            n20192;
wire            n20193;
wire            n20194;
wire            n20195;
wire            n20196;
wire            n20197;
wire            n20198;
wire            n20199;
wire            n20200;
wire            n20201;
wire            n20202;
wire            n20203;
wire            n20204;
wire            n20205;
wire            n20206;
wire            n20207;
wire            n20208;
wire            n20209;
wire            n20210;
wire            n20211;
wire            n20212;
wire            n20213;
wire            n20214;
wire            n20215;
wire            n20216;
wire            n20217;
wire            n20218;
wire            n20219;
wire            n20220;
wire            n20221;
wire            n20222;
wire            n20223;
wire            n20224;
wire            n20225;
wire            n20226;
wire            n20227;
wire            n20228;
wire            n20229;
wire            n20230;
wire            n20231;
wire            n20232;
wire            n20233;
wire            n20234;
wire            n20235;
wire            n20236;
wire            n20237;
wire            n20238;
wire            n20239;
wire            n20240;
wire            n20241;
wire            n20242;
wire            n20243;
wire            n20244;
wire            n20245;
wire            n20246;
wire            n20247;
wire            n20248;
wire            n20249;
wire            n20250;
wire            n20251;
wire            n20252;
wire            n20253;
wire            n20254;
wire            n20255;
wire            n20256;
wire            n20257;
wire            n20258;
wire            n20259;
wire            n20260;
wire            n20261;
wire            n20262;
wire            n20263;
wire            n20264;
wire            n20265;
wire            n20266;
wire            n20267;
wire            n20268;
wire            n20269;
wire            n20270;
wire            n20271;
wire            n20272;
wire            n20273;
wire            n20274;
wire            n20275;
wire            n20276;
wire            n20277;
wire            n20278;
wire            n20279;
wire            n20280;
wire            n20281;
wire            n20282;
wire            n20283;
wire            n20284;
wire            n20285;
wire            n20286;
wire            n20287;
wire            n20288;
wire            n20289;
wire            n20290;
wire            n20291;
wire            n20292;
wire            n20293;
wire            n20294;
wire            n20295;
wire            n20296;
wire            n20297;
wire            n20298;
wire            n20299;
wire            n20300;
wire            n20301;
wire            n20302;
wire            n20303;
wire            n20304;
wire            n20305;
wire            n20306;
wire            n20307;
wire            n20308;
wire            n20309;
wire            n20310;
wire            n20311;
wire            n20312;
wire            n20313;
wire            n20314;
wire            n20315;
wire            n20316;
wire            n20317;
wire            n20318;
wire            n20319;
wire            n20320;
wire            n20321;
wire            n20322;
wire            n20323;
wire            n20324;
wire            n20325;
wire            n20326;
wire            n20327;
wire            n20328;
wire            n20329;
wire            n20330;
wire            n20331;
wire            n20332;
wire            n20333;
wire            n20334;
wire            n20335;
wire            n20336;
wire            n20337;
wire            n20338;
wire            n20339;
wire            n20340;
wire            n20341;
wire            n20342;
wire            n20343;
wire            n20344;
wire            n20345;
wire            n20346;
wire            n20347;
wire            n20348;
wire            n20349;
wire            n20350;
wire            n20351;
wire            n20352;
wire            n20353;
wire            n20354;
wire            n20355;
wire            n20356;
wire            n20357;
wire            n20358;
wire            n20359;
wire            n20360;
wire            n20361;
wire            n20362;
wire            n20363;
wire            n20364;
wire            n20365;
wire            n20366;
wire            n20367;
wire            n20368;
wire            n20369;
wire            n20370;
wire            n20371;
wire            n20372;
wire            n20373;
wire            n20374;
wire            n20375;
wire            n20376;
wire            n20377;
wire            n20378;
wire            n20379;
wire            n20380;
wire            n20381;
wire            n20382;
wire            n20383;
wire            n20384;
wire            n20385;
wire            n20386;
wire            n20387;
wire            n20388;
wire            n20389;
wire            n20390;
wire            n20391;
wire            n20392;
wire            n20393;
wire            n20394;
wire            n20395;
wire            n20396;
wire            n20397;
wire            n20398;
wire            n20399;
wire            n20400;
wire            n20401;
wire            n20402;
wire            n20403;
wire            n20404;
wire            n20405;
wire            n20406;
wire            n20407;
wire            n20408;
wire            n20409;
wire            n20410;
wire            n20411;
wire            n20412;
wire            n20413;
wire            n20414;
wire            n20415;
wire            n20416;
wire            n20417;
wire            n20418;
wire            n20419;
wire            n20420;
wire            n20421;
wire            n20422;
wire            n20423;
wire            n20424;
wire            n20425;
wire            n20426;
wire            n20427;
wire            n20428;
wire            n20429;
wire            n20430;
wire            n20431;
wire            n20432;
wire            n20433;
wire            n20434;
wire            n20435;
wire            n20436;
wire            n20437;
wire            n20438;
wire            n20439;
wire            n20440;
wire            n20441;
wire            n20442;
wire            n20443;
wire            n20444;
wire            n20445;
wire            n20446;
wire            n20447;
wire            n20448;
wire            n20449;
wire            n20450;
wire            n20451;
wire            n20452;
wire            n20453;
wire            n20454;
wire            n20455;
wire            n20456;
wire            n20457;
wire            n20458;
wire            n20459;
wire            n20460;
wire            n20461;
wire            n20462;
wire            n20463;
wire            n20464;
wire            n20465;
wire            n20466;
wire            n20467;
wire            n20468;
wire            n20469;
wire            n20470;
wire            n20471;
wire            n20472;
wire            n20473;
wire            n20474;
wire            n20475;
wire            n20476;
wire            n20477;
wire            n20478;
wire            n20479;
wire            n20480;
wire            n20481;
wire            n20482;
wire            n20483;
wire            n20484;
wire            n20485;
wire            n20486;
wire            n20487;
wire            n20488;
wire            n20489;
wire            n20490;
wire            n20491;
wire            n20492;
wire            n20493;
wire            n20494;
wire            n20495;
wire            n20496;
wire            n20497;
wire            n20498;
wire            n20499;
wire            n20500;
wire            n20501;
wire            n20502;
wire            n20503;
wire            n20504;
wire            n20505;
wire            n20506;
wire            n20507;
wire            n20508;
wire            n20509;
wire            n20510;
wire            n20511;
wire            n20512;
wire            n20513;
wire            n20514;
wire            n20515;
wire            n20516;
wire            n20517;
wire            n20518;
wire            n20519;
wire            n20520;
wire            n20521;
wire            n20522;
wire            n20523;
wire            n20524;
wire            n20525;
wire            n20526;
wire            n20527;
wire            n20528;
wire            n20529;
wire            n20530;
wire            n20531;
wire            n20532;
wire            n20533;
wire            n20534;
wire            n20535;
wire            n20536;
wire            n20537;
wire            n20538;
wire            n20539;
wire            n20540;
wire            n20541;
wire            n20542;
wire            n20543;
wire            n20544;
wire            n20545;
wire            n20546;
wire            n20547;
wire            n20548;
wire     [31:0] n20549;
wire     [31:0] n20550;
wire     [31:0] n20551;
wire     [31:0] n20552;
wire     [31:0] n20553;
wire     [31:0] n20554;
wire     [31:0] n20555;
wire     [31:0] n20556;
wire     [31:0] n20557;
wire     [31:0] n20558;
wire     [31:0] n20559;
wire     [31:0] n20560;
wire     [31:0] n20561;
wire     [31:0] n20562;
wire     [31:0] n20563;
wire     [31:0] n20564;
wire     [31:0] n20565;
wire     [31:0] n20566;
wire     [31:0] n20567;
wire     [31:0] n20568;
wire     [31:0] n20569;
wire     [31:0] n20570;
wire     [31:0] n20571;
wire     [31:0] n20572;
wire     [31:0] n20573;
wire     [31:0] n20574;
wire     [31:0] n20575;
wire     [31:0] n20576;
wire     [31:0] n20577;
wire     [31:0] n20578;
wire     [31:0] n20579;
wire     [31:0] n20580;
wire     [31:0] n20581;
wire     [31:0] n20582;
wire     [31:0] n20583;
wire     [31:0] n20584;
wire     [31:0] n20585;
wire     [31:0] n20586;
wire     [31:0] n20587;
wire     [31:0] n20588;
wire     [31:0] n20589;
wire     [31:0] n20590;
wire     [31:0] n20591;
wire     [31:0] n20592;
wire     [31:0] n20593;
wire     [31:0] n20594;
wire     [31:0] n20595;
wire     [31:0] n20596;
wire     [31:0] n20597;
wire     [31:0] n20598;
wire     [31:0] n20599;
wire     [31:0] n20600;
wire     [31:0] n20601;
wire     [31:0] n20602;
wire     [31:0] n20603;
wire     [31:0] n20604;
wire     [31:0] n20605;
wire     [31:0] n20606;
wire     [31:0] n20607;
wire     [31:0] n20608;
wire     [31:0] n20609;
wire     [31:0] n20610;
wire     [31:0] n20611;
wire     [31:0] n20612;
wire     [31:0] n20613;
wire     [31:0] n20614;
wire     [31:0] n20615;
wire     [31:0] n20616;
wire     [31:0] n20617;
wire     [31:0] n20618;
wire     [31:0] n20619;
wire     [31:0] n20620;
wire     [31:0] n20621;
wire     [31:0] n20622;
wire     [31:0] n20623;
wire     [31:0] n20624;
wire     [31:0] n20625;
wire     [31:0] n20626;
wire     [31:0] n20627;
wire     [31:0] n20628;
wire     [31:0] n20629;
wire     [31:0] n20630;
wire     [31:0] n20631;
wire     [31:0] n20632;
wire     [31:0] n20633;
wire     [31:0] n20634;
wire     [31:0] n20635;
wire     [31:0] n20636;
wire     [31:0] n20637;
wire     [31:0] n20638;
wire     [31:0] n20639;
wire     [31:0] n20640;
wire     [31:0] n20641;
wire     [31:0] n20642;
wire     [31:0] n20643;
wire     [31:0] n20644;
wire     [31:0] n20645;
wire     [31:0] n20646;
wire     [31:0] n20647;
wire     [31:0] n20648;
wire     [31:0] n20649;
wire     [31:0] n20650;
wire     [31:0] n20651;
wire     [31:0] n20652;
wire     [31:0] n20653;
wire     [31:0] n20654;
wire     [31:0] n20655;
wire     [31:0] n20656;
wire     [31:0] n20657;
wire     [31:0] n20658;
wire     [31:0] n20659;
wire     [31:0] n20660;
wire     [31:0] n20661;
wire     [31:0] n20662;
wire     [31:0] n20663;
wire     [31:0] n20664;
wire     [31:0] n20665;
wire     [31:0] n20666;
wire     [31:0] n20667;
wire     [31:0] n20668;
wire     [31:0] n20669;
wire     [31:0] n20670;
wire     [31:0] n20671;
wire     [31:0] n20672;
wire     [31:0] n20673;
wire     [31:0] n20674;
wire     [31:0] n20675;
wire     [31:0] n20676;
wire     [31:0] n20677;
wire     [31:0] n20678;
wire     [31:0] n20679;
wire     [31:0] n20680;
wire     [31:0] n20681;
wire     [31:0] n20682;
wire     [31:0] n20683;
wire     [31:0] n20684;
wire     [31:0] n20685;
wire     [31:0] n20686;
wire     [31:0] n20687;
wire     [31:0] n20688;
wire     [31:0] n20689;
wire     [31:0] n20690;
wire     [31:0] n20691;
wire     [31:0] n20692;
wire     [31:0] n20693;
wire     [31:0] n20694;
wire     [31:0] n20695;
wire     [31:0] n20696;
wire     [31:0] n20697;
wire     [31:0] n20698;
wire     [31:0] n20699;
wire     [31:0] n20700;
wire     [31:0] n20701;
wire     [31:0] n20702;
wire     [31:0] n20703;
wire     [31:0] n20704;
wire     [31:0] n20705;
wire     [31:0] n20706;
wire     [31:0] n20707;
wire     [31:0] n20708;
wire     [31:0] n20709;
wire     [31:0] n20710;
wire     [31:0] n20711;
wire     [31:0] n20712;
wire     [31:0] n20713;
wire     [31:0] n20714;
wire     [31:0] n20715;
wire     [31:0] n20716;
wire     [31:0] n20717;
wire     [31:0] n20718;
wire     [31:0] n20719;
wire     [31:0] n20720;
wire     [31:0] n20721;
wire     [31:0] n20722;
wire     [31:0] n20723;
wire     [31:0] n20724;
wire     [31:0] n20725;
wire     [31:0] n20726;
wire     [31:0] n20727;
wire     [31:0] n20728;
wire     [31:0] n20729;
wire     [31:0] n20730;
wire     [31:0] n20731;
wire     [31:0] n20732;
wire     [31:0] n20733;
wire     [31:0] n20734;
wire     [31:0] n20735;
wire     [31:0] n20736;
wire     [31:0] n20737;
wire     [31:0] n20738;
wire     [31:0] n20739;
wire     [31:0] n20740;
wire     [31:0] n20741;
wire     [31:0] n20742;
wire     [31:0] n20743;
wire     [31:0] n20744;
wire     [31:0] n20745;
wire     [31:0] n20746;
wire     [31:0] n20747;
wire     [31:0] n20748;
wire     [31:0] n20749;
wire     [31:0] n20750;
wire     [31:0] n20751;
wire     [31:0] n20752;
wire     [31:0] n20753;
wire     [31:0] n20754;
wire     [31:0] n20755;
wire     [31:0] n20756;
wire     [31:0] n20757;
wire     [31:0] n20758;
wire     [31:0] n20759;
wire     [31:0] n20760;
wire     [31:0] n20761;
wire     [31:0] n20762;
wire     [31:0] n20763;
wire     [31:0] n20764;
wire     [31:0] n20765;
wire     [31:0] n20766;
wire     [31:0] n20767;
wire     [31:0] n20768;
wire     [31:0] n20769;
wire     [31:0] n20770;
wire     [31:0] n20771;
wire     [31:0] n20772;
wire     [31:0] n20773;
wire     [31:0] n20774;
wire     [31:0] n20775;
wire     [31:0] n20776;
wire     [31:0] n20777;
wire     [31:0] n20778;
wire     [31:0] n20779;
wire     [31:0] n20780;
wire     [31:0] n20781;
wire     [31:0] n20782;
wire     [31:0] n20783;
wire     [31:0] n20784;
wire     [31:0] n20785;
wire     [31:0] n20786;
wire     [31:0] n20787;
wire     [31:0] n20788;
wire     [31:0] n20789;
wire     [31:0] n20790;
wire     [31:0] n20791;
wire     [31:0] n20792;
wire     [31:0] n20793;
wire     [31:0] n20794;
wire     [31:0] n20795;
wire     [31:0] n20796;
wire     [31:0] n20797;
wire     [31:0] n20798;
wire     [31:0] n20799;
wire     [31:0] n20800;
wire     [31:0] n20801;
wire     [31:0] n20802;
wire     [31:0] n20803;
wire     [31:0] n20804;
wire     [31:0] n20805;
wire     [31:0] n20806;
wire     [31:0] n20807;
wire     [31:0] n20808;
wire     [31:0] n20809;
wire     [31:0] n20810;
wire     [31:0] n20811;
wire     [31:0] n20812;
wire     [31:0] n20813;
wire     [31:0] n20814;
wire     [31:0] n20815;
wire     [31:0] n20816;
wire     [31:0] n20817;
wire     [31:0] n20818;
wire     [31:0] n20819;
wire     [31:0] n20820;
wire     [31:0] n20821;
wire     [31:0] n20822;
wire     [31:0] n20823;
wire     [31:0] n20824;
wire     [31:0] n20825;
wire     [31:0] n20826;
wire     [31:0] n20827;
wire     [31:0] n20828;
wire     [31:0] n20829;
wire     [31:0] n20830;
wire     [31:0] n20831;
wire     [31:0] n20832;
wire     [31:0] n20833;
wire     [31:0] n20834;
wire     [31:0] n20835;
wire     [31:0] n20836;
wire     [31:0] n20837;
wire     [31:0] n20838;
wire     [31:0] n20839;
wire     [31:0] n20840;
wire     [31:0] n20841;
wire     [31:0] n20842;
wire     [31:0] n20843;
wire     [31:0] n20844;
wire     [31:0] n20845;
wire     [31:0] n20846;
wire     [31:0] n20847;
wire     [31:0] n20848;
wire     [31:0] n20849;
wire     [31:0] n20850;
wire     [31:0] n20851;
wire     [31:0] n20852;
wire     [31:0] n20853;
wire     [31:0] n20854;
wire     [31:0] n20855;
wire     [31:0] n20856;
wire     [31:0] n20857;
wire     [31:0] n20858;
wire     [31:0] n20859;
wire     [31:0] n20860;
wire     [31:0] n20861;
wire     [31:0] n20862;
wire     [31:0] n20863;
wire     [31:0] n20864;
wire     [31:0] n20865;
wire     [31:0] n20866;
wire     [31:0] n20867;
wire     [31:0] n20868;
wire     [31:0] n20869;
wire     [31:0] n20870;
wire     [31:0] n20871;
wire     [31:0] n20872;
wire     [31:0] n20873;
wire     [31:0] n20874;
wire     [31:0] n20875;
wire     [31:0] n20876;
wire     [31:0] n20877;
wire     [31:0] n20878;
wire     [31:0] n20879;
wire     [31:0] n20880;
wire     [31:0] n20881;
wire     [31:0] n20882;
wire     [31:0] n20883;
wire     [31:0] n20884;
wire     [31:0] n20885;
wire     [31:0] n20886;
wire     [31:0] n20887;
wire     [31:0] n20888;
wire     [31:0] n20889;
wire     [31:0] n20890;
wire     [31:0] n20891;
wire     [31:0] n20892;
wire     [31:0] n20893;
wire     [31:0] n20894;
wire     [31:0] n20895;
wire     [31:0] n20896;
wire     [31:0] n20897;
wire     [31:0] n20898;
wire     [31:0] n20899;
wire     [31:0] n20900;
wire     [31:0] n20901;
wire     [31:0] n20902;
wire     [31:0] n20903;
wire     [31:0] n20904;
wire     [31:0] n20905;
wire     [31:0] n20906;
wire     [31:0] n20907;
wire     [31:0] n20908;
wire     [31:0] n20909;
wire     [31:0] n20910;
wire     [31:0] n20911;
wire     [31:0] n20912;
wire     [31:0] n20913;
wire     [31:0] n20914;
wire     [31:0] n20915;
wire     [31:0] n20916;
wire     [31:0] n20917;
wire     [31:0] n20918;
wire     [31:0] n20919;
wire     [31:0] n20920;
wire     [31:0] n20921;
wire     [31:0] n20922;
wire     [31:0] n20923;
wire     [31:0] n20924;
wire     [31:0] n20925;
wire     [31:0] n20926;
wire     [31:0] n20927;
wire     [31:0] n20928;
wire     [31:0] n20929;
wire     [31:0] n20930;
wire     [31:0] n20931;
wire     [31:0] n20932;
wire     [31:0] n20933;
wire     [31:0] n20934;
wire     [31:0] n20935;
wire     [31:0] n20936;
wire     [31:0] n20937;
wire     [31:0] n20938;
wire     [31:0] n20939;
wire     [31:0] n20940;
wire     [31:0] n20941;
wire     [31:0] n20942;
wire     [31:0] n20943;
wire     [31:0] n20944;
wire     [31:0] n20945;
wire     [31:0] n20946;
wire     [31:0] n20947;
wire     [31:0] n20948;
wire     [31:0] n20949;
wire     [31:0] n20950;
wire     [31:0] n20951;
wire     [31:0] n20952;
wire     [31:0] n20953;
wire     [31:0] n20954;
wire     [31:0] n20955;
wire     [31:0] n20956;
wire     [31:0] n20957;
wire     [31:0] n20958;
wire     [31:0] n20959;
wire     [31:0] n20960;
wire     [31:0] n20961;
wire     [31:0] n20962;
wire     [31:0] n20963;
wire     [31:0] n20964;
wire     [31:0] n20965;
wire     [31:0] n20966;
wire     [31:0] n20967;
wire     [31:0] n20968;
wire     [31:0] n20969;
wire     [31:0] n20970;
wire     [31:0] n20971;
wire     [31:0] n20972;
wire     [31:0] n20973;
wire     [31:0] n20974;
wire     [31:0] n20975;
wire     [31:0] n20976;
wire     [31:0] n20977;
wire     [31:0] n20978;
wire     [31:0] n20979;
wire     [31:0] n20980;
wire     [31:0] n20981;
wire     [31:0] n20982;
wire     [31:0] n20983;
wire     [31:0] n20984;
wire     [31:0] n20985;
wire     [31:0] n20986;
wire     [31:0] n20987;
wire     [31:0] n20988;
wire     [31:0] n20989;
wire     [31:0] n20990;
wire     [31:0] n20991;
wire     [31:0] n20992;
wire     [31:0] n20993;
wire     [31:0] n20994;
wire     [31:0] n20995;
wire     [31:0] n20996;
wire     [31:0] n20997;
wire     [31:0] n20998;
wire     [31:0] n20999;
wire     [31:0] n21000;
wire     [31:0] n21001;
wire     [31:0] n21002;
wire     [31:0] n21003;
wire     [31:0] n21004;
wire     [31:0] n21005;
wire     [31:0] n21006;
wire     [31:0] n21007;
wire     [31:0] n21008;
wire     [31:0] n21009;
wire     [31:0] n21010;
wire     [31:0] n21011;
wire     [31:0] n21012;
wire     [31:0] n21013;
wire     [31:0] n21014;
wire     [31:0] n21015;
wire     [31:0] n21016;
wire     [31:0] n21017;
wire     [31:0] n21018;
wire     [31:0] n21019;
wire     [31:0] n21020;
wire     [31:0] n21021;
wire     [31:0] n21022;
wire     [31:0] n21023;
wire     [31:0] n21024;
wire     [31:0] n21025;
wire     [31:0] n21026;
wire     [31:0] n21027;
wire     [31:0] n21028;
wire     [31:0] n21029;
wire     [31:0] n21030;
wire     [31:0] n21031;
wire     [31:0] n21032;
wire     [31:0] n21033;
wire     [31:0] n21034;
wire     [31:0] n21035;
wire     [31:0] n21036;
wire     [31:0] n21037;
wire     [31:0] n21038;
wire     [31:0] n21039;
wire     [31:0] n21040;
wire     [31:0] n21041;
wire     [31:0] n21042;
wire     [31:0] n21043;
wire     [31:0] n21044;
wire     [31:0] n21045;
wire     [31:0] n21046;
wire     [31:0] n21047;
wire     [31:0] n21048;
wire     [31:0] n21049;
wire     [31:0] n21050;
wire     [31:0] n21051;
wire     [31:0] n21052;
wire     [31:0] n21053;
wire     [31:0] n21054;
wire     [31:0] n21055;
wire     [31:0] n21056;
wire     [31:0] n21057;
wire     [31:0] n21058;
wire     [31:0] n21059;
wire     [31:0] n21060;
wire     [31:0] n21061;
wire     [31:0] n21062;
wire     [31:0] n21063;
wire     [31:0] n21064;
wire     [31:0] n21065;
wire     [31:0] n21066;
wire     [31:0] n21067;
wire     [31:0] n21068;
wire     [31:0] n21069;
wire     [31:0] n21070;
wire            n21071;
wire            n21072;
wire            n21073;
wire            n21074;
wire            n21075;
wire            n21076;
wire            n21077;
wire            n21078;
wire            n21079;
wire            n21080;
wire            n21081;
wire            n21082;
wire            n21083;
wire            n21084;
wire            n21085;
wire            n21086;
wire            n21087;
wire            n21088;
wire            n21089;
wire            n21090;
wire            n21091;
wire            n21092;
wire            n21093;
wire            n21094;
wire            n21095;
wire            n21096;
wire            n21097;
wire            n21098;
wire            n21099;
wire            n21100;
wire            n21101;
wire            n21102;
wire            n21103;
wire            n21104;
wire            n21105;
wire            n21106;
wire            n21107;
wire            n21108;
wire            n21109;
wire            n21110;
wire            n21111;
wire            n21112;
wire            n21113;
wire            n21114;
wire            n21115;
wire            n21116;
wire            n21117;
wire            n21118;
wire            n21119;
wire            n21120;
wire            n21121;
wire            n21122;
wire            n21123;
wire            n21124;
wire            n21125;
wire            n21126;
wire            n21127;
wire            n21128;
wire            n21129;
wire            n21130;
wire            n21131;
wire            n21132;
wire            n21133;
wire            n21134;
wire            n21135;
wire            n21136;
wire            n21137;
wire            n21138;
wire            n21139;
wire            n21140;
wire            n21141;
wire            n21142;
wire            n21143;
wire            n21144;
wire            n21145;
wire            n21146;
wire            n21147;
wire            n21148;
wire            n21149;
wire            n21150;
wire            n21151;
wire            n21152;
wire            n21153;
wire            n21154;
wire            n21155;
wire            n21156;
wire            n21157;
wire            n21158;
wire            n21159;
wire            n21160;
wire            n21161;
wire            n21162;
wire            n21163;
wire            n21164;
wire            n21165;
wire            n21166;
wire            n21167;
wire            n21168;
wire            n21169;
wire            n21170;
wire            n21171;
wire            n21172;
wire            n21173;
wire            n21174;
wire            n21175;
wire            n21176;
wire            n21177;
wire            n21178;
wire            n21179;
wire            n21180;
wire            n21181;
wire            n21182;
wire            n21183;
wire            n21184;
wire            n21185;
wire            n21186;
wire            n21187;
wire            n21188;
wire            n21189;
wire            n21190;
wire            n21191;
wire            n21192;
wire            n21193;
wire            n21194;
wire            n21195;
wire            n21196;
wire            n21197;
wire            n21198;
wire            n21199;
wire            n21200;
wire            n21201;
wire            n21202;
wire            n21203;
wire            n21204;
wire            n21205;
wire            n21206;
wire            n21207;
wire            n21208;
wire            n21209;
wire            n21210;
wire            n21211;
wire            n21212;
wire            n21213;
wire            n21214;
wire            n21215;
wire            n21216;
wire            n21217;
wire            n21218;
wire            n21219;
wire            n21220;
wire            n21221;
wire            n21222;
wire            n21223;
wire            n21224;
wire            n21225;
wire            n21226;
wire            n21227;
wire            n21228;
wire            n21229;
wire            n21230;
wire            n21231;
wire            n21232;
wire            n21233;
wire            n21234;
wire            n21235;
wire            n21236;
wire            n21237;
wire            n21238;
wire            n21239;
wire            n21240;
wire            n21241;
wire            n21242;
wire            n21243;
wire            n21244;
wire            n21245;
wire            n21246;
wire            n21247;
wire            n21248;
wire            n21249;
wire            n21250;
wire            n21251;
wire            n21252;
wire            n21253;
wire            n21254;
wire            n21255;
wire            n21256;
wire            n21257;
wire            n21258;
wire            n21259;
wire            n21260;
wire            n21261;
wire            n21262;
wire            n21263;
wire            n21264;
wire            n21265;
wire            n21266;
wire            n21267;
wire            n21268;
wire            n21269;
wire            n21270;
wire            n21271;
wire            n21272;
wire            n21273;
wire            n21274;
wire            n21275;
wire            n21276;
wire            n21277;
wire            n21278;
wire            n21279;
wire            n21280;
wire            n21281;
wire            n21282;
wire            n21283;
wire            n21284;
wire            n21285;
wire            n21286;
wire            n21287;
wire            n21288;
wire            n21289;
wire            n21290;
wire            n21291;
wire            n21292;
wire            n21293;
wire            n21294;
wire            n21295;
wire            n21296;
wire            n21297;
wire            n21298;
wire            n21299;
wire            n21300;
wire            n21301;
wire            n21302;
wire            n21303;
wire            n21304;
wire            n21305;
wire            n21306;
wire            n21307;
wire            n21308;
wire            n21309;
wire            n21310;
wire            n21311;
wire            n21312;
wire            n21313;
wire            n21314;
wire            n21315;
wire            n21316;
wire            n21317;
wire            n21318;
wire            n21319;
wire            n21320;
wire            n21321;
wire            n21322;
wire            n21323;
wire            n21324;
wire            n21325;
wire            n21326;
wire            n21327;
wire            n21328;
wire            n21329;
wire            n21330;
wire            n21331;
wire            n21332;
wire            n21333;
wire            n21334;
wire            n21335;
wire            n21336;
wire            n21337;
wire            n21338;
wire            n21339;
wire            n21340;
wire            n21341;
wire            n21342;
wire            n21343;
wire            n21344;
wire            n21345;
wire            n21346;
wire            n21347;
wire            n21348;
wire            n21349;
wire            n21350;
wire            n21351;
wire            n21352;
wire            n21353;
wire            n21354;
wire            n21355;
wire            n21356;
wire            n21357;
wire            n21358;
wire            n21359;
wire            n21360;
wire            n21361;
wire            n21362;
wire            n21363;
wire            n21364;
wire            n21365;
wire            n21366;
wire            n21367;
wire            n21368;
wire            n21369;
wire            n21370;
wire            n21371;
wire            n21372;
wire            n21373;
wire            n21374;
wire            n21375;
wire            n21376;
wire            n21377;
wire            n21378;
wire            n21379;
wire            n21380;
wire            n21381;
wire            n21382;
wire            n21383;
wire            n21384;
wire            n21385;
wire            n21386;
wire            n21387;
wire            n21388;
wire            n21389;
wire            n21390;
wire            n21391;
wire            n21392;
wire            n21393;
wire            n21394;
wire            n21395;
wire            n21396;
wire            n21397;
wire            n21398;
wire            n21399;
wire            n21400;
wire            n21401;
wire            n21402;
wire            n21403;
wire            n21404;
wire            n21405;
wire            n21406;
wire            n21407;
wire            n21408;
wire            n21409;
wire            n21410;
wire            n21411;
wire            n21412;
wire            n21413;
wire            n21414;
wire            n21415;
wire            n21416;
wire            n21417;
wire            n21418;
wire            n21419;
wire            n21420;
wire            n21421;
wire            n21422;
wire            n21423;
wire            n21424;
wire            n21425;
wire            n21426;
wire            n21427;
wire            n21428;
wire            n21429;
wire            n21430;
wire            n21431;
wire            n21432;
wire            n21433;
wire            n21434;
wire            n21435;
wire            n21436;
wire            n21437;
wire            n21438;
wire            n21439;
wire            n21440;
wire            n21441;
wire            n21442;
wire            n21443;
wire            n21444;
wire            n21445;
wire            n21446;
wire            n21447;
wire            n21448;
wire            n21449;
wire            n21450;
wire            n21451;
wire            n21452;
wire            n21453;
wire            n21454;
wire            n21455;
wire            n21456;
wire            n21457;
wire            n21458;
wire            n21459;
wire            n21460;
wire            n21461;
wire            n21462;
wire            n21463;
wire            n21464;
wire            n21465;
wire            n21466;
wire            n21467;
wire            n21468;
wire            n21469;
wire            n21470;
wire            n21471;
wire            n21472;
wire            n21473;
wire            n21474;
wire            n21475;
wire            n21476;
wire            n21477;
wire            n21478;
wire            n21479;
wire            n21480;
wire            n21481;
wire            n21482;
wire            n21483;
wire            n21484;
wire            n21485;
wire            n21486;
wire            n21487;
wire            n21488;
wire            n21489;
wire            n21490;
wire            n21491;
wire            n21492;
wire            n21493;
wire            n21494;
wire            n21495;
wire            n21496;
wire            n21497;
wire            n21498;
wire            n21499;
wire            n21500;
wire            n21501;
wire            n21502;
wire            n21503;
wire            n21504;
wire            n21505;
wire            n21506;
wire            n21507;
wire            n21508;
wire            n21509;
wire            n21510;
wire            n21511;
wire            n21512;
wire            n21513;
wire            n21514;
wire            n21515;
wire            n21516;
wire            n21517;
wire            n21518;
wire            n21519;
wire            n21520;
wire            n21521;
wire            n21522;
wire            n21523;
wire            n21524;
wire            n21525;
wire            n21526;
wire            n21527;
wire            n21528;
wire            n21529;
wire            n21530;
wire            n21531;
wire            n21532;
wire            n21533;
wire            n21534;
wire            n21535;
wire            n21536;
wire            n21537;
wire            n21538;
wire            n21539;
wire            n21540;
wire            n21541;
wire            n21542;
wire            n21543;
wire            n21544;
wire            n21545;
wire            n21546;
wire            n21547;
wire            n21548;
wire            n21549;
wire            n21550;
wire            n21551;
wire            n21552;
wire            n21553;
wire            n21554;
wire            n21555;
wire            n21556;
wire            n21557;
wire            n21558;
wire            n21559;
wire            n21560;
wire            n21561;
wire            n21562;
wire            n21563;
wire            n21564;
wire            n21565;
wire            n21566;
wire            n21567;
wire            n21568;
wire            n21569;
wire            n21570;
wire            n21571;
wire            n21572;
wire            n21573;
wire            n21574;
wire            n21575;
wire            n21576;
wire            n21577;
wire            n21578;
wire            n21579;
wire            n21580;
wire            n21581;
wire            n21582;
wire     [31:0] n21583;
wire     [31:0] n21584;
wire     [31:0] n21585;
wire     [31:0] n21586;
wire     [31:0] n21587;
wire     [31:0] n21588;
wire     [31:0] n21589;
wire     [31:0] n21590;
wire     [31:0] n21591;
wire     [31:0] n21592;
wire     [31:0] n21593;
wire     [31:0] n21594;
wire     [31:0] n21595;
wire     [31:0] n21596;
wire     [31:0] n21597;
wire     [31:0] n21598;
wire     [31:0] n21599;
wire     [31:0] n21600;
wire     [31:0] n21601;
wire     [31:0] n21602;
wire     [31:0] n21603;
wire     [31:0] n21604;
wire     [31:0] n21605;
wire     [31:0] n21606;
wire     [31:0] n21607;
wire     [31:0] n21608;
wire     [31:0] n21609;
wire     [31:0] n21610;
wire     [31:0] n21611;
wire     [31:0] n21612;
wire     [31:0] n21613;
wire     [31:0] n21614;
wire     [31:0] n21615;
wire     [31:0] n21616;
wire     [31:0] n21617;
wire     [31:0] n21618;
wire     [31:0] n21619;
wire     [31:0] n21620;
wire     [31:0] n21621;
wire     [31:0] n21622;
wire     [31:0] n21623;
wire     [31:0] n21624;
wire     [31:0] n21625;
wire     [31:0] n21626;
wire     [31:0] n21627;
wire     [31:0] n21628;
wire     [31:0] n21629;
wire     [31:0] n21630;
wire     [31:0] n21631;
wire     [31:0] n21632;
wire     [31:0] n21633;
wire     [31:0] n21634;
wire     [31:0] n21635;
wire     [31:0] n21636;
wire     [31:0] n21637;
wire     [31:0] n21638;
wire     [31:0] n21639;
wire     [31:0] n21640;
wire     [31:0] n21641;
wire     [31:0] n21642;
wire     [31:0] n21643;
wire     [31:0] n21644;
wire     [31:0] n21645;
wire     [31:0] n21646;
wire     [31:0] n21647;
wire     [31:0] n21648;
wire     [31:0] n21649;
wire     [31:0] n21650;
wire     [31:0] n21651;
wire     [31:0] n21652;
wire     [31:0] n21653;
wire     [31:0] n21654;
wire     [31:0] n21655;
wire     [31:0] n21656;
wire     [31:0] n21657;
wire     [31:0] n21658;
wire     [31:0] n21659;
wire     [31:0] n21660;
wire     [31:0] n21661;
wire     [31:0] n21662;
wire     [31:0] n21663;
wire     [31:0] n21664;
wire     [31:0] n21665;
wire     [31:0] n21666;
wire     [31:0] n21667;
wire     [31:0] n21668;
wire     [31:0] n21669;
wire     [31:0] n21670;
wire     [31:0] n21671;
wire     [31:0] n21672;
wire     [31:0] n21673;
wire     [31:0] n21674;
wire     [31:0] n21675;
wire     [31:0] n21676;
wire     [31:0] n21677;
wire     [31:0] n21678;
wire     [31:0] n21679;
wire     [31:0] n21680;
wire     [31:0] n21681;
wire     [31:0] n21682;
wire     [31:0] n21683;
wire     [31:0] n21684;
wire     [31:0] n21685;
wire     [31:0] n21686;
wire     [31:0] n21687;
wire     [31:0] n21688;
wire     [31:0] n21689;
wire     [31:0] n21690;
wire     [31:0] n21691;
wire     [31:0] n21692;
wire     [31:0] n21693;
wire     [31:0] n21694;
wire     [31:0] n21695;
wire     [31:0] n21696;
wire     [31:0] n21697;
wire     [31:0] n21698;
wire     [31:0] n21699;
wire     [31:0] n21700;
wire     [31:0] n21701;
wire     [31:0] n21702;
wire     [31:0] n21703;
wire     [31:0] n21704;
wire     [31:0] n21705;
wire     [31:0] n21706;
wire     [31:0] n21707;
wire     [31:0] n21708;
wire     [31:0] n21709;
wire     [31:0] n21710;
wire     [31:0] n21711;
wire     [31:0] n21712;
wire     [31:0] n21713;
wire     [31:0] n21714;
wire     [31:0] n21715;
wire     [31:0] n21716;
wire     [31:0] n21717;
wire     [31:0] n21718;
wire     [31:0] n21719;
wire     [31:0] n21720;
wire     [31:0] n21721;
wire     [31:0] n21722;
wire     [31:0] n21723;
wire     [31:0] n21724;
wire     [31:0] n21725;
wire     [31:0] n21726;
wire     [31:0] n21727;
wire     [31:0] n21728;
wire     [31:0] n21729;
wire     [31:0] n21730;
wire     [31:0] n21731;
wire     [31:0] n21732;
wire     [31:0] n21733;
wire     [31:0] n21734;
wire     [31:0] n21735;
wire     [31:0] n21736;
wire     [31:0] n21737;
wire     [31:0] n21738;
wire     [31:0] n21739;
wire     [31:0] n21740;
wire     [31:0] n21741;
wire     [31:0] n21742;
wire     [31:0] n21743;
wire     [31:0] n21744;
wire     [31:0] n21745;
wire     [31:0] n21746;
wire     [31:0] n21747;
wire     [31:0] n21748;
wire     [31:0] n21749;
wire     [31:0] n21750;
wire     [31:0] n21751;
wire     [31:0] n21752;
wire     [31:0] n21753;
wire     [31:0] n21754;
wire     [31:0] n21755;
wire     [31:0] n21756;
wire     [31:0] n21757;
wire     [31:0] n21758;
wire     [31:0] n21759;
wire     [31:0] n21760;
wire     [31:0] n21761;
wire     [31:0] n21762;
wire     [31:0] n21763;
wire     [31:0] n21764;
wire     [31:0] n21765;
wire     [31:0] n21766;
wire     [31:0] n21767;
wire     [31:0] n21768;
wire     [31:0] n21769;
wire     [31:0] n21770;
wire     [31:0] n21771;
wire     [31:0] n21772;
wire     [31:0] n21773;
wire     [31:0] n21774;
wire     [31:0] n21775;
wire     [31:0] n21776;
wire     [31:0] n21777;
wire     [31:0] n21778;
wire     [31:0] n21779;
wire     [31:0] n21780;
wire     [31:0] n21781;
wire     [31:0] n21782;
wire     [31:0] n21783;
wire     [31:0] n21784;
wire     [31:0] n21785;
wire     [31:0] n21786;
wire     [31:0] n21787;
wire     [31:0] n21788;
wire     [31:0] n21789;
wire     [31:0] n21790;
wire     [31:0] n21791;
wire     [31:0] n21792;
wire     [31:0] n21793;
wire     [31:0] n21794;
wire     [31:0] n21795;
wire     [31:0] n21796;
wire     [31:0] n21797;
wire     [31:0] n21798;
wire     [31:0] n21799;
wire     [31:0] n21800;
wire     [31:0] n21801;
wire     [31:0] n21802;
wire     [31:0] n21803;
wire     [31:0] n21804;
wire     [31:0] n21805;
wire     [31:0] n21806;
wire     [31:0] n21807;
wire     [31:0] n21808;
wire     [31:0] n21809;
wire     [31:0] n21810;
wire     [31:0] n21811;
wire     [31:0] n21812;
wire     [31:0] n21813;
wire     [31:0] n21814;
wire     [31:0] n21815;
wire     [31:0] n21816;
wire     [31:0] n21817;
wire     [31:0] n21818;
wire     [31:0] n21819;
wire     [31:0] n21820;
wire     [31:0] n21821;
wire     [31:0] n21822;
wire     [31:0] n21823;
wire     [31:0] n21824;
wire     [31:0] n21825;
wire     [31:0] n21826;
wire     [31:0] n21827;
wire     [31:0] n21828;
wire     [31:0] n21829;
wire     [31:0] n21830;
wire     [31:0] n21831;
wire     [31:0] n21832;
wire     [31:0] n21833;
wire     [31:0] n21834;
wire     [31:0] n21835;
wire     [31:0] n21836;
wire     [31:0] n21837;
wire     [31:0] n21838;
wire     [31:0] n21839;
wire     [31:0] n21840;
wire     [31:0] n21841;
wire     [31:0] n21842;
wire     [31:0] n21843;
wire     [31:0] n21844;
wire     [31:0] n21845;
wire     [31:0] n21846;
wire     [31:0] n21847;
wire     [31:0] n21848;
wire     [31:0] n21849;
wire     [31:0] n21850;
wire     [31:0] n21851;
wire     [31:0] n21852;
wire     [31:0] n21853;
wire     [31:0] n21854;
wire     [31:0] n21855;
wire     [31:0] n21856;
wire     [31:0] n21857;
wire     [31:0] n21858;
wire     [31:0] n21859;
wire     [31:0] n21860;
wire     [31:0] n21861;
wire     [31:0] n21862;
wire     [31:0] n21863;
wire     [31:0] n21864;
wire     [31:0] n21865;
wire     [31:0] n21866;
wire     [31:0] n21867;
wire     [31:0] n21868;
wire     [31:0] n21869;
wire     [31:0] n21870;
wire     [31:0] n21871;
wire     [31:0] n21872;
wire     [31:0] n21873;
wire     [31:0] n21874;
wire     [31:0] n21875;
wire     [31:0] n21876;
wire     [31:0] n21877;
wire     [31:0] n21878;
wire     [31:0] n21879;
wire     [31:0] n21880;
wire     [31:0] n21881;
wire     [31:0] n21882;
wire     [31:0] n21883;
wire     [31:0] n21884;
wire     [31:0] n21885;
wire     [31:0] n21886;
wire     [31:0] n21887;
wire     [31:0] n21888;
wire     [31:0] n21889;
wire     [31:0] n21890;
wire     [31:0] n21891;
wire     [31:0] n21892;
wire     [31:0] n21893;
wire     [31:0] n21894;
wire     [31:0] n21895;
wire     [31:0] n21896;
wire     [31:0] n21897;
wire     [31:0] n21898;
wire     [31:0] n21899;
wire     [31:0] n21900;
wire     [31:0] n21901;
wire     [31:0] n21902;
wire     [31:0] n21903;
wire     [31:0] n21904;
wire     [31:0] n21905;
wire     [31:0] n21906;
wire     [31:0] n21907;
wire     [31:0] n21908;
wire     [31:0] n21909;
wire     [31:0] n21910;
wire     [31:0] n21911;
wire     [31:0] n21912;
wire     [31:0] n21913;
wire     [31:0] n21914;
wire     [31:0] n21915;
wire     [31:0] n21916;
wire     [31:0] n21917;
wire     [31:0] n21918;
wire     [31:0] n21919;
wire     [31:0] n21920;
wire     [31:0] n21921;
wire     [31:0] n21922;
wire     [31:0] n21923;
wire     [31:0] n21924;
wire     [31:0] n21925;
wire     [31:0] n21926;
wire     [31:0] n21927;
wire     [31:0] n21928;
wire     [31:0] n21929;
wire     [31:0] n21930;
wire     [31:0] n21931;
wire     [31:0] n21932;
wire     [31:0] n21933;
wire     [31:0] n21934;
wire     [31:0] n21935;
wire     [31:0] n21936;
wire     [31:0] n21937;
wire     [31:0] n21938;
wire     [31:0] n21939;
wire     [31:0] n21940;
wire     [31:0] n21941;
wire     [31:0] n21942;
wire     [31:0] n21943;
wire     [31:0] n21944;
wire     [31:0] n21945;
wire     [31:0] n21946;
wire     [31:0] n21947;
wire     [31:0] n21948;
wire     [31:0] n21949;
wire     [31:0] n21950;
wire     [31:0] n21951;
wire     [31:0] n21952;
wire     [31:0] n21953;
wire     [31:0] n21954;
wire     [31:0] n21955;
wire     [31:0] n21956;
wire     [31:0] n21957;
wire     [31:0] n21958;
wire     [31:0] n21959;
wire     [31:0] n21960;
wire     [31:0] n21961;
wire     [31:0] n21962;
wire     [31:0] n21963;
wire     [31:0] n21964;
wire     [31:0] n21965;
wire     [31:0] n21966;
wire     [31:0] n21967;
wire     [31:0] n21968;
wire     [31:0] n21969;
wire     [31:0] n21970;
wire     [31:0] n21971;
wire     [31:0] n21972;
wire     [31:0] n21973;
wire     [31:0] n21974;
wire     [31:0] n21975;
wire     [31:0] n21976;
wire     [31:0] n21977;
wire     [31:0] n21978;
wire     [31:0] n21979;
wire     [31:0] n21980;
wire     [31:0] n21981;
wire     [31:0] n21982;
wire     [31:0] n21983;
wire     [31:0] n21984;
wire     [31:0] n21985;
wire     [31:0] n21986;
wire     [31:0] n21987;
wire     [31:0] n21988;
wire     [31:0] n21989;
wire     [31:0] n21990;
wire     [31:0] n21991;
wire     [31:0] n21992;
wire     [31:0] n21993;
wire     [31:0] n21994;
wire     [31:0] n21995;
wire     [31:0] n21996;
wire     [31:0] n21997;
wire     [31:0] n21998;
wire     [31:0] n21999;
wire     [31:0] n22000;
wire     [31:0] n22001;
wire     [31:0] n22002;
wire     [31:0] n22003;
wire     [31:0] n22004;
wire     [31:0] n22005;
wire     [31:0] n22006;
wire     [31:0] n22007;
wire     [31:0] n22008;
wire     [31:0] n22009;
wire     [31:0] n22010;
wire     [31:0] n22011;
wire     [31:0] n22012;
wire     [31:0] n22013;
wire     [31:0] n22014;
wire     [31:0] n22015;
wire     [31:0] n22016;
wire     [31:0] n22017;
wire     [31:0] n22018;
wire     [31:0] n22019;
wire     [31:0] n22020;
wire     [31:0] n22021;
wire     [31:0] n22022;
wire     [31:0] n22023;
wire     [31:0] n22024;
wire     [31:0] n22025;
wire     [31:0] n22026;
wire     [31:0] n22027;
wire     [31:0] n22028;
wire     [31:0] n22029;
wire     [31:0] n22030;
wire     [31:0] n22031;
wire     [31:0] n22032;
wire     [31:0] n22033;
wire     [31:0] n22034;
wire     [31:0] n22035;
wire     [31:0] n22036;
wire     [31:0] n22037;
wire     [31:0] n22038;
wire     [31:0] n22039;
wire     [31:0] n22040;
wire     [31:0] n22041;
wire     [31:0] n22042;
wire     [31:0] n22043;
wire     [31:0] n22044;
wire     [31:0] n22045;
wire     [31:0] n22046;
wire     [31:0] n22047;
wire     [31:0] n22048;
wire     [31:0] n22049;
wire     [31:0] n22050;
wire     [31:0] n22051;
wire     [31:0] n22052;
wire     [31:0] n22053;
wire     [31:0] n22054;
wire     [31:0] n22055;
wire     [31:0] n22056;
wire     [31:0] n22057;
wire     [31:0] n22058;
wire     [31:0] n22059;
wire     [31:0] n22060;
wire     [31:0] n22061;
wire     [31:0] n22062;
wire     [31:0] n22063;
wire     [31:0] n22064;
wire     [31:0] n22065;
wire     [31:0] n22066;
wire     [31:0] n22067;
wire     [31:0] n22068;
wire     [31:0] n22069;
wire     [31:0] n22070;
wire     [31:0] n22071;
wire     [31:0] n22072;
wire     [31:0] n22073;
wire     [31:0] n22074;
wire     [31:0] n22075;
wire     [31:0] n22076;
wire     [31:0] n22077;
wire     [31:0] n22078;
wire     [31:0] n22079;
wire     [31:0] n22080;
wire     [31:0] n22081;
wire     [31:0] n22082;
wire     [31:0] n22083;
wire     [31:0] n22084;
wire     [31:0] n22085;
wire     [31:0] n22086;
wire     [31:0] n22087;
wire     [31:0] n22088;
wire     [31:0] n22089;
wire     [31:0] n22090;
wire     [31:0] n22091;
wire     [31:0] n22092;
wire     [31:0] n22093;
wire     [31:0] n22094;
wire     [31:0] n22095;
wire     [31:0] n22096;
wire     [31:0] n22097;
wire     [31:0] n22098;
wire     [31:0] n22099;
wire     [31:0] n22100;
wire     [31:0] n22101;
wire     [31:0] n22102;
wire     [31:0] n22103;
wire     [31:0] n22104;
wire            n22105;
wire            n22106;
wire     [31:0] n22107;
wire     [31:0] n22108;
wire     [31:0] n22109;
wire     [31:0] n22110;
wire     [31:0] n22111;
wire     [31:0] n22112;
wire     [31:0] n22113;
wire     [31:0] n22114;
wire     [31:0] n22115;
wire     [31:0] n22116;
wire     [31:0] n22117;
wire     [31:0] n22118;
wire     [31:0] n22119;
wire     [31:0] n22120;
wire     [31:0] n22121;
wire     [31:0] n22122;
wire     [31:0] n22123;
wire     [31:0] n22124;
wire     [31:0] n22125;
wire     [31:0] n22126;
wire     [31:0] n22127;
wire     [31:0] n22128;
wire     [31:0] n22129;
wire     [31:0] n22130;
wire     [31:0] n22131;
wire     [31:0] n22132;
wire     [31:0] n22133;
wire     [31:0] n22134;
wire     [31:0] n22135;
wire     [31:0] n22136;
wire     [31:0] n22137;
wire     [31:0] n22138;
wire     [31:0] n22139;
wire            n22140;
wire            n22141;
wire            n22142;
wire            n22143;
wire            n22144;
wire            n22145;
wire            n22146;
wire            n22147;
wire            n22148;
wire            n22149;
wire            n22150;
wire            n22151;
wire            n22152;
wire            n22153;
wire            n22154;
wire            n22155;
wire            n22156;
wire            n22157;
wire            n22158;
wire            n22159;
wire            n22160;
wire            n22161;
wire            n22162;
wire            n22163;
wire            n22164;
wire            n22165;
wire            n22166;
wire            n22167;
wire            n22168;
wire            n22169;
wire            n22170;
wire            n22171;
wire            n22172;
wire            n22173;
wire            n22174;
wire            n22175;
wire            n22176;
wire            n22177;
wire            n22178;
wire            n22179;
wire            n22180;
wire            n22181;
wire            n22182;
wire            n22183;
wire            n22184;
wire            n22185;
wire            n22186;
wire            n22187;
wire            n22188;
wire            n22189;
wire            n22190;
wire            n22191;
wire            n22192;
wire            n22193;
wire            n22194;
wire            n22195;
wire            n22196;
wire            n22197;
wire            n22198;
wire            n22199;
wire            n22200;
wire            n22201;
wire            n22202;
wire            n22203;
wire            n22204;
wire            n22205;
wire            n22206;
wire            n22207;
wire            n22208;
wire            n22209;
wire            n22210;
wire            n22211;
wire            n22212;
wire            n22213;
wire            n22214;
wire            n22215;
wire            n22216;
wire            n22217;
wire            n22218;
wire            n22219;
wire            n22220;
wire            n22221;
wire            n22222;
wire            n22223;
wire            n22224;
wire            n22225;
wire            n22226;
wire            n22227;
wire            n22228;
wire            n22229;
wire            n22230;
wire            n22231;
wire            n22232;
wire            n22233;
wire            n22234;
wire            n22235;
wire            n22236;
wire            n22237;
wire            n22238;
wire            n22239;
wire            n22240;
wire            n22241;
wire            n22242;
wire            n22243;
wire            n22244;
wire            n22245;
wire            n22246;
wire            n22247;
wire            n22248;
wire            n22249;
wire            n22250;
wire            n22251;
wire            n22252;
wire            n22253;
wire            n22254;
wire            n22255;
wire            n22256;
wire            n22257;
wire            n22258;
wire            n22259;
wire            n22260;
wire            n22261;
wire            n22262;
wire            n22263;
wire            n22264;
wire            n22265;
wire            n22266;
wire            n22267;
wire            n22268;
wire            n22269;
wire            n22270;
wire            n22271;
wire            n22272;
wire            n22273;
wire            n22274;
wire            n22275;
wire            n22276;
wire            n22277;
wire            n22278;
wire            n22279;
wire            n22280;
wire            n22281;
wire            n22282;
wire            n22283;
wire            n22284;
wire            n22285;
wire            n22286;
wire            n22287;
wire            n22288;
wire            n22289;
wire            n22290;
wire            n22291;
wire            n22292;
wire            n22293;
wire            n22294;
wire            n22295;
wire            n22296;
wire            n22297;
wire            n22298;
wire            n22299;
wire            n22300;
wire            n22301;
wire            n22302;
wire            n22303;
wire            n22304;
wire            n22305;
wire            n22306;
wire            n22307;
wire            n22308;
wire            n22309;
wire            n22310;
wire            n22311;
wire            n22312;
wire            n22313;
wire            n22314;
wire            n22315;
wire            n22316;
wire            n22317;
wire            n22318;
wire            n22319;
wire            n22320;
wire            n22321;
wire            n22322;
wire            n22323;
wire            n22324;
wire            n22325;
wire            n22326;
wire            n22327;
wire            n22328;
wire            n22329;
wire            n22330;
wire            n22331;
wire            n22332;
wire            n22333;
wire            n22334;
wire            n22335;
wire            n22336;
wire            n22337;
wire            n22338;
wire            n22339;
wire            n22340;
wire            n22341;
wire            n22342;
wire            n22343;
wire            n22344;
wire            n22345;
wire            n22346;
wire            n22347;
wire            n22348;
wire            n22349;
wire            n22350;
wire            n22351;
wire            n22352;
wire            n22353;
wire            n22354;
wire            n22355;
wire            n22356;
wire            n22357;
wire            n22358;
wire            n22359;
wire            n22360;
wire            n22361;
wire            n22362;
wire            n22363;
wire            n22364;
wire            n22365;
wire            n22366;
wire            n22367;
wire            n22368;
wire            n22369;
wire            n22370;
wire            n22371;
wire            n22372;
wire            n22373;
wire            n22374;
wire            n22375;
wire            n22376;
wire            n22377;
wire            n22378;
wire            n22379;
wire            n22380;
wire            n22381;
wire            n22382;
wire            n22383;
wire            n22384;
wire            n22385;
wire            n22386;
wire            n22387;
wire            n22388;
wire            n22389;
wire            n22390;
wire            n22391;
wire            n22392;
wire            n22393;
wire            n22394;
wire            n22395;
wire            n22396;
wire            n22397;
wire            n22398;
wire            n22399;
wire            n22400;
wire            n22401;
wire            n22402;
wire            n22403;
wire            n22404;
wire            n22405;
wire            n22406;
wire            n22407;
wire            n22408;
wire            n22409;
wire            n22410;
wire            n22411;
wire            n22412;
wire            n22413;
wire            n22414;
wire            n22415;
wire            n22416;
wire            n22417;
wire            n22418;
wire            n22419;
wire            n22420;
wire            n22421;
wire            n22422;
wire            n22423;
wire            n22424;
wire            n22425;
wire            n22426;
wire            n22427;
wire            n22428;
wire            n22429;
wire            n22430;
wire            n22431;
wire            n22432;
wire            n22433;
wire            n22434;
wire            n22435;
wire            n22436;
wire            n22437;
wire            n22438;
wire            n22439;
wire            n22440;
wire            n22441;
wire            n22442;
wire            n22443;
wire            n22444;
wire            n22445;
wire            n22446;
wire            n22447;
wire            n22448;
wire            n22449;
wire            n22450;
wire            n22451;
wire            n22452;
wire            n22453;
wire            n22454;
wire            n22455;
wire            n22456;
wire            n22457;
wire            n22458;
wire            n22459;
wire            n22460;
wire            n22461;
wire            n22462;
wire            n22463;
wire            n22464;
wire            n22465;
wire            n22466;
wire            n22467;
wire            n22468;
wire            n22469;
wire            n22470;
wire            n22471;
wire            n22472;
wire            n22473;
wire            n22474;
wire            n22475;
wire            n22476;
wire            n22477;
wire            n22478;
wire            n22479;
wire            n22480;
wire            n22481;
wire            n22482;
wire            n22483;
wire            n22484;
wire            n22485;
wire            n22486;
wire            n22487;
wire            n22488;
wire            n22489;
wire            n22490;
wire            n22491;
wire            n22492;
wire            n22493;
wire            n22494;
wire            n22495;
wire            n22496;
wire            n22497;
wire            n22498;
wire            n22499;
wire            n22500;
wire            n22501;
wire            n22502;
wire            n22503;
wire            n22504;
wire            n22505;
wire            n22506;
wire            n22507;
wire            n22508;
wire            n22509;
wire            n22510;
wire            n22511;
wire            n22512;
wire            n22513;
wire            n22514;
wire            n22515;
wire            n22516;
wire            n22517;
wire            n22518;
wire            n22519;
wire            n22520;
wire            n22521;
wire            n22522;
wire            n22523;
wire            n22524;
wire            n22525;
wire            n22526;
wire            n22527;
wire            n22528;
wire            n22529;
wire            n22530;
wire            n22531;
wire            n22532;
wire            n22533;
wire            n22534;
wire            n22535;
wire            n22536;
wire            n22537;
wire            n22538;
wire            n22539;
wire            n22540;
wire            n22541;
wire            n22542;
wire            n22543;
wire            n22544;
wire            n22545;
wire            n22546;
wire            n22547;
wire            n22548;
wire            n22549;
wire            n22550;
wire            n22551;
wire            n22552;
wire            n22553;
wire            n22554;
wire            n22555;
wire            n22556;
wire            n22557;
wire            n22558;
wire            n22559;
wire            n22560;
wire            n22561;
wire            n22562;
wire            n22563;
wire            n22564;
wire            n22565;
wire            n22566;
wire            n22567;
wire            n22568;
wire            n22569;
wire            n22570;
wire            n22571;
wire            n22572;
wire            n22573;
wire            n22574;
wire            n22575;
wire            n22576;
wire            n22577;
wire            n22578;
wire            n22579;
wire            n22580;
wire            n22581;
wire            n22582;
wire            n22583;
wire            n22584;
wire            n22585;
wire            n22586;
wire            n22587;
wire            n22588;
wire            n22589;
wire            n22590;
wire            n22591;
wire            n22592;
wire            n22593;
wire            n22594;
wire            n22595;
wire            n22596;
wire            n22597;
wire            n22598;
wire            n22599;
wire            n22600;
wire            n22601;
wire            n22602;
wire            n22603;
wire            n22604;
wire            n22605;
wire            n22606;
wire            n22607;
wire            n22608;
wire            n22609;
wire            n22610;
wire            n22611;
wire            n22612;
wire            n22613;
wire            n22614;
wire            n22615;
wire            n22616;
wire            n22617;
wire            n22618;
wire            n22619;
wire            n22620;
wire            n22621;
wire            n22622;
wire            n22623;
wire            n22624;
wire            n22625;
wire            n22626;
wire            n22627;
wire            n22628;
wire            n22629;
wire            n22630;
wire            n22631;
wire            n22632;
wire            n22633;
wire            n22634;
wire            n22635;
wire            n22636;
wire            n22637;
wire            n22638;
wire            n22639;
wire            n22640;
wire            n22641;
wire            n22642;
wire            n22643;
wire            n22644;
wire            n22645;
wire            n22646;
wire            n22647;
wire            n22648;
wire            n22649;
wire            n22650;
wire            n22651;
wire            n22652;
wire            n22653;
wire            n22654;
wire            n22655;
wire            n22656;
wire            n22657;
wire            n22658;
wire            n22659;
wire            n22660;
wire            n22661;
wire            n22662;
wire            n22663;
wire            n22664;
wire            n22665;
wire            n22666;
wire            n22667;
wire     [31:0] n22668;
wire     [31:0] n22669;
wire     [31:0] n22670;
wire     [31:0] n22671;
wire     [31:0] n22672;
wire     [31:0] n22673;
wire     [31:0] n22674;
wire     [31:0] n22675;
wire     [31:0] n22676;
wire     [31:0] n22677;
wire     [31:0] n22678;
wire     [31:0] n22679;
wire     [31:0] n22680;
wire     [31:0] n22681;
wire     [31:0] n22682;
wire     [31:0] n22683;
wire     [31:0] n22684;
wire     [31:0] n22685;
wire     [31:0] n22686;
wire     [31:0] n22687;
wire     [31:0] n22688;
wire     [31:0] n22689;
wire     [31:0] n22690;
wire     [31:0] n22691;
wire     [31:0] n22692;
wire     [31:0] n22693;
wire     [31:0] n22694;
wire     [31:0] n22695;
wire     [31:0] n22696;
wire     [31:0] n22697;
wire     [31:0] n22698;
wire     [31:0] n22699;
wire     [31:0] n22700;
wire     [31:0] n22701;
wire     [31:0] n22702;
wire     [31:0] n22703;
wire     [31:0] n22704;
wire     [31:0] n22705;
wire     [31:0] n22706;
wire     [31:0] n22707;
wire     [31:0] n22708;
wire     [31:0] n22709;
wire     [31:0] n22710;
wire     [31:0] n22711;
wire     [31:0] n22712;
wire     [31:0] n22713;
wire     [31:0] n22714;
wire     [31:0] n22715;
wire     [31:0] n22716;
wire     [31:0] n22717;
wire     [31:0] n22718;
wire     [31:0] n22719;
wire     [31:0] n22720;
wire     [31:0] n22721;
wire     [31:0] n22722;
wire     [31:0] n22723;
wire     [31:0] n22724;
wire     [31:0] n22725;
wire     [31:0] n22726;
wire     [31:0] n22727;
wire     [31:0] n22728;
wire     [31:0] n22729;
wire     [31:0] n22730;
wire     [31:0] n22731;
wire     [31:0] n22732;
wire     [31:0] n22733;
wire     [31:0] n22734;
wire     [31:0] n22735;
wire     [31:0] n22736;
wire     [31:0] n22737;
wire     [31:0] n22738;
wire     [31:0] n22739;
wire     [31:0] n22740;
wire     [31:0] n22741;
wire     [31:0] n22742;
wire     [31:0] n22743;
wire     [31:0] n22744;
wire     [31:0] n22745;
wire     [31:0] n22746;
wire     [31:0] n22747;
wire     [31:0] n22748;
wire     [31:0] n22749;
wire     [31:0] n22750;
wire     [31:0] n22751;
wire     [31:0] n22752;
wire     [31:0] n22753;
wire     [31:0] n22754;
wire     [31:0] n22755;
wire     [31:0] n22756;
wire     [31:0] n22757;
wire     [31:0] n22758;
wire     [31:0] n22759;
wire     [31:0] n22760;
wire     [31:0] n22761;
wire     [31:0] n22762;
wire     [31:0] n22763;
wire     [31:0] n22764;
wire     [31:0] n22765;
wire     [31:0] n22766;
wire     [31:0] n22767;
wire     [31:0] n22768;
wire     [31:0] n22769;
wire     [31:0] n22770;
wire     [31:0] n22771;
wire     [31:0] n22772;
wire     [31:0] n22773;
wire     [31:0] n22774;
wire     [31:0] n22775;
wire     [31:0] n22776;
wire     [31:0] n22777;
wire     [31:0] n22778;
wire     [31:0] n22779;
wire     [31:0] n22780;
wire     [31:0] n22781;
wire     [31:0] n22782;
wire     [31:0] n22783;
wire     [31:0] n22784;
wire     [31:0] n22785;
wire     [31:0] n22786;
wire     [31:0] n22787;
wire     [31:0] n22788;
wire     [31:0] n22789;
wire     [31:0] n22790;
wire     [31:0] n22791;
wire     [31:0] n22792;
wire     [31:0] n22793;
wire     [31:0] n22794;
wire     [31:0] n22795;
wire     [31:0] n22796;
wire     [31:0] n22797;
wire     [31:0] n22798;
wire     [31:0] n22799;
wire     [31:0] n22800;
wire     [31:0] n22801;
wire     [31:0] n22802;
wire     [31:0] n22803;
wire     [31:0] n22804;
wire     [31:0] n22805;
wire     [31:0] n22806;
wire     [31:0] n22807;
wire     [31:0] n22808;
wire     [31:0] n22809;
wire     [31:0] n22810;
wire     [31:0] n22811;
wire     [31:0] n22812;
wire     [31:0] n22813;
wire     [31:0] n22814;
wire     [31:0] n22815;
wire     [31:0] n22816;
wire     [31:0] n22817;
wire     [31:0] n22818;
wire     [31:0] n22819;
wire     [31:0] n22820;
wire     [31:0] n22821;
wire     [31:0] n22822;
wire     [31:0] n22823;
wire     [31:0] n22824;
wire     [31:0] n22825;
wire     [31:0] n22826;
wire     [31:0] n22827;
wire     [31:0] n22828;
wire     [31:0] n22829;
wire     [31:0] n22830;
wire     [31:0] n22831;
wire     [31:0] n22832;
wire     [31:0] n22833;
wire     [31:0] n22834;
wire     [31:0] n22835;
wire     [31:0] n22836;
wire     [31:0] n22837;
wire     [31:0] n22838;
wire     [31:0] n22839;
wire     [31:0] n22840;
wire     [31:0] n22841;
wire     [31:0] n22842;
wire     [31:0] n22843;
wire     [31:0] n22844;
wire     [31:0] n22845;
wire     [31:0] n22846;
wire     [31:0] n22847;
wire     [31:0] n22848;
wire     [31:0] n22849;
wire     [31:0] n22850;
wire     [31:0] n22851;
wire     [31:0] n22852;
wire     [31:0] n22853;
wire     [31:0] n22854;
wire     [31:0] n22855;
wire     [31:0] n22856;
wire     [31:0] n22857;
wire     [31:0] n22858;
wire     [31:0] n22859;
wire     [31:0] n22860;
wire     [31:0] n22861;
wire     [31:0] n22862;
wire     [31:0] n22863;
wire     [31:0] n22864;
wire     [31:0] n22865;
wire     [31:0] n22866;
wire     [31:0] n22867;
wire     [31:0] n22868;
wire     [31:0] n22869;
wire     [31:0] n22870;
wire     [31:0] n22871;
wire     [31:0] n22872;
wire     [31:0] n22873;
wire     [31:0] n22874;
wire     [31:0] n22875;
wire     [31:0] n22876;
wire     [31:0] n22877;
wire     [31:0] n22878;
wire     [31:0] n22879;
wire     [31:0] n22880;
wire     [31:0] n22881;
wire     [31:0] n22882;
wire     [31:0] n22883;
wire     [31:0] n22884;
wire     [31:0] n22885;
wire     [31:0] n22886;
wire     [31:0] n22887;
wire     [31:0] n22888;
wire     [31:0] n22889;
wire     [31:0] n22890;
wire     [31:0] n22891;
wire     [31:0] n22892;
wire     [31:0] n22893;
wire     [31:0] n22894;
wire     [31:0] n22895;
wire     [31:0] n22896;
wire     [31:0] n22897;
wire     [31:0] n22898;
wire     [31:0] n22899;
wire     [31:0] n22900;
wire     [31:0] n22901;
wire     [31:0] n22902;
wire     [31:0] n22903;
wire     [31:0] n22904;
wire     [31:0] n22905;
wire     [31:0] n22906;
wire     [31:0] n22907;
wire     [31:0] n22908;
wire     [31:0] n22909;
wire     [31:0] n22910;
wire     [31:0] n22911;
wire     [31:0] n22912;
wire     [31:0] n22913;
wire     [31:0] n22914;
wire     [31:0] n22915;
wire     [31:0] n22916;
wire     [31:0] n22917;
wire     [31:0] n22918;
wire     [31:0] n22919;
wire     [31:0] n22920;
wire     [31:0] n22921;
wire     [31:0] n22922;
wire     [31:0] n22923;
wire     [31:0] n22924;
wire     [31:0] n22925;
wire     [31:0] n22926;
wire     [31:0] n22927;
wire     [31:0] n22928;
wire     [31:0] n22929;
wire     [31:0] n22930;
wire     [31:0] n22931;
wire     [31:0] n22932;
wire     [31:0] n22933;
wire     [31:0] n22934;
wire     [31:0] n22935;
wire     [31:0] n22936;
wire     [31:0] n22937;
wire     [31:0] n22938;
wire     [31:0] n22939;
wire     [31:0] n22940;
wire     [31:0] n22941;
wire     [31:0] n22942;
wire     [31:0] n22943;
wire     [31:0] n22944;
wire     [31:0] n22945;
wire     [31:0] n22946;
wire     [31:0] n22947;
wire     [31:0] n22948;
wire     [31:0] n22949;
wire     [31:0] n22950;
wire     [31:0] n22951;
wire     [31:0] n22952;
wire     [31:0] n22953;
wire     [31:0] n22954;
wire     [31:0] n22955;
wire     [31:0] n22956;
wire     [31:0] n22957;
wire     [31:0] n22958;
wire     [31:0] n22959;
wire     [31:0] n22960;
wire     [31:0] n22961;
wire     [31:0] n22962;
wire     [31:0] n22963;
wire     [31:0] n22964;
wire     [31:0] n22965;
wire     [31:0] n22966;
wire     [31:0] n22967;
wire     [31:0] n22968;
wire     [31:0] n22969;
wire     [31:0] n22970;
wire     [31:0] n22971;
wire     [31:0] n22972;
wire     [31:0] n22973;
wire     [31:0] n22974;
wire     [31:0] n22975;
wire     [31:0] n22976;
wire     [31:0] n22977;
wire     [31:0] n22978;
wire     [31:0] n22979;
wire     [31:0] n22980;
wire     [31:0] n22981;
wire     [31:0] n22982;
wire     [31:0] n22983;
wire     [31:0] n22984;
wire     [31:0] n22985;
wire     [31:0] n22986;
wire     [31:0] n22987;
wire     [31:0] n22988;
wire     [31:0] n22989;
wire     [31:0] n22990;
wire     [31:0] n22991;
wire     [31:0] n22992;
wire     [31:0] n22993;
wire     [31:0] n22994;
wire     [31:0] n22995;
wire     [31:0] n22996;
wire     [31:0] n22997;
wire     [31:0] n22998;
wire     [31:0] n22999;
wire     [31:0] n23000;
wire     [31:0] n23001;
wire     [31:0] n23002;
wire     [31:0] n23003;
wire     [31:0] n23004;
wire     [31:0] n23005;
wire     [31:0] n23006;
wire     [31:0] n23007;
wire     [31:0] n23008;
wire     [31:0] n23009;
wire     [31:0] n23010;
wire     [31:0] n23011;
wire     [31:0] n23012;
wire     [31:0] n23013;
wire     [31:0] n23014;
wire     [31:0] n23015;
wire     [31:0] n23016;
wire     [31:0] n23017;
wire     [31:0] n23018;
wire     [31:0] n23019;
wire     [31:0] n23020;
wire     [31:0] n23021;
wire     [31:0] n23022;
wire     [31:0] n23023;
wire     [31:0] n23024;
wire     [31:0] n23025;
wire     [31:0] n23026;
wire     [31:0] n23027;
wire     [31:0] n23028;
wire     [31:0] n23029;
wire     [31:0] n23030;
wire     [31:0] n23031;
wire     [31:0] n23032;
wire     [31:0] n23033;
wire     [31:0] n23034;
wire     [31:0] n23035;
wire     [31:0] n23036;
wire     [31:0] n23037;
wire     [31:0] n23038;
wire     [31:0] n23039;
wire     [31:0] n23040;
wire     [31:0] n23041;
wire     [31:0] n23042;
wire     [31:0] n23043;
wire     [31:0] n23044;
wire     [31:0] n23045;
wire     [31:0] n23046;
wire     [31:0] n23047;
wire     [31:0] n23048;
wire     [31:0] n23049;
wire     [31:0] n23050;
wire     [31:0] n23051;
wire     [31:0] n23052;
wire     [31:0] n23053;
wire     [31:0] n23054;
wire     [31:0] n23055;
wire     [31:0] n23056;
wire     [31:0] n23057;
wire     [31:0] n23058;
wire     [31:0] n23059;
wire     [31:0] n23060;
wire     [31:0] n23061;
wire     [31:0] n23062;
wire     [31:0] n23063;
wire     [31:0] n23064;
wire     [31:0] n23065;
wire     [31:0] n23066;
wire     [31:0] n23067;
wire     [31:0] n23068;
wire     [31:0] n23069;
wire     [31:0] n23070;
wire     [31:0] n23071;
wire     [31:0] n23072;
wire     [31:0] n23073;
wire     [31:0] n23074;
wire     [31:0] n23075;
wire     [31:0] n23076;
wire     [31:0] n23077;
wire     [31:0] n23078;
wire     [31:0] n23079;
wire     [31:0] n23080;
wire     [31:0] n23081;
wire     [31:0] n23082;
wire     [31:0] n23083;
wire     [31:0] n23084;
wire     [31:0] n23085;
wire     [31:0] n23086;
wire     [31:0] n23087;
wire     [31:0] n23088;
wire     [31:0] n23089;
wire     [31:0] n23090;
wire     [31:0] n23091;
wire     [31:0] n23092;
wire     [31:0] n23093;
wire     [31:0] n23094;
wire     [31:0] n23095;
wire     [31:0] n23096;
wire     [31:0] n23097;
wire     [31:0] n23098;
wire     [31:0] n23099;
wire     [31:0] n23100;
wire     [31:0] n23101;
wire     [31:0] n23102;
wire     [31:0] n23103;
wire     [31:0] n23104;
wire     [31:0] n23105;
wire     [31:0] n23106;
wire     [31:0] n23107;
wire     [31:0] n23108;
wire     [31:0] n23109;
wire     [31:0] n23110;
wire     [31:0] n23111;
wire     [31:0] n23112;
wire     [31:0] n23113;
wire     [31:0] n23114;
wire     [31:0] n23115;
wire     [31:0] n23116;
wire     [31:0] n23117;
wire     [31:0] n23118;
wire     [31:0] n23119;
wire     [31:0] n23120;
wire     [31:0] n23121;
wire     [31:0] n23122;
wire     [31:0] n23123;
wire     [31:0] n23124;
wire     [31:0] n23125;
wire     [31:0] n23126;
wire     [31:0] n23127;
wire     [31:0] n23128;
wire     [31:0] n23129;
wire     [31:0] n23130;
wire     [31:0] n23131;
wire     [31:0] n23132;
wire     [31:0] n23133;
wire     [31:0] n23134;
wire     [31:0] n23135;
wire     [31:0] n23136;
wire     [31:0] n23137;
wire     [31:0] n23138;
wire     [31:0] n23139;
wire     [31:0] n23140;
wire     [31:0] n23141;
wire     [31:0] n23142;
wire     [31:0] n23143;
wire     [31:0] n23144;
wire     [31:0] n23145;
wire     [31:0] n23146;
wire     [31:0] n23147;
wire     [31:0] n23148;
wire     [31:0] n23149;
wire     [31:0] n23150;
wire     [31:0] n23151;
wire     [31:0] n23152;
wire     [31:0] n23153;
wire     [31:0] n23154;
wire     [31:0] n23155;
wire     [31:0] n23156;
wire     [31:0] n23157;
wire     [31:0] n23158;
wire     [31:0] n23159;
wire     [31:0] n23160;
wire     [31:0] n23161;
wire     [31:0] n23162;
wire     [31:0] n23163;
wire     [31:0] n23164;
wire     [31:0] n23165;
wire     [31:0] n23166;
wire     [31:0] n23167;
wire     [31:0] n23168;
wire     [31:0] n23169;
wire     [31:0] n23170;
wire     [31:0] n23171;
wire     [31:0] n23172;
wire     [31:0] n23173;
wire     [31:0] n23174;
wire     [31:0] n23175;
wire     [31:0] n23176;
wire     [31:0] n23177;
wire     [31:0] n23178;
wire     [31:0] n23179;
wire     [31:0] n23180;
wire     [31:0] n23181;
wire     [31:0] n23182;
wire     [31:0] n23183;
wire     [31:0] n23184;
wire     [31:0] n23185;
wire     [31:0] n23186;
wire     [31:0] n23187;
wire     [31:0] n23188;
wire     [31:0] n23189;
wire            n23190;
wire            n23191;
wire            n23192;
wire            n23193;
wire            n23194;
wire            n23195;
wire            n23196;
wire            n23197;
wire            n23198;
wire            n23199;
wire            n23200;
wire            n23201;
wire            n23202;
wire            n23203;
wire            n23204;
wire            n23205;
wire            n23206;
wire            n23207;
wire            n23208;
wire            n23209;
wire            n23210;
wire            n23211;
wire            n23212;
wire            n23213;
wire            n23214;
wire            n23215;
wire            n23216;
wire            n23217;
wire            n23218;
wire            n23219;
wire            n23220;
wire            n23221;
wire            n23222;
wire            n23223;
wire            n23224;
wire            n23225;
wire            n23226;
wire            n23227;
wire            n23228;
wire            n23229;
wire            n23230;
wire            n23231;
wire            n23232;
wire            n23233;
wire            n23234;
wire            n23235;
wire            n23236;
wire            n23237;
wire            n23238;
wire            n23239;
wire            n23240;
wire            n23241;
wire            n23242;
wire            n23243;
wire            n23244;
wire            n23245;
wire            n23246;
wire            n23247;
wire            n23248;
wire            n23249;
wire            n23250;
wire            n23251;
wire            n23252;
wire            n23253;
wire            n23254;
wire            n23255;
wire            n23256;
wire            n23257;
wire            n23258;
wire            n23259;
wire            n23260;
wire            n23261;
wire            n23262;
wire            n23263;
wire            n23264;
wire            n23265;
wire            n23266;
wire            n23267;
wire            n23268;
wire            n23269;
wire            n23270;
wire            n23271;
wire            n23272;
wire            n23273;
wire            n23274;
wire            n23275;
wire            n23276;
wire            n23277;
wire            n23278;
wire            n23279;
wire            n23280;
wire            n23281;
wire            n23282;
wire            n23283;
wire            n23284;
wire            n23285;
wire            n23286;
wire            n23287;
wire            n23288;
wire            n23289;
wire            n23290;
wire            n23291;
wire            n23292;
wire            n23293;
wire            n23294;
wire            n23295;
wire            n23296;
wire            n23297;
wire            n23298;
wire            n23299;
wire            n23300;
wire            n23301;
wire            n23302;
wire            n23303;
wire            n23304;
wire            n23305;
wire            n23306;
wire            n23307;
wire            n23308;
wire            n23309;
wire            n23310;
wire            n23311;
wire            n23312;
wire            n23313;
wire            n23314;
wire            n23315;
wire            n23316;
wire            n23317;
wire            n23318;
wire            n23319;
wire            n23320;
wire            n23321;
wire            n23322;
wire            n23323;
wire            n23324;
wire            n23325;
wire            n23326;
wire            n23327;
wire            n23328;
wire            n23329;
wire            n23330;
wire            n23331;
wire            n23332;
wire            n23333;
wire            n23334;
wire            n23335;
wire            n23336;
wire            n23337;
wire            n23338;
wire            n23339;
wire            n23340;
wire            n23341;
wire            n23342;
wire            n23343;
wire            n23344;
wire            n23345;
wire            n23346;
wire            n23347;
wire            n23348;
wire            n23349;
wire            n23350;
wire            n23351;
wire            n23352;
wire            n23353;
wire            n23354;
wire            n23355;
wire            n23356;
wire            n23357;
wire            n23358;
wire            n23359;
wire            n23360;
wire            n23361;
wire            n23362;
wire            n23363;
wire            n23364;
wire            n23365;
wire            n23366;
wire            n23367;
wire            n23368;
wire            n23369;
wire            n23370;
wire            n23371;
wire            n23372;
wire            n23373;
wire            n23374;
wire            n23375;
wire            n23376;
wire            n23377;
wire            n23378;
wire            n23379;
wire            n23380;
wire            n23381;
wire            n23382;
wire            n23383;
wire            n23384;
wire            n23385;
wire            n23386;
wire            n23387;
wire            n23388;
wire            n23389;
wire            n23390;
wire            n23391;
wire            n23392;
wire            n23393;
wire            n23394;
wire            n23395;
wire            n23396;
wire            n23397;
wire            n23398;
wire            n23399;
wire            n23400;
wire            n23401;
wire            n23402;
wire            n23403;
wire            n23404;
wire            n23405;
wire            n23406;
wire            n23407;
wire            n23408;
wire            n23409;
wire            n23410;
wire            n23411;
wire            n23412;
wire            n23413;
wire            n23414;
wire            n23415;
wire            n23416;
wire            n23417;
wire            n23418;
wire            n23419;
wire            n23420;
wire            n23421;
wire            n23422;
wire            n23423;
wire            n23424;
wire            n23425;
wire            n23426;
wire            n23427;
wire            n23428;
wire            n23429;
wire            n23430;
wire            n23431;
wire            n23432;
wire            n23433;
wire            n23434;
wire            n23435;
wire            n23436;
wire            n23437;
wire            n23438;
wire            n23439;
wire            n23440;
wire            n23441;
wire            n23442;
wire            n23443;
wire            n23444;
wire            n23445;
wire            n23446;
wire            n23447;
wire            n23448;
wire            n23449;
wire            n23450;
wire            n23451;
wire            n23452;
wire            n23453;
wire            n23454;
wire            n23455;
wire            n23456;
wire            n23457;
wire            n23458;
wire            n23459;
wire            n23460;
wire            n23461;
wire            n23462;
wire            n23463;
wire            n23464;
wire            n23465;
wire            n23466;
wire            n23467;
wire            n23468;
wire            n23469;
wire            n23470;
wire            n23471;
wire            n23472;
wire            n23473;
wire            n23474;
wire            n23475;
wire            n23476;
wire            n23477;
wire            n23478;
wire            n23479;
wire            n23480;
wire            n23481;
wire            n23482;
wire            n23483;
wire            n23484;
wire            n23485;
wire            n23486;
wire            n23487;
wire            n23488;
wire            n23489;
wire            n23490;
wire            n23491;
wire            n23492;
wire            n23493;
wire            n23494;
wire            n23495;
wire            n23496;
wire            n23497;
wire            n23498;
wire            n23499;
wire            n23500;
wire            n23501;
wire            n23502;
wire            n23503;
wire            n23504;
wire            n23505;
wire            n23506;
wire            n23507;
wire            n23508;
wire            n23509;
wire            n23510;
wire            n23511;
wire            n23512;
wire            n23513;
wire            n23514;
wire            n23515;
wire            n23516;
wire            n23517;
wire            n23518;
wire            n23519;
wire            n23520;
wire            n23521;
wire            n23522;
wire            n23523;
wire            n23524;
wire            n23525;
wire            n23526;
wire            n23527;
wire            n23528;
wire            n23529;
wire            n23530;
wire            n23531;
wire            n23532;
wire            n23533;
wire            n23534;
wire            n23535;
wire            n23536;
wire            n23537;
wire            n23538;
wire            n23539;
wire            n23540;
wire            n23541;
wire            n23542;
wire            n23543;
wire            n23544;
wire            n23545;
wire            n23546;
wire            n23547;
wire            n23548;
wire            n23549;
wire            n23550;
wire            n23551;
wire            n23552;
wire            n23553;
wire            n23554;
wire            n23555;
wire            n23556;
wire            n23557;
wire            n23558;
wire            n23559;
wire            n23560;
wire            n23561;
wire            n23562;
wire            n23563;
wire            n23564;
wire            n23565;
wire            n23566;
wire            n23567;
wire            n23568;
wire            n23569;
wire            n23570;
wire            n23571;
wire            n23572;
wire            n23573;
wire            n23574;
wire            n23575;
wire            n23576;
wire            n23577;
wire            n23578;
wire            n23579;
wire            n23580;
wire            n23581;
wire            n23582;
wire            n23583;
wire            n23584;
wire            n23585;
wire            n23586;
wire            n23587;
wire            n23588;
wire            n23589;
wire            n23590;
wire            n23591;
wire            n23592;
wire            n23593;
wire            n23594;
wire            n23595;
wire            n23596;
wire            n23597;
wire            n23598;
wire            n23599;
wire            n23600;
wire            n23601;
wire            n23602;
wire            n23603;
wire            n23604;
wire            n23605;
wire            n23606;
wire            n23607;
wire            n23608;
wire            n23609;
wire            n23610;
wire            n23611;
wire            n23612;
wire            n23613;
wire            n23614;
wire            n23615;
wire            n23616;
wire            n23617;
wire            n23618;
wire            n23619;
wire            n23620;
wire            n23621;
wire            n23622;
wire            n23623;
wire            n23624;
wire            n23625;
wire            n23626;
wire            n23627;
wire            n23628;
wire            n23629;
wire            n23630;
wire            n23631;
wire            n23632;
wire            n23633;
wire            n23634;
wire            n23635;
wire            n23636;
wire            n23637;
wire            n23638;
wire            n23639;
wire            n23640;
wire            n23641;
wire            n23642;
wire            n23643;
wire            n23644;
wire            n23645;
wire            n23646;
wire            n23647;
wire            n23648;
wire            n23649;
wire            n23650;
wire            n23651;
wire            n23652;
wire            n23653;
wire            n23654;
wire            n23655;
wire            n23656;
wire            n23657;
wire            n23658;
wire            n23659;
wire            n23660;
wire            n23661;
wire            n23662;
wire            n23663;
wire            n23664;
wire            n23665;
wire            n23666;
wire            n23667;
wire            n23668;
wire            n23669;
wire            n23670;
wire            n23671;
wire            n23672;
wire            n23673;
wire            n23674;
wire            n23675;
wire            n23676;
wire            n23677;
wire            n23678;
wire            n23679;
wire            n23680;
wire            n23681;
wire            n23682;
wire            n23683;
wire            n23684;
wire            n23685;
wire            n23686;
wire            n23687;
wire            n23688;
wire            n23689;
wire            n23690;
wire            n23691;
wire            n23692;
wire            n23693;
wire            n23694;
wire            n23695;
wire            n23696;
wire            n23697;
wire            n23698;
wire            n23699;
wire            n23700;
wire            n23701;
wire     [31:0] n23702;
wire     [31:0] n23703;
wire     [31:0] n23704;
wire     [31:0] n23705;
wire     [31:0] n23706;
wire     [31:0] n23707;
wire     [31:0] n23708;
wire     [31:0] n23709;
wire     [31:0] n23710;
wire     [31:0] n23711;
wire     [31:0] n23712;
wire     [31:0] n23713;
wire     [31:0] n23714;
wire     [31:0] n23715;
wire     [31:0] n23716;
wire     [31:0] n23717;
wire     [31:0] n23718;
wire     [31:0] n23719;
wire     [31:0] n23720;
wire     [31:0] n23721;
wire     [31:0] n23722;
wire     [31:0] n23723;
wire     [31:0] n23724;
wire     [31:0] n23725;
wire     [31:0] n23726;
wire     [31:0] n23727;
wire     [31:0] n23728;
wire     [31:0] n23729;
wire     [31:0] n23730;
wire     [31:0] n23731;
wire     [31:0] n23732;
wire     [31:0] n23733;
wire     [31:0] n23734;
wire     [31:0] n23735;
wire     [31:0] n23736;
wire     [31:0] n23737;
wire     [31:0] n23738;
wire     [31:0] n23739;
wire     [31:0] n23740;
wire     [31:0] n23741;
wire     [31:0] n23742;
wire     [31:0] n23743;
wire     [31:0] n23744;
wire     [31:0] n23745;
wire     [31:0] n23746;
wire     [31:0] n23747;
wire     [31:0] n23748;
wire     [31:0] n23749;
wire     [31:0] n23750;
wire     [31:0] n23751;
wire     [31:0] n23752;
wire     [31:0] n23753;
wire     [31:0] n23754;
wire     [31:0] n23755;
wire     [31:0] n23756;
wire     [31:0] n23757;
wire     [31:0] n23758;
wire     [31:0] n23759;
wire     [31:0] n23760;
wire     [31:0] n23761;
wire     [31:0] n23762;
wire     [31:0] n23763;
wire     [31:0] n23764;
wire     [31:0] n23765;
wire     [31:0] n23766;
wire     [31:0] n23767;
wire     [31:0] n23768;
wire     [31:0] n23769;
wire     [31:0] n23770;
wire     [31:0] n23771;
wire     [31:0] n23772;
wire     [31:0] n23773;
wire     [31:0] n23774;
wire     [31:0] n23775;
wire     [31:0] n23776;
wire     [31:0] n23777;
wire     [31:0] n23778;
wire     [31:0] n23779;
wire     [31:0] n23780;
wire     [31:0] n23781;
wire     [31:0] n23782;
wire     [31:0] n23783;
wire     [31:0] n23784;
wire     [31:0] n23785;
wire     [31:0] n23786;
wire     [31:0] n23787;
wire     [31:0] n23788;
wire     [31:0] n23789;
wire     [31:0] n23790;
wire     [31:0] n23791;
wire     [31:0] n23792;
wire     [31:0] n23793;
wire     [31:0] n23794;
wire     [31:0] n23795;
wire     [31:0] n23796;
wire     [31:0] n23797;
wire     [31:0] n23798;
wire     [31:0] n23799;
wire     [31:0] n23800;
wire     [31:0] n23801;
wire     [31:0] n23802;
wire     [31:0] n23803;
wire     [31:0] n23804;
wire     [31:0] n23805;
wire     [31:0] n23806;
wire     [31:0] n23807;
wire     [31:0] n23808;
wire     [31:0] n23809;
wire     [31:0] n23810;
wire     [31:0] n23811;
wire     [31:0] n23812;
wire     [31:0] n23813;
wire     [31:0] n23814;
wire     [31:0] n23815;
wire     [31:0] n23816;
wire     [31:0] n23817;
wire     [31:0] n23818;
wire     [31:0] n23819;
wire     [31:0] n23820;
wire     [31:0] n23821;
wire     [31:0] n23822;
wire     [31:0] n23823;
wire     [31:0] n23824;
wire     [31:0] n23825;
wire     [31:0] n23826;
wire     [31:0] n23827;
wire     [31:0] n23828;
wire     [31:0] n23829;
wire     [31:0] n23830;
wire     [31:0] n23831;
wire     [31:0] n23832;
wire     [31:0] n23833;
wire     [31:0] n23834;
wire     [31:0] n23835;
wire     [31:0] n23836;
wire     [31:0] n23837;
wire     [31:0] n23838;
wire     [31:0] n23839;
wire     [31:0] n23840;
wire     [31:0] n23841;
wire     [31:0] n23842;
wire     [31:0] n23843;
wire     [31:0] n23844;
wire     [31:0] n23845;
wire     [31:0] n23846;
wire     [31:0] n23847;
wire     [31:0] n23848;
wire     [31:0] n23849;
wire     [31:0] n23850;
wire     [31:0] n23851;
wire     [31:0] n23852;
wire     [31:0] n23853;
wire     [31:0] n23854;
wire     [31:0] n23855;
wire     [31:0] n23856;
wire     [31:0] n23857;
wire     [31:0] n23858;
wire     [31:0] n23859;
wire     [31:0] n23860;
wire     [31:0] n23861;
wire     [31:0] n23862;
wire     [31:0] n23863;
wire     [31:0] n23864;
wire     [31:0] n23865;
wire     [31:0] n23866;
wire     [31:0] n23867;
wire     [31:0] n23868;
wire     [31:0] n23869;
wire     [31:0] n23870;
wire     [31:0] n23871;
wire     [31:0] n23872;
wire     [31:0] n23873;
wire     [31:0] n23874;
wire     [31:0] n23875;
wire     [31:0] n23876;
wire     [31:0] n23877;
wire     [31:0] n23878;
wire     [31:0] n23879;
wire     [31:0] n23880;
wire     [31:0] n23881;
wire     [31:0] n23882;
wire     [31:0] n23883;
wire     [31:0] n23884;
wire     [31:0] n23885;
wire     [31:0] n23886;
wire     [31:0] n23887;
wire     [31:0] n23888;
wire     [31:0] n23889;
wire     [31:0] n23890;
wire     [31:0] n23891;
wire     [31:0] n23892;
wire     [31:0] n23893;
wire     [31:0] n23894;
wire     [31:0] n23895;
wire     [31:0] n23896;
wire     [31:0] n23897;
wire     [31:0] n23898;
wire     [31:0] n23899;
wire     [31:0] n23900;
wire     [31:0] n23901;
wire     [31:0] n23902;
wire     [31:0] n23903;
wire     [31:0] n23904;
wire     [31:0] n23905;
wire     [31:0] n23906;
wire     [31:0] n23907;
wire     [31:0] n23908;
wire     [31:0] n23909;
wire     [31:0] n23910;
wire     [31:0] n23911;
wire     [31:0] n23912;
wire     [31:0] n23913;
wire     [31:0] n23914;
wire     [31:0] n23915;
wire     [31:0] n23916;
wire     [31:0] n23917;
wire     [31:0] n23918;
wire     [31:0] n23919;
wire     [31:0] n23920;
wire     [31:0] n23921;
wire     [31:0] n23922;
wire     [31:0] n23923;
wire     [31:0] n23924;
wire     [31:0] n23925;
wire     [31:0] n23926;
wire     [31:0] n23927;
wire     [31:0] n23928;
wire     [31:0] n23929;
wire     [31:0] n23930;
wire     [31:0] n23931;
wire     [31:0] n23932;
wire     [31:0] n23933;
wire     [31:0] n23934;
wire     [31:0] n23935;
wire     [31:0] n23936;
wire     [31:0] n23937;
wire     [31:0] n23938;
wire     [31:0] n23939;
wire     [31:0] n23940;
wire     [31:0] n23941;
wire     [31:0] n23942;
wire     [31:0] n23943;
wire     [31:0] n23944;
wire     [31:0] n23945;
wire     [31:0] n23946;
wire     [31:0] n23947;
wire     [31:0] n23948;
wire     [31:0] n23949;
wire     [31:0] n23950;
wire     [31:0] n23951;
wire     [31:0] n23952;
wire     [31:0] n23953;
wire     [31:0] n23954;
wire     [31:0] n23955;
wire     [31:0] n23956;
wire     [31:0] n23957;
wire     [31:0] n23958;
wire     [31:0] n23959;
wire     [31:0] n23960;
wire     [31:0] n23961;
wire     [31:0] n23962;
wire     [31:0] n23963;
wire     [31:0] n23964;
wire     [31:0] n23965;
wire     [31:0] n23966;
wire     [31:0] n23967;
wire     [31:0] n23968;
wire     [31:0] n23969;
wire     [31:0] n23970;
wire     [31:0] n23971;
wire     [31:0] n23972;
wire     [31:0] n23973;
wire     [31:0] n23974;
wire     [31:0] n23975;
wire     [31:0] n23976;
wire     [31:0] n23977;
wire     [31:0] n23978;
wire     [31:0] n23979;
wire     [31:0] n23980;
wire     [31:0] n23981;
wire     [31:0] n23982;
wire     [31:0] n23983;
wire     [31:0] n23984;
wire     [31:0] n23985;
wire     [31:0] n23986;
wire     [31:0] n23987;
wire     [31:0] n23988;
wire     [31:0] n23989;
wire     [31:0] n23990;
wire     [31:0] n23991;
wire     [31:0] n23992;
wire     [31:0] n23993;
wire     [31:0] n23994;
wire     [31:0] n23995;
wire     [31:0] n23996;
wire     [31:0] n23997;
wire     [31:0] n23998;
wire     [31:0] n23999;
wire     [31:0] n24000;
wire     [31:0] n24001;
wire     [31:0] n24002;
wire     [31:0] n24003;
wire     [31:0] n24004;
wire     [31:0] n24005;
wire     [31:0] n24006;
wire     [31:0] n24007;
wire     [31:0] n24008;
wire     [31:0] n24009;
wire     [31:0] n24010;
wire     [31:0] n24011;
wire     [31:0] n24012;
wire     [31:0] n24013;
wire     [31:0] n24014;
wire     [31:0] n24015;
wire     [31:0] n24016;
wire     [31:0] n24017;
wire     [31:0] n24018;
wire     [31:0] n24019;
wire     [31:0] n24020;
wire     [31:0] n24021;
wire     [31:0] n24022;
wire     [31:0] n24023;
wire     [31:0] n24024;
wire     [31:0] n24025;
wire     [31:0] n24026;
wire     [31:0] n24027;
wire     [31:0] n24028;
wire     [31:0] n24029;
wire     [31:0] n24030;
wire     [31:0] n24031;
wire     [31:0] n24032;
wire     [31:0] n24033;
wire     [31:0] n24034;
wire     [31:0] n24035;
wire     [31:0] n24036;
wire     [31:0] n24037;
wire     [31:0] n24038;
wire     [31:0] n24039;
wire     [31:0] n24040;
wire     [31:0] n24041;
wire     [31:0] n24042;
wire     [31:0] n24043;
wire     [31:0] n24044;
wire     [31:0] n24045;
wire     [31:0] n24046;
wire     [31:0] n24047;
wire     [31:0] n24048;
wire     [31:0] n24049;
wire     [31:0] n24050;
wire     [31:0] n24051;
wire     [31:0] n24052;
wire     [31:0] n24053;
wire     [31:0] n24054;
wire     [31:0] n24055;
wire     [31:0] n24056;
wire     [31:0] n24057;
wire     [31:0] n24058;
wire     [31:0] n24059;
wire     [31:0] n24060;
wire     [31:0] n24061;
wire     [31:0] n24062;
wire     [31:0] n24063;
wire     [31:0] n24064;
wire     [31:0] n24065;
wire     [31:0] n24066;
wire     [31:0] n24067;
wire     [31:0] n24068;
wire     [31:0] n24069;
wire     [31:0] n24070;
wire     [31:0] n24071;
wire     [31:0] n24072;
wire     [31:0] n24073;
wire     [31:0] n24074;
wire     [31:0] n24075;
wire     [31:0] n24076;
wire     [31:0] n24077;
wire     [31:0] n24078;
wire     [31:0] n24079;
wire     [31:0] n24080;
wire     [31:0] n24081;
wire     [31:0] n24082;
wire     [31:0] n24083;
wire     [31:0] n24084;
wire     [31:0] n24085;
wire     [31:0] n24086;
wire     [31:0] n24087;
wire     [31:0] n24088;
wire     [31:0] n24089;
wire     [31:0] n24090;
wire     [31:0] n24091;
wire     [31:0] n24092;
wire     [31:0] n24093;
wire     [31:0] n24094;
wire     [31:0] n24095;
wire     [31:0] n24096;
wire     [31:0] n24097;
wire     [31:0] n24098;
wire     [31:0] n24099;
wire     [31:0] n24100;
wire     [31:0] n24101;
wire     [31:0] n24102;
wire     [31:0] n24103;
wire     [31:0] n24104;
wire     [31:0] n24105;
wire     [31:0] n24106;
wire     [31:0] n24107;
wire     [31:0] n24108;
wire     [31:0] n24109;
wire     [31:0] n24110;
wire     [31:0] n24111;
wire     [31:0] n24112;
wire     [31:0] n24113;
wire     [31:0] n24114;
wire     [31:0] n24115;
wire     [31:0] n24116;
wire     [31:0] n24117;
wire     [31:0] n24118;
wire     [31:0] n24119;
wire     [31:0] n24120;
wire     [31:0] n24121;
wire     [31:0] n24122;
wire     [31:0] n24123;
wire     [31:0] n24124;
wire     [31:0] n24125;
wire     [31:0] n24126;
wire     [31:0] n24127;
wire     [31:0] n24128;
wire     [31:0] n24129;
wire     [31:0] n24130;
wire     [31:0] n24131;
wire     [31:0] n24132;
wire     [31:0] n24133;
wire     [31:0] n24134;
wire     [31:0] n24135;
wire     [31:0] n24136;
wire     [31:0] n24137;
wire     [31:0] n24138;
wire     [31:0] n24139;
wire     [31:0] n24140;
wire     [31:0] n24141;
wire     [31:0] n24142;
wire     [31:0] n24143;
wire     [31:0] n24144;
wire     [31:0] n24145;
wire     [31:0] n24146;
wire     [31:0] n24147;
wire     [31:0] n24148;
wire     [31:0] n24149;
wire     [31:0] n24150;
wire     [31:0] n24151;
wire     [31:0] n24152;
wire     [31:0] n24153;
wire     [31:0] n24154;
wire     [31:0] n24155;
wire     [31:0] n24156;
wire     [31:0] n24157;
wire     [31:0] n24158;
wire     [31:0] n24159;
wire     [31:0] n24160;
wire     [31:0] n24161;
wire     [31:0] n24162;
wire     [31:0] n24163;
wire     [31:0] n24164;
wire     [31:0] n24165;
wire     [31:0] n24166;
wire     [31:0] n24167;
wire     [31:0] n24168;
wire     [31:0] n24169;
wire     [31:0] n24170;
wire     [31:0] n24171;
wire     [31:0] n24172;
wire     [31:0] n24173;
wire     [31:0] n24174;
wire     [31:0] n24175;
wire     [31:0] n24176;
wire     [31:0] n24177;
wire     [31:0] n24178;
wire     [31:0] n24179;
wire     [31:0] n24180;
wire     [31:0] n24181;
wire     [31:0] n24182;
wire     [31:0] n24183;
wire     [31:0] n24184;
wire     [31:0] n24185;
wire     [31:0] n24186;
wire     [31:0] n24187;
wire     [31:0] n24188;
wire     [31:0] n24189;
wire     [31:0] n24190;
wire     [31:0] n24191;
wire     [31:0] n24192;
wire     [31:0] n24193;
wire     [31:0] n24194;
wire     [31:0] n24195;
wire     [31:0] n24196;
wire     [31:0] n24197;
wire     [31:0] n24198;
wire     [31:0] n24199;
wire     [31:0] n24200;
wire     [31:0] n24201;
wire     [31:0] n24202;
wire     [31:0] n24203;
wire     [31:0] n24204;
wire     [31:0] n24205;
wire     [31:0] n24206;
wire     [31:0] n24207;
wire     [31:0] n24208;
wire     [31:0] n24209;
wire     [31:0] n24210;
wire     [31:0] n24211;
wire     [31:0] n24212;
wire     [31:0] n24213;
wire     [31:0] n24214;
wire     [31:0] n24215;
wire     [31:0] n24216;
wire     [31:0] n24217;
wire     [31:0] n24218;
wire     [31:0] n24219;
wire     [31:0] n24220;
wire     [31:0] n24221;
wire     [31:0] n24222;
wire     [31:0] n24223;
wire            n24224;
wire            n24225;
wire     [31:0] n24226;
wire     [31:0] n24227;
wire     [31:0] n24228;
wire     [31:0] n24229;
wire     [31:0] n24230;
wire     [31:0] n24231;
wire     [31:0] n24232;
wire     [31:0] n24233;
wire     [31:0] n24234;
wire     [31:0] n24235;
wire     [31:0] n24236;
wire     [31:0] n24237;
wire     [31:0] n24238;
wire     [31:0] n24239;
wire     [31:0] n24240;
wire     [31:0] n24241;
wire     [31:0] n24242;
wire     [31:0] n24243;
wire     [31:0] n24244;
wire     [31:0] n24245;
wire     [31:0] n24246;
wire     [31:0] n24247;
wire     [31:0] n24248;
wire     [31:0] n24249;
wire     [31:0] n24250;
wire     [31:0] n24251;
wire     [31:0] n24252;
wire     [31:0] n24253;
wire     [31:0] n24254;
wire     [31:0] n24255;
wire     [31:0] n24256;
wire     [31:0] n24257;
wire     [31:0] n24258;
wire            n24259;
wire            n24260;
wire            n24261;
wire            n24262;
wire            n24263;
wire            n24264;
wire            n24265;
wire            n24266;
wire            n24267;
wire            n24268;
wire            n24269;
wire            n24270;
wire            n24271;
wire            n24272;
wire            n24273;
wire            n24274;
wire            n24275;
wire            n24276;
wire            n24277;
wire            n24278;
wire            n24279;
wire            n24280;
wire            n24281;
wire            n24282;
wire            n24283;
wire            n24284;
wire            n24285;
wire            n24286;
wire            n24287;
wire            n24288;
wire            n24289;
wire            n24290;
wire            n24291;
wire            n24292;
wire            n24293;
wire            n24294;
wire            n24295;
wire            n24296;
wire            n24297;
wire            n24298;
wire            n24299;
wire            n24300;
wire            n24301;
wire            n24302;
wire            n24303;
wire            n24304;
wire            n24305;
wire            n24306;
wire            n24307;
wire            n24308;
wire            n24309;
wire            n24310;
wire            n24311;
wire            n24312;
wire            n24313;
wire            n24314;
wire            n24315;
wire            n24316;
wire            n24317;
wire            n24318;
wire            n24319;
wire            n24320;
wire            n24321;
wire            n24322;
wire            n24323;
wire            n24324;
wire            n24325;
wire            n24326;
wire            n24327;
wire            n24328;
wire            n24329;
wire            n24330;
wire            n24331;
wire            n24332;
wire            n24333;
wire            n24334;
wire            n24335;
wire            n24336;
wire            n24337;
wire            n24338;
wire            n24339;
wire            n24340;
wire            n24341;
wire            n24342;
wire            n24343;
wire            n24344;
wire            n24345;
wire            n24346;
wire            n24347;
wire            n24348;
wire            n24349;
wire            n24350;
wire            n24351;
wire            n24352;
wire            n24353;
wire            n24354;
wire            n24355;
wire            n24356;
wire            n24357;
wire            n24358;
wire            n24359;
wire            n24360;
wire            n24361;
wire            n24362;
wire            n24363;
wire            n24364;
wire            n24365;
wire            n24366;
wire            n24367;
wire            n24368;
wire            n24369;
wire            n24370;
wire            n24371;
wire            n24372;
wire            n24373;
wire            n24374;
wire            n24375;
wire            n24376;
wire            n24377;
wire            n24378;
wire            n24379;
wire            n24380;
wire            n24381;
wire            n24382;
wire            n24383;
wire            n24384;
wire            n24385;
wire            n24386;
wire            n24387;
wire            n24388;
wire            n24389;
wire            n24390;
wire            n24391;
wire            n24392;
wire            n24393;
wire            n24394;
wire            n24395;
wire            n24396;
wire            n24397;
wire            n24398;
wire            n24399;
wire            n24400;
wire            n24401;
wire            n24402;
wire            n24403;
wire            n24404;
wire            n24405;
wire            n24406;
wire            n24407;
wire            n24408;
wire            n24409;
wire            n24410;
wire            n24411;
wire            n24412;
wire            n24413;
wire            n24414;
wire            n24415;
wire            n24416;
wire            n24417;
wire            n24418;
wire            n24419;
wire            n24420;
wire            n24421;
wire            n24422;
wire            n24423;
wire            n24424;
wire            n24425;
wire            n24426;
wire            n24427;
wire            n24428;
wire            n24429;
wire            n24430;
wire            n24431;
wire            n24432;
wire            n24433;
wire            n24434;
wire            n24435;
wire            n24436;
wire            n24437;
wire            n24438;
wire            n24439;
wire            n24440;
wire            n24441;
wire            n24442;
wire            n24443;
wire            n24444;
wire            n24445;
wire            n24446;
wire            n24447;
wire            n24448;
wire            n24449;
wire            n24450;
wire            n24451;
wire            n24452;
wire            n24453;
wire            n24454;
wire            n24455;
wire            n24456;
wire            n24457;
wire            n24458;
wire            n24459;
wire            n24460;
wire            n24461;
wire            n24462;
wire            n24463;
wire            n24464;
wire            n24465;
wire            n24466;
wire            n24467;
wire            n24468;
wire            n24469;
wire            n24470;
wire            n24471;
wire            n24472;
wire            n24473;
wire            n24474;
wire            n24475;
wire            n24476;
wire            n24477;
wire            n24478;
wire            n24479;
wire            n24480;
wire            n24481;
wire            n24482;
wire            n24483;
wire            n24484;
wire            n24485;
wire            n24486;
wire            n24487;
wire            n24488;
wire            n24489;
wire            n24490;
wire            n24491;
wire            n24492;
wire            n24493;
wire            n24494;
wire            n24495;
wire            n24496;
wire            n24497;
wire            n24498;
wire            n24499;
wire            n24500;
wire            n24501;
wire            n24502;
wire            n24503;
wire            n24504;
wire            n24505;
wire            n24506;
wire            n24507;
wire            n24508;
wire            n24509;
wire            n24510;
wire            n24511;
wire            n24512;
wire            n24513;
wire            n24514;
wire            n24515;
wire            n24516;
wire            n24517;
wire            n24518;
wire            n24519;
wire            n24520;
wire            n24521;
wire            n24522;
wire            n24523;
wire            n24524;
wire            n24525;
wire            n24526;
wire            n24527;
wire            n24528;
wire            n24529;
wire            n24530;
wire            n24531;
wire            n24532;
wire            n24533;
wire            n24534;
wire            n24535;
wire            n24536;
wire            n24537;
wire            n24538;
wire            n24539;
wire            n24540;
wire            n24541;
wire            n24542;
wire            n24543;
wire            n24544;
wire            n24545;
wire            n24546;
wire            n24547;
wire            n24548;
wire            n24549;
wire            n24550;
wire            n24551;
wire            n24552;
wire            n24553;
wire            n24554;
wire            n24555;
wire            n24556;
wire            n24557;
wire            n24558;
wire            n24559;
wire            n24560;
wire            n24561;
wire            n24562;
wire            n24563;
wire            n24564;
wire            n24565;
wire            n24566;
wire            n24567;
wire            n24568;
wire            n24569;
wire            n24570;
wire            n24571;
wire            n24572;
wire            n24573;
wire            n24574;
wire            n24575;
wire            n24576;
wire            n24577;
wire            n24578;
wire            n24579;
wire            n24580;
wire            n24581;
wire            n24582;
wire            n24583;
wire            n24584;
wire            n24585;
wire            n24586;
wire            n24587;
wire            n24588;
wire            n24589;
wire            n24590;
wire            n24591;
wire            n24592;
wire            n24593;
wire            n24594;
wire            n24595;
wire            n24596;
wire            n24597;
wire            n24598;
wire            n24599;
wire            n24600;
wire            n24601;
wire            n24602;
wire            n24603;
wire            n24604;
wire            n24605;
wire            n24606;
wire            n24607;
wire            n24608;
wire            n24609;
wire            n24610;
wire            n24611;
wire            n24612;
wire            n24613;
wire            n24614;
wire            n24615;
wire            n24616;
wire            n24617;
wire            n24618;
wire            n24619;
wire            n24620;
wire            n24621;
wire            n24622;
wire            n24623;
wire            n24624;
wire            n24625;
wire            n24626;
wire            n24627;
wire            n24628;
wire            n24629;
wire            n24630;
wire            n24631;
wire            n24632;
wire            n24633;
wire            n24634;
wire            n24635;
wire            n24636;
wire            n24637;
wire            n24638;
wire            n24639;
wire            n24640;
wire            n24641;
wire            n24642;
wire            n24643;
wire            n24644;
wire            n24645;
wire            n24646;
wire            n24647;
wire            n24648;
wire            n24649;
wire            n24650;
wire            n24651;
wire            n24652;
wire            n24653;
wire            n24654;
wire            n24655;
wire            n24656;
wire            n24657;
wire            n24658;
wire            n24659;
wire            n24660;
wire            n24661;
wire            n24662;
wire            n24663;
wire            n24664;
wire            n24665;
wire            n24666;
wire            n24667;
wire            n24668;
wire            n24669;
wire            n24670;
wire            n24671;
wire            n24672;
wire            n24673;
wire            n24674;
wire            n24675;
wire            n24676;
wire            n24677;
wire            n24678;
wire            n24679;
wire            n24680;
wire            n24681;
wire            n24682;
wire            n24683;
wire            n24684;
wire            n24685;
wire            n24686;
wire            n24687;
wire            n24688;
wire            n24689;
wire            n24690;
wire            n24691;
wire            n24692;
wire            n24693;
wire            n24694;
wire            n24695;
wire            n24696;
wire            n24697;
wire            n24698;
wire            n24699;
wire            n24700;
wire            n24701;
wire            n24702;
wire            n24703;
wire            n24704;
wire            n24705;
wire            n24706;
wire            n24707;
wire            n24708;
wire            n24709;
wire            n24710;
wire            n24711;
wire            n24712;
wire            n24713;
wire            n24714;
wire            n24715;
wire            n24716;
wire            n24717;
wire            n24718;
wire            n24719;
wire            n24720;
wire            n24721;
wire            n24722;
wire            n24723;
wire            n24724;
wire            n24725;
wire            n24726;
wire            n24727;
wire            n24728;
wire            n24729;
wire            n24730;
wire            n24731;
wire            n24732;
wire            n24733;
wire            n24734;
wire            n24735;
wire            n24736;
wire            n24737;
wire            n24738;
wire            n24739;
wire            n24740;
wire            n24741;
wire            n24742;
wire            n24743;
wire            n24744;
wire            n24745;
wire            n24746;
wire            n24747;
wire            n24748;
wire            n24749;
wire            n24750;
wire            n24751;
wire            n24752;
wire            n24753;
wire            n24754;
wire            n24755;
wire            n24756;
wire            n24757;
wire            n24758;
wire            n24759;
wire            n24760;
wire            n24761;
wire            n24762;
wire            n24763;
wire            n24764;
wire            n24765;
wire            n24766;
wire            n24767;
wire            n24768;
wire            n24769;
wire            n24770;
wire            n24771;
wire            n24772;
wire            n24773;
wire            n24774;
wire            n24775;
wire            n24776;
wire            n24777;
wire            n24778;
wire            n24779;
wire            n24780;
wire            n24781;
wire            n24782;
wire            n24783;
wire            n24784;
wire            n24785;
wire            n24786;
wire     [31:0] n24787;
wire     [31:0] n24788;
wire     [31:0] n24789;
wire     [31:0] n24790;
wire     [31:0] n24791;
wire     [31:0] n24792;
wire     [31:0] n24793;
wire     [31:0] n24794;
wire     [31:0] n24795;
wire     [31:0] n24796;
wire     [31:0] n24797;
wire     [31:0] n24798;
wire     [31:0] n24799;
wire     [31:0] n24800;
wire     [31:0] n24801;
wire     [31:0] n24802;
wire     [31:0] n24803;
wire     [31:0] n24804;
wire     [31:0] n24805;
wire     [31:0] n24806;
wire     [31:0] n24807;
wire     [31:0] n24808;
wire     [31:0] n24809;
wire     [31:0] n24810;
wire     [31:0] n24811;
wire     [31:0] n24812;
wire     [31:0] n24813;
wire     [31:0] n24814;
wire     [31:0] n24815;
wire     [31:0] n24816;
wire     [31:0] n24817;
wire     [31:0] n24818;
wire     [31:0] n24819;
wire     [31:0] n24820;
wire     [31:0] n24821;
wire     [31:0] n24822;
wire     [31:0] n24823;
wire     [31:0] n24824;
wire     [31:0] n24825;
wire     [31:0] n24826;
wire     [31:0] n24827;
wire     [31:0] n24828;
wire     [31:0] n24829;
wire     [31:0] n24830;
wire     [31:0] n24831;
wire     [31:0] n24832;
wire     [31:0] n24833;
wire     [31:0] n24834;
wire     [31:0] n24835;
wire     [31:0] n24836;
wire     [31:0] n24837;
wire     [31:0] n24838;
wire     [31:0] n24839;
wire     [31:0] n24840;
wire     [31:0] n24841;
wire     [31:0] n24842;
wire     [31:0] n24843;
wire     [31:0] n24844;
wire     [31:0] n24845;
wire     [31:0] n24846;
wire     [31:0] n24847;
wire     [31:0] n24848;
wire     [31:0] n24849;
wire     [31:0] n24850;
wire     [31:0] n24851;
wire     [31:0] n24852;
wire     [31:0] n24853;
wire     [31:0] n24854;
wire     [31:0] n24855;
wire     [31:0] n24856;
wire     [31:0] n24857;
wire     [31:0] n24858;
wire     [31:0] n24859;
wire     [31:0] n24860;
wire     [31:0] n24861;
wire     [31:0] n24862;
wire     [31:0] n24863;
wire     [31:0] n24864;
wire     [31:0] n24865;
wire     [31:0] n24866;
wire     [31:0] n24867;
wire     [31:0] n24868;
wire     [31:0] n24869;
wire     [31:0] n24870;
wire     [31:0] n24871;
wire     [31:0] n24872;
wire     [31:0] n24873;
wire     [31:0] n24874;
wire     [31:0] n24875;
wire     [31:0] n24876;
wire     [31:0] n24877;
wire     [31:0] n24878;
wire     [31:0] n24879;
wire     [31:0] n24880;
wire     [31:0] n24881;
wire     [31:0] n24882;
wire     [31:0] n24883;
wire     [31:0] n24884;
wire     [31:0] n24885;
wire     [31:0] n24886;
wire     [31:0] n24887;
wire     [31:0] n24888;
wire     [31:0] n24889;
wire     [31:0] n24890;
wire     [31:0] n24891;
wire     [31:0] n24892;
wire     [31:0] n24893;
wire     [31:0] n24894;
wire     [31:0] n24895;
wire     [31:0] n24896;
wire     [31:0] n24897;
wire     [31:0] n24898;
wire     [31:0] n24899;
wire     [31:0] n24900;
wire     [31:0] n24901;
wire     [31:0] n24902;
wire     [31:0] n24903;
wire     [31:0] n24904;
wire     [31:0] n24905;
wire     [31:0] n24906;
wire     [31:0] n24907;
wire     [31:0] n24908;
wire     [31:0] n24909;
wire     [31:0] n24910;
wire     [31:0] n24911;
wire     [31:0] n24912;
wire     [31:0] n24913;
wire     [31:0] n24914;
wire     [31:0] n24915;
wire     [31:0] n24916;
wire     [31:0] n24917;
wire     [31:0] n24918;
wire     [31:0] n24919;
wire     [31:0] n24920;
wire     [31:0] n24921;
wire     [31:0] n24922;
wire     [31:0] n24923;
wire     [31:0] n24924;
wire     [31:0] n24925;
wire     [31:0] n24926;
wire     [31:0] n24927;
wire     [31:0] n24928;
wire     [31:0] n24929;
wire     [31:0] n24930;
wire     [31:0] n24931;
wire     [31:0] n24932;
wire     [31:0] n24933;
wire     [31:0] n24934;
wire     [31:0] n24935;
wire     [31:0] n24936;
wire     [31:0] n24937;
wire     [31:0] n24938;
wire     [31:0] n24939;
wire     [31:0] n24940;
wire     [31:0] n24941;
wire     [31:0] n24942;
wire     [31:0] n24943;
wire     [31:0] n24944;
wire     [31:0] n24945;
wire     [31:0] n24946;
wire     [31:0] n24947;
wire     [31:0] n24948;
wire     [31:0] n24949;
wire     [31:0] n24950;
wire     [31:0] n24951;
wire     [31:0] n24952;
wire     [31:0] n24953;
wire     [31:0] n24954;
wire     [31:0] n24955;
wire     [31:0] n24956;
wire     [31:0] n24957;
wire     [31:0] n24958;
wire     [31:0] n24959;
wire     [31:0] n24960;
wire     [31:0] n24961;
wire     [31:0] n24962;
wire     [31:0] n24963;
wire     [31:0] n24964;
wire     [31:0] n24965;
wire     [31:0] n24966;
wire     [31:0] n24967;
wire     [31:0] n24968;
wire     [31:0] n24969;
wire     [31:0] n24970;
wire     [31:0] n24971;
wire     [31:0] n24972;
wire     [31:0] n24973;
wire     [31:0] n24974;
wire     [31:0] n24975;
wire     [31:0] n24976;
wire     [31:0] n24977;
wire     [31:0] n24978;
wire     [31:0] n24979;
wire     [31:0] n24980;
wire     [31:0] n24981;
wire     [31:0] n24982;
wire     [31:0] n24983;
wire     [31:0] n24984;
wire     [31:0] n24985;
wire     [31:0] n24986;
wire     [31:0] n24987;
wire     [31:0] n24988;
wire     [31:0] n24989;
wire     [31:0] n24990;
wire     [31:0] n24991;
wire     [31:0] n24992;
wire     [31:0] n24993;
wire     [31:0] n24994;
wire     [31:0] n24995;
wire     [31:0] n24996;
wire     [31:0] n24997;
wire     [31:0] n24998;
wire     [31:0] n24999;
wire     [31:0] n25000;
wire     [31:0] n25001;
wire     [31:0] n25002;
wire     [31:0] n25003;
wire     [31:0] n25004;
wire     [31:0] n25005;
wire     [31:0] n25006;
wire     [31:0] n25007;
wire     [31:0] n25008;
wire     [31:0] n25009;
wire     [31:0] n25010;
wire     [31:0] n25011;
wire     [31:0] n25012;
wire     [31:0] n25013;
wire     [31:0] n25014;
wire     [31:0] n25015;
wire     [31:0] n25016;
wire     [31:0] n25017;
wire     [31:0] n25018;
wire     [31:0] n25019;
wire     [31:0] n25020;
wire     [31:0] n25021;
wire     [31:0] n25022;
wire     [31:0] n25023;
wire     [31:0] n25024;
wire     [31:0] n25025;
wire     [31:0] n25026;
wire     [31:0] n25027;
wire     [31:0] n25028;
wire     [31:0] n25029;
wire     [31:0] n25030;
wire     [31:0] n25031;
wire     [31:0] n25032;
wire     [31:0] n25033;
wire     [31:0] n25034;
wire     [31:0] n25035;
wire     [31:0] n25036;
wire     [31:0] n25037;
wire     [31:0] n25038;
wire     [31:0] n25039;
wire     [31:0] n25040;
wire     [31:0] n25041;
wire     [31:0] n25042;
wire     [31:0] n25043;
wire     [31:0] n25044;
wire     [31:0] n25045;
wire     [31:0] n25046;
wire     [31:0] n25047;
wire     [31:0] n25048;
wire     [31:0] n25049;
wire     [31:0] n25050;
wire     [31:0] n25051;
wire     [31:0] n25052;
wire     [31:0] n25053;
wire     [31:0] n25054;
wire     [31:0] n25055;
wire     [31:0] n25056;
wire     [31:0] n25057;
wire     [31:0] n25058;
wire     [31:0] n25059;
wire     [31:0] n25060;
wire     [31:0] n25061;
wire     [31:0] n25062;
wire     [31:0] n25063;
wire     [31:0] n25064;
wire     [31:0] n25065;
wire     [31:0] n25066;
wire     [31:0] n25067;
wire     [31:0] n25068;
wire     [31:0] n25069;
wire     [31:0] n25070;
wire     [31:0] n25071;
wire     [31:0] n25072;
wire     [31:0] n25073;
wire     [31:0] n25074;
wire     [31:0] n25075;
wire     [31:0] n25076;
wire     [31:0] n25077;
wire     [31:0] n25078;
wire     [31:0] n25079;
wire     [31:0] n25080;
wire     [31:0] n25081;
wire     [31:0] n25082;
wire     [31:0] n25083;
wire     [31:0] n25084;
wire     [31:0] n25085;
wire     [31:0] n25086;
wire     [31:0] n25087;
wire     [31:0] n25088;
wire     [31:0] n25089;
wire     [31:0] n25090;
wire     [31:0] n25091;
wire     [31:0] n25092;
wire     [31:0] n25093;
wire     [31:0] n25094;
wire     [31:0] n25095;
wire     [31:0] n25096;
wire     [31:0] n25097;
wire     [31:0] n25098;
wire     [31:0] n25099;
wire     [31:0] n25100;
wire     [31:0] n25101;
wire     [31:0] n25102;
wire     [31:0] n25103;
wire     [31:0] n25104;
wire     [31:0] n25105;
wire     [31:0] n25106;
wire     [31:0] n25107;
wire     [31:0] n25108;
wire     [31:0] n25109;
wire     [31:0] n25110;
wire     [31:0] n25111;
wire     [31:0] n25112;
wire     [31:0] n25113;
wire     [31:0] n25114;
wire     [31:0] n25115;
wire     [31:0] n25116;
wire     [31:0] n25117;
wire     [31:0] n25118;
wire     [31:0] n25119;
wire     [31:0] n25120;
wire     [31:0] n25121;
wire     [31:0] n25122;
wire     [31:0] n25123;
wire     [31:0] n25124;
wire     [31:0] n25125;
wire     [31:0] n25126;
wire     [31:0] n25127;
wire     [31:0] n25128;
wire     [31:0] n25129;
wire     [31:0] n25130;
wire     [31:0] n25131;
wire     [31:0] n25132;
wire     [31:0] n25133;
wire     [31:0] n25134;
wire     [31:0] n25135;
wire     [31:0] n25136;
wire     [31:0] n25137;
wire     [31:0] n25138;
wire     [31:0] n25139;
wire     [31:0] n25140;
wire     [31:0] n25141;
wire     [31:0] n25142;
wire     [31:0] n25143;
wire     [31:0] n25144;
wire     [31:0] n25145;
wire     [31:0] n25146;
wire     [31:0] n25147;
wire     [31:0] n25148;
wire     [31:0] n25149;
wire     [31:0] n25150;
wire     [31:0] n25151;
wire     [31:0] n25152;
wire     [31:0] n25153;
wire     [31:0] n25154;
wire     [31:0] n25155;
wire     [31:0] n25156;
wire     [31:0] n25157;
wire     [31:0] n25158;
wire     [31:0] n25159;
wire     [31:0] n25160;
wire     [31:0] n25161;
wire     [31:0] n25162;
wire     [31:0] n25163;
wire     [31:0] n25164;
wire     [31:0] n25165;
wire     [31:0] n25166;
wire     [31:0] n25167;
wire     [31:0] n25168;
wire     [31:0] n25169;
wire     [31:0] n25170;
wire     [31:0] n25171;
wire     [31:0] n25172;
wire     [31:0] n25173;
wire     [31:0] n25174;
wire     [31:0] n25175;
wire     [31:0] n25176;
wire     [31:0] n25177;
wire     [31:0] n25178;
wire     [31:0] n25179;
wire     [31:0] n25180;
wire     [31:0] n25181;
wire     [31:0] n25182;
wire     [31:0] n25183;
wire     [31:0] n25184;
wire     [31:0] n25185;
wire     [31:0] n25186;
wire     [31:0] n25187;
wire     [31:0] n25188;
wire     [31:0] n25189;
wire     [31:0] n25190;
wire     [31:0] n25191;
wire     [31:0] n25192;
wire     [31:0] n25193;
wire     [31:0] n25194;
wire     [31:0] n25195;
wire     [31:0] n25196;
wire     [31:0] n25197;
wire     [31:0] n25198;
wire     [31:0] n25199;
wire     [31:0] n25200;
wire     [31:0] n25201;
wire     [31:0] n25202;
wire     [31:0] n25203;
wire     [31:0] n25204;
wire     [31:0] n25205;
wire     [31:0] n25206;
wire     [31:0] n25207;
wire     [31:0] n25208;
wire     [31:0] n25209;
wire     [31:0] n25210;
wire     [31:0] n25211;
wire     [31:0] n25212;
wire     [31:0] n25213;
wire     [31:0] n25214;
wire     [31:0] n25215;
wire     [31:0] n25216;
wire     [31:0] n25217;
wire     [31:0] n25218;
wire     [31:0] n25219;
wire     [31:0] n25220;
wire     [31:0] n25221;
wire     [31:0] n25222;
wire     [31:0] n25223;
wire     [31:0] n25224;
wire     [31:0] n25225;
wire     [31:0] n25226;
wire     [31:0] n25227;
wire     [31:0] n25228;
wire     [31:0] n25229;
wire     [31:0] n25230;
wire     [31:0] n25231;
wire     [31:0] n25232;
wire     [31:0] n25233;
wire     [31:0] n25234;
wire     [31:0] n25235;
wire     [31:0] n25236;
wire     [31:0] n25237;
wire     [31:0] n25238;
wire     [31:0] n25239;
wire     [31:0] n25240;
wire     [31:0] n25241;
wire     [31:0] n25242;
wire     [31:0] n25243;
wire     [31:0] n25244;
wire     [31:0] n25245;
wire     [31:0] n25246;
wire     [31:0] n25247;
wire     [31:0] n25248;
wire     [31:0] n25249;
wire     [31:0] n25250;
wire     [31:0] n25251;
wire     [31:0] n25252;
wire     [31:0] n25253;
wire     [31:0] n25254;
wire     [31:0] n25255;
wire     [31:0] n25256;
wire     [31:0] n25257;
wire     [31:0] n25258;
wire     [31:0] n25259;
wire     [31:0] n25260;
wire     [31:0] n25261;
wire     [31:0] n25262;
wire     [31:0] n25263;
wire     [31:0] n25264;
wire     [31:0] n25265;
wire     [31:0] n25266;
wire     [31:0] n25267;
wire     [31:0] n25268;
wire     [31:0] n25269;
wire     [31:0] n25270;
wire     [31:0] n25271;
wire     [31:0] n25272;
wire     [31:0] n25273;
wire     [31:0] n25274;
wire     [31:0] n25275;
wire     [31:0] n25276;
wire     [31:0] n25277;
wire     [31:0] n25278;
wire     [31:0] n25279;
wire     [31:0] n25280;
wire     [31:0] n25281;
wire     [31:0] n25282;
wire     [31:0] n25283;
wire     [31:0] n25284;
wire     [31:0] n25285;
wire     [31:0] n25286;
wire     [31:0] n25287;
wire     [31:0] n25288;
wire     [31:0] n25289;
wire     [31:0] n25290;
wire     [31:0] n25291;
wire     [31:0] n25292;
wire     [31:0] n25293;
wire     [31:0] n25294;
wire     [31:0] n25295;
wire     [31:0] n25296;
wire     [31:0] n25297;
wire     [31:0] n25298;
wire     [31:0] n25299;
wire     [31:0] n25300;
wire     [31:0] n25301;
wire     [31:0] n25302;
wire     [31:0] n25303;
wire     [31:0] n25304;
wire     [31:0] n25305;
wire     [31:0] n25306;
wire     [31:0] n25307;
wire     [31:0] n25308;
wire            n25309;
wire            n25310;
wire            n25311;
wire            n25312;
wire            n25313;
wire            n25314;
wire            n25315;
wire            n25316;
wire            n25317;
wire            n25318;
wire            n25319;
wire            n25320;
wire            n25321;
wire            n25322;
wire            n25323;
wire            n25324;
wire            n25325;
wire            n25326;
wire            n25327;
wire            n25328;
wire            n25329;
wire            n25330;
wire            n25331;
wire            n25332;
wire            n25333;
wire            n25334;
wire            n25335;
wire            n25336;
wire            n25337;
wire            n25338;
wire            n25339;
wire            n25340;
wire            n25341;
wire            n25342;
wire            n25343;
wire            n25344;
wire            n25345;
wire            n25346;
wire            n25347;
wire            n25348;
wire            n25349;
wire            n25350;
wire            n25351;
wire            n25352;
wire            n25353;
wire            n25354;
wire            n25355;
wire            n25356;
wire            n25357;
wire            n25358;
wire            n25359;
wire            n25360;
wire            n25361;
wire            n25362;
wire            n25363;
wire            n25364;
wire            n25365;
wire            n25366;
wire            n25367;
wire            n25368;
wire            n25369;
wire            n25370;
wire            n25371;
wire            n25372;
wire            n25373;
wire            n25374;
wire            n25375;
wire            n25376;
wire            n25377;
wire            n25378;
wire            n25379;
wire            n25380;
wire            n25381;
wire            n25382;
wire            n25383;
wire            n25384;
wire            n25385;
wire            n25386;
wire            n25387;
wire            n25388;
wire            n25389;
wire            n25390;
wire            n25391;
wire            n25392;
wire            n25393;
wire            n25394;
wire            n25395;
wire            n25396;
wire            n25397;
wire            n25398;
wire            n25399;
wire            n25400;
wire            n25401;
wire            n25402;
wire            n25403;
wire            n25404;
wire            n25405;
wire            n25406;
wire            n25407;
wire            n25408;
wire            n25409;
wire            n25410;
wire            n25411;
wire            n25412;
wire            n25413;
wire            n25414;
wire            n25415;
wire            n25416;
wire            n25417;
wire            n25418;
wire            n25419;
wire            n25420;
wire            n25421;
wire            n25422;
wire            n25423;
wire            n25424;
wire            n25425;
wire            n25426;
wire            n25427;
wire            n25428;
wire            n25429;
wire            n25430;
wire            n25431;
wire            n25432;
wire            n25433;
wire            n25434;
wire            n25435;
wire            n25436;
wire            n25437;
wire            n25438;
wire            n25439;
wire            n25440;
wire            n25441;
wire            n25442;
wire            n25443;
wire            n25444;
wire            n25445;
wire            n25446;
wire            n25447;
wire            n25448;
wire            n25449;
wire            n25450;
wire            n25451;
wire            n25452;
wire            n25453;
wire            n25454;
wire            n25455;
wire            n25456;
wire            n25457;
wire            n25458;
wire            n25459;
wire            n25460;
wire            n25461;
wire            n25462;
wire            n25463;
wire            n25464;
wire            n25465;
wire            n25466;
wire            n25467;
wire            n25468;
wire            n25469;
wire            n25470;
wire            n25471;
wire            n25472;
wire            n25473;
wire            n25474;
wire            n25475;
wire            n25476;
wire            n25477;
wire            n25478;
wire            n25479;
wire            n25480;
wire            n25481;
wire            n25482;
wire            n25483;
wire            n25484;
wire            n25485;
wire            n25486;
wire            n25487;
wire            n25488;
wire            n25489;
wire            n25490;
wire            n25491;
wire            n25492;
wire            n25493;
wire            n25494;
wire            n25495;
wire            n25496;
wire            n25497;
wire            n25498;
wire            n25499;
wire            n25500;
wire            n25501;
wire            n25502;
wire            n25503;
wire            n25504;
wire            n25505;
wire            n25506;
wire            n25507;
wire            n25508;
wire            n25509;
wire            n25510;
wire            n25511;
wire            n25512;
wire            n25513;
wire            n25514;
wire            n25515;
wire            n25516;
wire            n25517;
wire            n25518;
wire            n25519;
wire            n25520;
wire            n25521;
wire            n25522;
wire            n25523;
wire            n25524;
wire            n25525;
wire            n25526;
wire            n25527;
wire            n25528;
wire            n25529;
wire            n25530;
wire            n25531;
wire            n25532;
wire            n25533;
wire            n25534;
wire            n25535;
wire            n25536;
wire            n25537;
wire            n25538;
wire            n25539;
wire            n25540;
wire            n25541;
wire            n25542;
wire            n25543;
wire            n25544;
wire            n25545;
wire            n25546;
wire            n25547;
wire            n25548;
wire            n25549;
wire            n25550;
wire            n25551;
wire            n25552;
wire            n25553;
wire            n25554;
wire            n25555;
wire            n25556;
wire            n25557;
wire            n25558;
wire            n25559;
wire            n25560;
wire            n25561;
wire            n25562;
wire            n25563;
wire            n25564;
wire            n25565;
wire            n25566;
wire            n25567;
wire            n25568;
wire            n25569;
wire            n25570;
wire            n25571;
wire            n25572;
wire            n25573;
wire            n25574;
wire            n25575;
wire            n25576;
wire            n25577;
wire            n25578;
wire            n25579;
wire            n25580;
wire            n25581;
wire            n25582;
wire            n25583;
wire            n25584;
wire            n25585;
wire            n25586;
wire            n25587;
wire            n25588;
wire            n25589;
wire            n25590;
wire            n25591;
wire            n25592;
wire            n25593;
wire            n25594;
wire            n25595;
wire            n25596;
wire            n25597;
wire            n25598;
wire            n25599;
wire            n25600;
wire            n25601;
wire            n25602;
wire            n25603;
wire            n25604;
wire            n25605;
wire            n25606;
wire            n25607;
wire            n25608;
wire            n25609;
wire            n25610;
wire            n25611;
wire            n25612;
wire            n25613;
wire            n25614;
wire            n25615;
wire            n25616;
wire            n25617;
wire            n25618;
wire            n25619;
wire            n25620;
wire            n25621;
wire            n25622;
wire            n25623;
wire            n25624;
wire            n25625;
wire            n25626;
wire            n25627;
wire            n25628;
wire            n25629;
wire            n25630;
wire            n25631;
wire            n25632;
wire            n25633;
wire            n25634;
wire            n25635;
wire            n25636;
wire            n25637;
wire            n25638;
wire            n25639;
wire            n25640;
wire            n25641;
wire            n25642;
wire            n25643;
wire            n25644;
wire            n25645;
wire            n25646;
wire            n25647;
wire            n25648;
wire            n25649;
wire            n25650;
wire            n25651;
wire            n25652;
wire            n25653;
wire            n25654;
wire            n25655;
wire            n25656;
wire            n25657;
wire            n25658;
wire            n25659;
wire            n25660;
wire            n25661;
wire            n25662;
wire            n25663;
wire            n25664;
wire            n25665;
wire            n25666;
wire            n25667;
wire            n25668;
wire            n25669;
wire            n25670;
wire            n25671;
wire            n25672;
wire            n25673;
wire            n25674;
wire            n25675;
wire            n25676;
wire            n25677;
wire            n25678;
wire            n25679;
wire            n25680;
wire            n25681;
wire            n25682;
wire            n25683;
wire            n25684;
wire            n25685;
wire            n25686;
wire            n25687;
wire            n25688;
wire            n25689;
wire            n25690;
wire            n25691;
wire            n25692;
wire            n25693;
wire            n25694;
wire            n25695;
wire            n25696;
wire            n25697;
wire            n25698;
wire            n25699;
wire            n25700;
wire            n25701;
wire            n25702;
wire            n25703;
wire            n25704;
wire            n25705;
wire            n25706;
wire            n25707;
wire            n25708;
wire            n25709;
wire            n25710;
wire            n25711;
wire            n25712;
wire            n25713;
wire            n25714;
wire            n25715;
wire            n25716;
wire            n25717;
wire            n25718;
wire            n25719;
wire            n25720;
wire            n25721;
wire            n25722;
wire            n25723;
wire            n25724;
wire            n25725;
wire            n25726;
wire            n25727;
wire            n25728;
wire            n25729;
wire            n25730;
wire            n25731;
wire            n25732;
wire            n25733;
wire            n25734;
wire            n25735;
wire            n25736;
wire            n25737;
wire            n25738;
wire            n25739;
wire            n25740;
wire            n25741;
wire            n25742;
wire            n25743;
wire            n25744;
wire            n25745;
wire            n25746;
wire            n25747;
wire            n25748;
wire            n25749;
wire            n25750;
wire            n25751;
wire            n25752;
wire            n25753;
wire            n25754;
wire            n25755;
wire            n25756;
wire            n25757;
wire            n25758;
wire            n25759;
wire            n25760;
wire            n25761;
wire            n25762;
wire            n25763;
wire            n25764;
wire            n25765;
wire            n25766;
wire            n25767;
wire            n25768;
wire            n25769;
wire            n25770;
wire            n25771;
wire            n25772;
wire            n25773;
wire            n25774;
wire            n25775;
wire            n25776;
wire            n25777;
wire            n25778;
wire            n25779;
wire            n25780;
wire            n25781;
wire            n25782;
wire            n25783;
wire            n25784;
wire            n25785;
wire            n25786;
wire            n25787;
wire            n25788;
wire            n25789;
wire            n25790;
wire            n25791;
wire            n25792;
wire            n25793;
wire            n25794;
wire            n25795;
wire            n25796;
wire            n25797;
wire            n25798;
wire            n25799;
wire            n25800;
wire            n25801;
wire            n25802;
wire            n25803;
wire            n25804;
wire            n25805;
wire            n25806;
wire            n25807;
wire            n25808;
wire            n25809;
wire            n25810;
wire            n25811;
wire            n25812;
wire            n25813;
wire            n25814;
wire            n25815;
wire            n25816;
wire            n25817;
wire            n25818;
wire            n25819;
wire            n25820;
wire     [31:0] n25821;
wire     [31:0] n25822;
wire     [31:0] n25823;
wire     [31:0] n25824;
wire     [31:0] n25825;
wire     [31:0] n25826;
wire     [31:0] n25827;
wire     [31:0] n25828;
wire     [31:0] n25829;
wire     [31:0] n25830;
wire     [31:0] n25831;
wire     [31:0] n25832;
wire     [31:0] n25833;
wire     [31:0] n25834;
wire     [31:0] n25835;
wire     [31:0] n25836;
wire     [31:0] n25837;
wire     [31:0] n25838;
wire     [31:0] n25839;
wire     [31:0] n25840;
wire     [31:0] n25841;
wire     [31:0] n25842;
wire     [31:0] n25843;
wire     [31:0] n25844;
wire     [31:0] n25845;
wire     [31:0] n25846;
wire     [31:0] n25847;
wire     [31:0] n25848;
wire     [31:0] n25849;
wire     [31:0] n25850;
wire     [31:0] n25851;
wire     [31:0] n25852;
wire     [31:0] n25853;
wire     [31:0] n25854;
wire     [31:0] n25855;
wire     [31:0] n25856;
wire     [31:0] n25857;
wire     [31:0] n25858;
wire     [31:0] n25859;
wire     [31:0] n25860;
wire     [31:0] n25861;
wire     [31:0] n25862;
wire     [31:0] n25863;
wire     [31:0] n25864;
wire     [31:0] n25865;
wire     [31:0] n25866;
wire     [31:0] n25867;
wire     [31:0] n25868;
wire     [31:0] n25869;
wire     [31:0] n25870;
wire     [31:0] n25871;
wire     [31:0] n25872;
wire     [31:0] n25873;
wire     [31:0] n25874;
wire     [31:0] n25875;
wire     [31:0] n25876;
wire     [31:0] n25877;
wire     [31:0] n25878;
wire     [31:0] n25879;
wire     [31:0] n25880;
wire     [31:0] n25881;
wire     [31:0] n25882;
wire     [31:0] n25883;
wire     [31:0] n25884;
wire     [31:0] n25885;
wire     [31:0] n25886;
wire     [31:0] n25887;
wire     [31:0] n25888;
wire     [31:0] n25889;
wire     [31:0] n25890;
wire     [31:0] n25891;
wire     [31:0] n25892;
wire     [31:0] n25893;
wire     [31:0] n25894;
wire     [31:0] n25895;
wire     [31:0] n25896;
wire     [31:0] n25897;
wire     [31:0] n25898;
wire     [31:0] n25899;
wire     [31:0] n25900;
wire     [31:0] n25901;
wire     [31:0] n25902;
wire     [31:0] n25903;
wire     [31:0] n25904;
wire     [31:0] n25905;
wire     [31:0] n25906;
wire     [31:0] n25907;
wire     [31:0] n25908;
wire     [31:0] n25909;
wire     [31:0] n25910;
wire     [31:0] n25911;
wire     [31:0] n25912;
wire     [31:0] n25913;
wire     [31:0] n25914;
wire     [31:0] n25915;
wire     [31:0] n25916;
wire     [31:0] n25917;
wire     [31:0] n25918;
wire     [31:0] n25919;
wire     [31:0] n25920;
wire     [31:0] n25921;
wire     [31:0] n25922;
wire     [31:0] n25923;
wire     [31:0] n25924;
wire     [31:0] n25925;
wire     [31:0] n25926;
wire     [31:0] n25927;
wire     [31:0] n25928;
wire     [31:0] n25929;
wire     [31:0] n25930;
wire     [31:0] n25931;
wire     [31:0] n25932;
wire     [31:0] n25933;
wire     [31:0] n25934;
wire     [31:0] n25935;
wire     [31:0] n25936;
wire     [31:0] n25937;
wire     [31:0] n25938;
wire     [31:0] n25939;
wire     [31:0] n25940;
wire     [31:0] n25941;
wire     [31:0] n25942;
wire     [31:0] n25943;
wire     [31:0] n25944;
wire     [31:0] n25945;
wire     [31:0] n25946;
wire     [31:0] n25947;
wire     [31:0] n25948;
wire     [31:0] n25949;
wire     [31:0] n25950;
wire     [31:0] n25951;
wire     [31:0] n25952;
wire     [31:0] n25953;
wire     [31:0] n25954;
wire     [31:0] n25955;
wire     [31:0] n25956;
wire     [31:0] n25957;
wire     [31:0] n25958;
wire     [31:0] n25959;
wire     [31:0] n25960;
wire     [31:0] n25961;
wire     [31:0] n25962;
wire     [31:0] n25963;
wire     [31:0] n25964;
wire     [31:0] n25965;
wire     [31:0] n25966;
wire     [31:0] n25967;
wire     [31:0] n25968;
wire     [31:0] n25969;
wire     [31:0] n25970;
wire     [31:0] n25971;
wire     [31:0] n25972;
wire     [31:0] n25973;
wire     [31:0] n25974;
wire     [31:0] n25975;
wire     [31:0] n25976;
wire     [31:0] n25977;
wire     [31:0] n25978;
wire     [31:0] n25979;
wire     [31:0] n25980;
wire     [31:0] n25981;
wire     [31:0] n25982;
wire     [31:0] n25983;
wire     [31:0] n25984;
wire     [31:0] n25985;
wire     [31:0] n25986;
wire     [31:0] n25987;
wire     [31:0] n25988;
wire     [31:0] n25989;
wire     [31:0] n25990;
wire     [31:0] n25991;
wire     [31:0] n25992;
wire     [31:0] n25993;
wire     [31:0] n25994;
wire     [31:0] n25995;
wire     [31:0] n25996;
wire     [31:0] n25997;
wire     [31:0] n25998;
wire     [31:0] n25999;
wire     [31:0] n26000;
wire     [31:0] n26001;
wire     [31:0] n26002;
wire     [31:0] n26003;
wire     [31:0] n26004;
wire     [31:0] n26005;
wire     [31:0] n26006;
wire     [31:0] n26007;
wire     [31:0] n26008;
wire     [31:0] n26009;
wire     [31:0] n26010;
wire     [31:0] n26011;
wire     [31:0] n26012;
wire     [31:0] n26013;
wire     [31:0] n26014;
wire     [31:0] n26015;
wire     [31:0] n26016;
wire     [31:0] n26017;
wire     [31:0] n26018;
wire     [31:0] n26019;
wire     [31:0] n26020;
wire     [31:0] n26021;
wire     [31:0] n26022;
wire     [31:0] n26023;
wire     [31:0] n26024;
wire     [31:0] n26025;
wire     [31:0] n26026;
wire     [31:0] n26027;
wire     [31:0] n26028;
wire     [31:0] n26029;
wire     [31:0] n26030;
wire     [31:0] n26031;
wire     [31:0] n26032;
wire     [31:0] n26033;
wire     [31:0] n26034;
wire     [31:0] n26035;
wire     [31:0] n26036;
wire     [31:0] n26037;
wire     [31:0] n26038;
wire     [31:0] n26039;
wire     [31:0] n26040;
wire     [31:0] n26041;
wire     [31:0] n26042;
wire     [31:0] n26043;
wire     [31:0] n26044;
wire     [31:0] n26045;
wire     [31:0] n26046;
wire     [31:0] n26047;
wire     [31:0] n26048;
wire     [31:0] n26049;
wire     [31:0] n26050;
wire     [31:0] n26051;
wire     [31:0] n26052;
wire     [31:0] n26053;
wire     [31:0] n26054;
wire     [31:0] n26055;
wire     [31:0] n26056;
wire     [31:0] n26057;
wire     [31:0] n26058;
wire     [31:0] n26059;
wire     [31:0] n26060;
wire     [31:0] n26061;
wire     [31:0] n26062;
wire     [31:0] n26063;
wire     [31:0] n26064;
wire     [31:0] n26065;
wire     [31:0] n26066;
wire     [31:0] n26067;
wire     [31:0] n26068;
wire     [31:0] n26069;
wire     [31:0] n26070;
wire     [31:0] n26071;
wire     [31:0] n26072;
wire     [31:0] n26073;
wire     [31:0] n26074;
wire     [31:0] n26075;
wire     [31:0] n26076;
wire     [31:0] n26077;
wire     [31:0] n26078;
wire     [31:0] n26079;
wire     [31:0] n26080;
wire     [31:0] n26081;
wire     [31:0] n26082;
wire     [31:0] n26083;
wire     [31:0] n26084;
wire     [31:0] n26085;
wire     [31:0] n26086;
wire     [31:0] n26087;
wire     [31:0] n26088;
wire     [31:0] n26089;
wire     [31:0] n26090;
wire     [31:0] n26091;
wire     [31:0] n26092;
wire     [31:0] n26093;
wire     [31:0] n26094;
wire     [31:0] n26095;
wire     [31:0] n26096;
wire     [31:0] n26097;
wire     [31:0] n26098;
wire     [31:0] n26099;
wire     [31:0] n26100;
wire     [31:0] n26101;
wire     [31:0] n26102;
wire     [31:0] n26103;
wire     [31:0] n26104;
wire     [31:0] n26105;
wire     [31:0] n26106;
wire     [31:0] n26107;
wire     [31:0] n26108;
wire     [31:0] n26109;
wire     [31:0] n26110;
wire     [31:0] n26111;
wire     [31:0] n26112;
wire     [31:0] n26113;
wire     [31:0] n26114;
wire     [31:0] n26115;
wire     [31:0] n26116;
wire     [31:0] n26117;
wire     [31:0] n26118;
wire     [31:0] n26119;
wire     [31:0] n26120;
wire     [31:0] n26121;
wire     [31:0] n26122;
wire     [31:0] n26123;
wire     [31:0] n26124;
wire     [31:0] n26125;
wire     [31:0] n26126;
wire     [31:0] n26127;
wire     [31:0] n26128;
wire     [31:0] n26129;
wire     [31:0] n26130;
wire     [31:0] n26131;
wire     [31:0] n26132;
wire     [31:0] n26133;
wire     [31:0] n26134;
wire     [31:0] n26135;
wire     [31:0] n26136;
wire     [31:0] n26137;
wire     [31:0] n26138;
wire     [31:0] n26139;
wire     [31:0] n26140;
wire     [31:0] n26141;
wire     [31:0] n26142;
wire     [31:0] n26143;
wire     [31:0] n26144;
wire     [31:0] n26145;
wire     [31:0] n26146;
wire     [31:0] n26147;
wire     [31:0] n26148;
wire     [31:0] n26149;
wire     [31:0] n26150;
wire     [31:0] n26151;
wire     [31:0] n26152;
wire     [31:0] n26153;
wire     [31:0] n26154;
wire     [31:0] n26155;
wire     [31:0] n26156;
wire     [31:0] n26157;
wire     [31:0] n26158;
wire     [31:0] n26159;
wire     [31:0] n26160;
wire     [31:0] n26161;
wire     [31:0] n26162;
wire     [31:0] n26163;
wire     [31:0] n26164;
wire     [31:0] n26165;
wire     [31:0] n26166;
wire     [31:0] n26167;
wire     [31:0] n26168;
wire     [31:0] n26169;
wire     [31:0] n26170;
wire     [31:0] n26171;
wire     [31:0] n26172;
wire     [31:0] n26173;
wire     [31:0] n26174;
wire     [31:0] n26175;
wire     [31:0] n26176;
wire     [31:0] n26177;
wire     [31:0] n26178;
wire     [31:0] n26179;
wire     [31:0] n26180;
wire     [31:0] n26181;
wire     [31:0] n26182;
wire     [31:0] n26183;
wire     [31:0] n26184;
wire     [31:0] n26185;
wire     [31:0] n26186;
wire     [31:0] n26187;
wire     [31:0] n26188;
wire     [31:0] n26189;
wire     [31:0] n26190;
wire     [31:0] n26191;
wire     [31:0] n26192;
wire     [31:0] n26193;
wire     [31:0] n26194;
wire     [31:0] n26195;
wire     [31:0] n26196;
wire     [31:0] n26197;
wire     [31:0] n26198;
wire     [31:0] n26199;
wire     [31:0] n26200;
wire     [31:0] n26201;
wire     [31:0] n26202;
wire     [31:0] n26203;
wire     [31:0] n26204;
wire     [31:0] n26205;
wire     [31:0] n26206;
wire     [31:0] n26207;
wire     [31:0] n26208;
wire     [31:0] n26209;
wire     [31:0] n26210;
wire     [31:0] n26211;
wire     [31:0] n26212;
wire     [31:0] n26213;
wire     [31:0] n26214;
wire     [31:0] n26215;
wire     [31:0] n26216;
wire     [31:0] n26217;
wire     [31:0] n26218;
wire     [31:0] n26219;
wire     [31:0] n26220;
wire     [31:0] n26221;
wire     [31:0] n26222;
wire     [31:0] n26223;
wire     [31:0] n26224;
wire     [31:0] n26225;
wire     [31:0] n26226;
wire     [31:0] n26227;
wire     [31:0] n26228;
wire     [31:0] n26229;
wire     [31:0] n26230;
wire     [31:0] n26231;
wire     [31:0] n26232;
wire     [31:0] n26233;
wire     [31:0] n26234;
wire     [31:0] n26235;
wire     [31:0] n26236;
wire     [31:0] n26237;
wire     [31:0] n26238;
wire     [31:0] n26239;
wire     [31:0] n26240;
wire     [31:0] n26241;
wire     [31:0] n26242;
wire     [31:0] n26243;
wire     [31:0] n26244;
wire     [31:0] n26245;
wire     [31:0] n26246;
wire     [31:0] n26247;
wire     [31:0] n26248;
wire     [31:0] n26249;
wire     [31:0] n26250;
wire     [31:0] n26251;
wire     [31:0] n26252;
wire     [31:0] n26253;
wire     [31:0] n26254;
wire     [31:0] n26255;
wire     [31:0] n26256;
wire     [31:0] n26257;
wire     [31:0] n26258;
wire     [31:0] n26259;
wire     [31:0] n26260;
wire     [31:0] n26261;
wire     [31:0] n26262;
wire     [31:0] n26263;
wire     [31:0] n26264;
wire     [31:0] n26265;
wire     [31:0] n26266;
wire     [31:0] n26267;
wire     [31:0] n26268;
wire     [31:0] n26269;
wire     [31:0] n26270;
wire     [31:0] n26271;
wire     [31:0] n26272;
wire     [31:0] n26273;
wire     [31:0] n26274;
wire     [31:0] n26275;
wire     [31:0] n26276;
wire     [31:0] n26277;
wire     [31:0] n26278;
wire     [31:0] n26279;
wire     [31:0] n26280;
wire     [31:0] n26281;
wire     [31:0] n26282;
wire     [31:0] n26283;
wire     [31:0] n26284;
wire     [31:0] n26285;
wire     [31:0] n26286;
wire     [31:0] n26287;
wire     [31:0] n26288;
wire     [31:0] n26289;
wire     [31:0] n26290;
wire     [31:0] n26291;
wire     [31:0] n26292;
wire     [31:0] n26293;
wire     [31:0] n26294;
wire     [31:0] n26295;
wire     [31:0] n26296;
wire     [31:0] n26297;
wire     [31:0] n26298;
wire     [31:0] n26299;
wire     [31:0] n26300;
wire     [31:0] n26301;
wire     [31:0] n26302;
wire     [31:0] n26303;
wire     [31:0] n26304;
wire     [31:0] n26305;
wire     [31:0] n26306;
wire     [31:0] n26307;
wire     [31:0] n26308;
wire     [31:0] n26309;
wire     [31:0] n26310;
wire     [31:0] n26311;
wire     [31:0] n26312;
wire     [31:0] n26313;
wire     [31:0] n26314;
wire     [31:0] n26315;
wire     [31:0] n26316;
wire     [31:0] n26317;
wire     [31:0] n26318;
wire     [31:0] n26319;
wire     [31:0] n26320;
wire     [31:0] n26321;
wire     [31:0] n26322;
wire     [31:0] n26323;
wire     [31:0] n26324;
wire     [31:0] n26325;
wire     [31:0] n26326;
wire     [31:0] n26327;
wire     [31:0] n26328;
wire     [31:0] n26329;
wire     [31:0] n26330;
wire     [31:0] n26331;
wire     [31:0] n26332;
wire     [31:0] n26333;
wire     [31:0] n26334;
wire     [31:0] n26335;
wire     [31:0] n26336;
wire     [31:0] n26337;
wire     [31:0] n26338;
wire     [31:0] n26339;
wire     [31:0] n26340;
wire     [31:0] n26341;
wire     [31:0] n26342;
wire            n26343;
wire            n26344;
wire     [31:0] n26345;
wire     [31:0] n26346;
wire     [31:0] n26347;
wire     [31:0] n26348;
wire     [31:0] n26349;
wire     [31:0] n26350;
wire     [31:0] n26351;
wire     [31:0] n26352;
wire     [31:0] n26353;
wire     [31:0] n26354;
wire     [31:0] n26355;
wire     [31:0] n26356;
wire     [31:0] n26357;
wire     [31:0] n26358;
wire     [31:0] n26359;
wire     [31:0] n26360;
wire     [31:0] n26361;
wire     [31:0] n26362;
wire     [31:0] n26363;
wire     [31:0] n26364;
wire     [31:0] n26365;
wire     [31:0] n26366;
wire     [31:0] n26367;
wire     [31:0] n26368;
wire     [31:0] n26369;
wire     [31:0] n26370;
wire     [31:0] n26371;
wire     [31:0] n26372;
wire     [31:0] n26373;
wire     [31:0] n26374;
wire     [31:0] n26375;
wire     [31:0] n26376;
wire     [31:0] n26377;
wire            n26378;
wire            n26379;
wire            n26380;
wire            n26381;
wire            n26382;
wire            n26383;
wire            n26384;
wire            n26385;
wire            n26386;
wire            n26387;
wire            n26388;
wire            n26389;
wire            n26390;
wire            n26391;
wire            n26392;
wire            n26393;
wire            n26394;
wire            n26395;
wire            n26396;
wire            n26397;
wire            n26398;
wire            n26399;
wire            n26400;
wire            n26401;
wire            n26402;
wire            n26403;
wire            n26404;
wire            n26405;
wire            n26406;
wire            n26407;
wire            n26408;
wire            n26409;
wire            n26410;
wire            n26411;
wire            n26412;
wire            n26413;
wire            n26414;
wire            n26415;
wire            n26416;
wire            n26417;
wire            n26418;
wire            n26419;
wire            n26420;
wire            n26421;
wire            n26422;
wire            n26423;
wire            n26424;
wire            n26425;
wire            n26426;
wire            n26427;
wire            n26428;
wire            n26429;
wire            n26430;
wire            n26431;
wire            n26432;
wire            n26433;
wire            n26434;
wire            n26435;
wire            n26436;
wire            n26437;
wire            n26438;
wire            n26439;
wire            n26440;
wire            n26441;
wire            n26442;
wire            n26443;
wire            n26444;
wire            n26445;
wire            n26446;
wire            n26447;
wire            n26448;
wire            n26449;
wire            n26450;
wire            n26451;
wire            n26452;
wire            n26453;
wire            n26454;
wire            n26455;
wire            n26456;
wire            n26457;
wire            n26458;
wire            n26459;
wire            n26460;
wire            n26461;
wire            n26462;
wire            n26463;
wire            n26464;
wire            n26465;
wire            n26466;
wire            n26467;
wire            n26468;
wire            n26469;
wire            n26470;
wire            n26471;
wire            n26472;
wire            n26473;
wire            n26474;
wire            n26475;
wire            n26476;
wire            n26477;
wire            n26478;
wire            n26479;
wire            n26480;
wire            n26481;
wire            n26482;
wire            n26483;
wire            n26484;
wire            n26485;
wire            n26486;
wire            n26487;
wire            n26488;
wire            n26489;
wire            n26490;
wire            n26491;
wire            n26492;
wire            n26493;
wire            n26494;
wire            n26495;
wire            n26496;
wire            n26497;
wire            n26498;
wire            n26499;
wire            n26500;
wire            n26501;
wire            n26502;
wire            n26503;
wire            n26504;
wire            n26505;
wire            n26506;
wire            n26507;
wire            n26508;
wire            n26509;
wire            n26510;
wire            n26511;
wire            n26512;
wire            n26513;
wire            n26514;
wire            n26515;
wire            n26516;
wire            n26517;
wire            n26518;
wire            n26519;
wire            n26520;
wire            n26521;
wire            n26522;
wire            n26523;
wire            n26524;
wire            n26525;
wire            n26526;
wire            n26527;
wire            n26528;
wire            n26529;
wire            n26530;
wire            n26531;
wire            n26532;
wire            n26533;
wire            n26534;
wire            n26535;
wire            n26536;
wire            n26537;
wire            n26538;
wire            n26539;
wire            n26540;
wire            n26541;
wire            n26542;
wire            n26543;
wire            n26544;
wire            n26545;
wire            n26546;
wire            n26547;
wire            n26548;
wire            n26549;
wire            n26550;
wire            n26551;
wire            n26552;
wire            n26553;
wire            n26554;
wire            n26555;
wire            n26556;
wire            n26557;
wire            n26558;
wire            n26559;
wire            n26560;
wire            n26561;
wire            n26562;
wire            n26563;
wire            n26564;
wire            n26565;
wire            n26566;
wire            n26567;
wire            n26568;
wire            n26569;
wire            n26570;
wire            n26571;
wire            n26572;
wire            n26573;
wire            n26574;
wire            n26575;
wire            n26576;
wire            n26577;
wire            n26578;
wire            n26579;
wire            n26580;
wire            n26581;
wire            n26582;
wire            n26583;
wire            n26584;
wire            n26585;
wire            n26586;
wire            n26587;
wire            n26588;
wire            n26589;
wire            n26590;
wire            n26591;
wire            n26592;
wire            n26593;
wire            n26594;
wire            n26595;
wire            n26596;
wire            n26597;
wire            n26598;
wire            n26599;
wire            n26600;
wire            n26601;
wire            n26602;
wire            n26603;
wire            n26604;
wire            n26605;
wire            n26606;
wire            n26607;
wire            n26608;
wire            n26609;
wire            n26610;
wire            n26611;
wire            n26612;
wire            n26613;
wire            n26614;
wire            n26615;
wire            n26616;
wire            n26617;
wire            n26618;
wire            n26619;
wire            n26620;
wire            n26621;
wire            n26622;
wire            n26623;
wire            n26624;
wire            n26625;
wire            n26626;
wire            n26627;
wire            n26628;
wire            n26629;
wire            n26630;
wire            n26631;
wire            n26632;
wire            n26633;
wire            n26634;
wire            n26635;
wire            n26636;
wire            n26637;
wire            n26638;
wire            n26639;
wire            n26640;
wire            n26641;
wire            n26642;
wire            n26643;
wire            n26644;
wire            n26645;
wire            n26646;
wire            n26647;
wire            n26648;
wire            n26649;
wire            n26650;
wire            n26651;
wire            n26652;
wire            n26653;
wire            n26654;
wire            n26655;
wire            n26656;
wire            n26657;
wire            n26658;
wire            n26659;
wire            n26660;
wire            n26661;
wire            n26662;
wire            n26663;
wire            n26664;
wire            n26665;
wire            n26666;
wire            n26667;
wire            n26668;
wire            n26669;
wire            n26670;
wire            n26671;
wire            n26672;
wire            n26673;
wire            n26674;
wire            n26675;
wire            n26676;
wire            n26677;
wire            n26678;
wire            n26679;
wire            n26680;
wire            n26681;
wire            n26682;
wire            n26683;
wire            n26684;
wire            n26685;
wire            n26686;
wire            n26687;
wire            n26688;
wire            n26689;
wire            n26690;
wire            n26691;
wire            n26692;
wire            n26693;
wire            n26694;
wire            n26695;
wire            n26696;
wire            n26697;
wire            n26698;
wire            n26699;
wire            n26700;
wire            n26701;
wire            n26702;
wire            n26703;
wire            n26704;
wire            n26705;
wire            n26706;
wire            n26707;
wire            n26708;
wire            n26709;
wire            n26710;
wire            n26711;
wire            n26712;
wire            n26713;
wire            n26714;
wire            n26715;
wire            n26716;
wire            n26717;
wire            n26718;
wire            n26719;
wire            n26720;
wire            n26721;
wire            n26722;
wire            n26723;
wire            n26724;
wire            n26725;
wire            n26726;
wire            n26727;
wire            n26728;
wire            n26729;
wire            n26730;
wire            n26731;
wire            n26732;
wire            n26733;
wire            n26734;
wire            n26735;
wire            n26736;
wire            n26737;
wire            n26738;
wire            n26739;
wire            n26740;
wire            n26741;
wire            n26742;
wire            n26743;
wire            n26744;
wire            n26745;
wire            n26746;
wire            n26747;
wire            n26748;
wire            n26749;
wire            n26750;
wire            n26751;
wire            n26752;
wire            n26753;
wire            n26754;
wire            n26755;
wire            n26756;
wire            n26757;
wire            n26758;
wire            n26759;
wire            n26760;
wire            n26761;
wire            n26762;
wire            n26763;
wire            n26764;
wire            n26765;
wire            n26766;
wire            n26767;
wire            n26768;
wire            n26769;
wire            n26770;
wire            n26771;
wire            n26772;
wire            n26773;
wire            n26774;
wire            n26775;
wire            n26776;
wire            n26777;
wire            n26778;
wire            n26779;
wire            n26780;
wire            n26781;
wire            n26782;
wire            n26783;
wire            n26784;
wire            n26785;
wire            n26786;
wire            n26787;
wire            n26788;
wire            n26789;
wire            n26790;
wire            n26791;
wire            n26792;
wire            n26793;
wire            n26794;
wire            n26795;
wire            n26796;
wire            n26797;
wire            n26798;
wire            n26799;
wire            n26800;
wire            n26801;
wire            n26802;
wire            n26803;
wire            n26804;
wire            n26805;
wire            n26806;
wire            n26807;
wire            n26808;
wire            n26809;
wire            n26810;
wire            n26811;
wire            n26812;
wire            n26813;
wire            n26814;
wire            n26815;
wire            n26816;
wire            n26817;
wire            n26818;
wire            n26819;
wire            n26820;
wire            n26821;
wire            n26822;
wire            n26823;
wire            n26824;
wire            n26825;
wire            n26826;
wire            n26827;
wire            n26828;
wire            n26829;
wire            n26830;
wire            n26831;
wire            n26832;
wire            n26833;
wire            n26834;
wire            n26835;
wire            n26836;
wire            n26837;
wire            n26838;
wire            n26839;
wire            n26840;
wire            n26841;
wire            n26842;
wire            n26843;
wire            n26844;
wire            n26845;
wire            n26846;
wire            n26847;
wire            n26848;
wire            n26849;
wire            n26850;
wire            n26851;
wire            n26852;
wire            n26853;
wire            n26854;
wire            n26855;
wire            n26856;
wire            n26857;
wire            n26858;
wire            n26859;
wire            n26860;
wire            n26861;
wire            n26862;
wire            n26863;
wire            n26864;
wire            n26865;
wire            n26866;
wire            n26867;
wire            n26868;
wire            n26869;
wire            n26870;
wire            n26871;
wire            n26872;
wire            n26873;
wire            n26874;
wire            n26875;
wire            n26876;
wire            n26877;
wire            n26878;
wire            n26879;
wire            n26880;
wire            n26881;
wire            n26882;
wire            n26883;
wire            n26884;
wire            n26885;
wire            n26886;
wire            n26887;
wire            n26888;
wire            n26889;
wire            n26890;
wire            n26891;
wire            n26892;
wire            n26893;
wire            n26894;
wire            n26895;
wire            n26896;
wire            n26897;
wire            n26898;
wire            n26899;
wire            n26900;
wire            n26901;
wire            n26902;
wire            n26903;
wire            n26904;
wire            n26905;
wire     [31:0] n26906;
wire     [31:0] n26907;
wire     [31:0] n26908;
wire     [31:0] n26909;
wire     [31:0] n26910;
wire     [31:0] n26911;
wire     [31:0] n26912;
wire     [31:0] n26913;
wire     [31:0] n26914;
wire     [31:0] n26915;
wire     [31:0] n26916;
wire     [31:0] n26917;
wire     [31:0] n26918;
wire     [31:0] n26919;
wire     [31:0] n26920;
wire     [31:0] n26921;
wire     [31:0] n26922;
wire     [31:0] n26923;
wire     [31:0] n26924;
wire     [31:0] n26925;
wire     [31:0] n26926;
wire     [31:0] n26927;
wire     [31:0] n26928;
wire     [31:0] n26929;
wire     [31:0] n26930;
wire     [31:0] n26931;
wire     [31:0] n26932;
wire     [31:0] n26933;
wire     [31:0] n26934;
wire     [31:0] n26935;
wire     [31:0] n26936;
wire     [31:0] n26937;
wire     [31:0] n26938;
wire     [31:0] n26939;
wire     [31:0] n26940;
wire     [31:0] n26941;
wire     [31:0] n26942;
wire     [31:0] n26943;
wire     [31:0] n26944;
wire     [31:0] n26945;
wire     [31:0] n26946;
wire     [31:0] n26947;
wire     [31:0] n26948;
wire     [31:0] n26949;
wire     [31:0] n26950;
wire     [31:0] n26951;
wire     [31:0] n26952;
wire     [31:0] n26953;
wire     [31:0] n26954;
wire     [31:0] n26955;
wire     [31:0] n26956;
wire     [31:0] n26957;
wire     [31:0] n26958;
wire     [31:0] n26959;
wire     [31:0] n26960;
wire     [31:0] n26961;
wire     [31:0] n26962;
wire     [31:0] n26963;
wire     [31:0] n26964;
wire     [31:0] n26965;
wire     [31:0] n26966;
wire     [31:0] n26967;
wire     [31:0] n26968;
wire     [31:0] n26969;
wire     [31:0] n26970;
wire     [31:0] n26971;
wire     [31:0] n26972;
wire     [31:0] n26973;
wire     [31:0] n26974;
wire     [31:0] n26975;
wire     [31:0] n26976;
wire     [31:0] n26977;
wire     [31:0] n26978;
wire     [31:0] n26979;
wire     [31:0] n26980;
wire     [31:0] n26981;
wire     [31:0] n26982;
wire     [31:0] n26983;
wire     [31:0] n26984;
wire     [31:0] n26985;
wire     [31:0] n26986;
wire     [31:0] n26987;
wire     [31:0] n26988;
wire     [31:0] n26989;
wire     [31:0] n26990;
wire     [31:0] n26991;
wire     [31:0] n26992;
wire     [31:0] n26993;
wire     [31:0] n26994;
wire     [31:0] n26995;
wire     [31:0] n26996;
wire     [31:0] n26997;
wire     [31:0] n26998;
wire     [31:0] n26999;
wire     [31:0] n27000;
wire     [31:0] n27001;
wire     [31:0] n27002;
wire     [31:0] n27003;
wire     [31:0] n27004;
wire     [31:0] n27005;
wire     [31:0] n27006;
wire     [31:0] n27007;
wire     [31:0] n27008;
wire     [31:0] n27009;
wire     [31:0] n27010;
wire     [31:0] n27011;
wire     [31:0] n27012;
wire     [31:0] n27013;
wire     [31:0] n27014;
wire     [31:0] n27015;
wire     [31:0] n27016;
wire     [31:0] n27017;
wire     [31:0] n27018;
wire     [31:0] n27019;
wire     [31:0] n27020;
wire     [31:0] n27021;
wire     [31:0] n27022;
wire     [31:0] n27023;
wire     [31:0] n27024;
wire     [31:0] n27025;
wire     [31:0] n27026;
wire     [31:0] n27027;
wire     [31:0] n27028;
wire     [31:0] n27029;
wire     [31:0] n27030;
wire     [31:0] n27031;
wire     [31:0] n27032;
wire     [31:0] n27033;
wire     [31:0] n27034;
wire     [31:0] n27035;
wire     [31:0] n27036;
wire     [31:0] n27037;
wire     [31:0] n27038;
wire     [31:0] n27039;
wire     [31:0] n27040;
wire     [31:0] n27041;
wire     [31:0] n27042;
wire     [31:0] n27043;
wire     [31:0] n27044;
wire     [31:0] n27045;
wire     [31:0] n27046;
wire     [31:0] n27047;
wire     [31:0] n27048;
wire     [31:0] n27049;
wire     [31:0] n27050;
wire     [31:0] n27051;
wire     [31:0] n27052;
wire     [31:0] n27053;
wire     [31:0] n27054;
wire     [31:0] n27055;
wire     [31:0] n27056;
wire     [31:0] n27057;
wire     [31:0] n27058;
wire     [31:0] n27059;
wire     [31:0] n27060;
wire     [31:0] n27061;
wire     [31:0] n27062;
wire     [31:0] n27063;
wire     [31:0] n27064;
wire     [31:0] n27065;
wire     [31:0] n27066;
wire     [31:0] n27067;
wire     [31:0] n27068;
wire     [31:0] n27069;
wire     [31:0] n27070;
wire     [31:0] n27071;
wire     [31:0] n27072;
wire     [31:0] n27073;
wire     [31:0] n27074;
wire     [31:0] n27075;
wire     [31:0] n27076;
wire     [31:0] n27077;
wire     [31:0] n27078;
wire     [31:0] n27079;
wire     [31:0] n27080;
wire     [31:0] n27081;
wire     [31:0] n27082;
wire     [31:0] n27083;
wire     [31:0] n27084;
wire     [31:0] n27085;
wire     [31:0] n27086;
wire     [31:0] n27087;
wire     [31:0] n27088;
wire     [31:0] n27089;
wire     [31:0] n27090;
wire     [31:0] n27091;
wire     [31:0] n27092;
wire     [31:0] n27093;
wire     [31:0] n27094;
wire     [31:0] n27095;
wire     [31:0] n27096;
wire     [31:0] n27097;
wire     [31:0] n27098;
wire     [31:0] n27099;
wire     [31:0] n27100;
wire     [31:0] n27101;
wire     [31:0] n27102;
wire     [31:0] n27103;
wire     [31:0] n27104;
wire     [31:0] n27105;
wire     [31:0] n27106;
wire     [31:0] n27107;
wire     [31:0] n27108;
wire     [31:0] n27109;
wire     [31:0] n27110;
wire     [31:0] n27111;
wire     [31:0] n27112;
wire     [31:0] n27113;
wire     [31:0] n27114;
wire     [31:0] n27115;
wire     [31:0] n27116;
wire     [31:0] n27117;
wire     [31:0] n27118;
wire     [31:0] n27119;
wire     [31:0] n27120;
wire     [31:0] n27121;
wire     [31:0] n27122;
wire     [31:0] n27123;
wire     [31:0] n27124;
wire     [31:0] n27125;
wire     [31:0] n27126;
wire     [31:0] n27127;
wire     [31:0] n27128;
wire     [31:0] n27129;
wire     [31:0] n27130;
wire     [31:0] n27131;
wire     [31:0] n27132;
wire     [31:0] n27133;
wire     [31:0] n27134;
wire     [31:0] n27135;
wire     [31:0] n27136;
wire     [31:0] n27137;
wire     [31:0] n27138;
wire     [31:0] n27139;
wire     [31:0] n27140;
wire     [31:0] n27141;
wire     [31:0] n27142;
wire     [31:0] n27143;
wire     [31:0] n27144;
wire     [31:0] n27145;
wire     [31:0] n27146;
wire     [31:0] n27147;
wire     [31:0] n27148;
wire     [31:0] n27149;
wire     [31:0] n27150;
wire     [31:0] n27151;
wire     [31:0] n27152;
wire     [31:0] n27153;
wire     [31:0] n27154;
wire     [31:0] n27155;
wire     [31:0] n27156;
wire     [31:0] n27157;
wire     [31:0] n27158;
wire     [31:0] n27159;
wire     [31:0] n27160;
wire     [31:0] n27161;
wire     [31:0] n27162;
wire     [31:0] n27163;
wire     [31:0] n27164;
wire     [31:0] n27165;
wire     [31:0] n27166;
wire     [31:0] n27167;
wire     [31:0] n27168;
wire     [31:0] n27169;
wire     [31:0] n27170;
wire     [31:0] n27171;
wire     [31:0] n27172;
wire     [31:0] n27173;
wire     [31:0] n27174;
wire     [31:0] n27175;
wire     [31:0] n27176;
wire     [31:0] n27177;
wire     [31:0] n27178;
wire     [31:0] n27179;
wire     [31:0] n27180;
wire     [31:0] n27181;
wire     [31:0] n27182;
wire     [31:0] n27183;
wire     [31:0] n27184;
wire     [31:0] n27185;
wire     [31:0] n27186;
wire     [31:0] n27187;
wire     [31:0] n27188;
wire     [31:0] n27189;
wire     [31:0] n27190;
wire     [31:0] n27191;
wire     [31:0] n27192;
wire     [31:0] n27193;
wire     [31:0] n27194;
wire     [31:0] n27195;
wire     [31:0] n27196;
wire     [31:0] n27197;
wire     [31:0] n27198;
wire     [31:0] n27199;
wire     [31:0] n27200;
wire     [31:0] n27201;
wire     [31:0] n27202;
wire     [31:0] n27203;
wire     [31:0] n27204;
wire     [31:0] n27205;
wire     [31:0] n27206;
wire     [31:0] n27207;
wire     [31:0] n27208;
wire     [31:0] n27209;
wire     [31:0] n27210;
wire     [31:0] n27211;
wire     [31:0] n27212;
wire     [31:0] n27213;
wire     [31:0] n27214;
wire     [31:0] n27215;
wire     [31:0] n27216;
wire     [31:0] n27217;
wire     [31:0] n27218;
wire     [31:0] n27219;
wire     [31:0] n27220;
wire     [31:0] n27221;
wire     [31:0] n27222;
wire     [31:0] n27223;
wire     [31:0] n27224;
wire     [31:0] n27225;
wire     [31:0] n27226;
wire     [31:0] n27227;
wire     [31:0] n27228;
wire     [31:0] n27229;
wire     [31:0] n27230;
wire     [31:0] n27231;
wire     [31:0] n27232;
wire     [31:0] n27233;
wire     [31:0] n27234;
wire     [31:0] n27235;
wire     [31:0] n27236;
wire     [31:0] n27237;
wire     [31:0] n27238;
wire     [31:0] n27239;
wire     [31:0] n27240;
wire     [31:0] n27241;
wire     [31:0] n27242;
wire     [31:0] n27243;
wire     [31:0] n27244;
wire     [31:0] n27245;
wire     [31:0] n27246;
wire     [31:0] n27247;
wire     [31:0] n27248;
wire     [31:0] n27249;
wire     [31:0] n27250;
wire     [31:0] n27251;
wire     [31:0] n27252;
wire     [31:0] n27253;
wire     [31:0] n27254;
wire     [31:0] n27255;
wire     [31:0] n27256;
wire     [31:0] n27257;
wire     [31:0] n27258;
wire     [31:0] n27259;
wire     [31:0] n27260;
wire     [31:0] n27261;
wire     [31:0] n27262;
wire     [31:0] n27263;
wire     [31:0] n27264;
wire     [31:0] n27265;
wire     [31:0] n27266;
wire     [31:0] n27267;
wire     [31:0] n27268;
wire     [31:0] n27269;
wire     [31:0] n27270;
wire     [31:0] n27271;
wire     [31:0] n27272;
wire     [31:0] n27273;
wire     [31:0] n27274;
wire     [31:0] n27275;
wire     [31:0] n27276;
wire     [31:0] n27277;
wire     [31:0] n27278;
wire     [31:0] n27279;
wire     [31:0] n27280;
wire     [31:0] n27281;
wire     [31:0] n27282;
wire     [31:0] n27283;
wire     [31:0] n27284;
wire     [31:0] n27285;
wire     [31:0] n27286;
wire     [31:0] n27287;
wire     [31:0] n27288;
wire     [31:0] n27289;
wire     [31:0] n27290;
wire     [31:0] n27291;
wire     [31:0] n27292;
wire     [31:0] n27293;
wire     [31:0] n27294;
wire     [31:0] n27295;
wire     [31:0] n27296;
wire     [31:0] n27297;
wire     [31:0] n27298;
wire     [31:0] n27299;
wire     [31:0] n27300;
wire     [31:0] n27301;
wire     [31:0] n27302;
wire     [31:0] n27303;
wire     [31:0] n27304;
wire     [31:0] n27305;
wire     [31:0] n27306;
wire     [31:0] n27307;
wire     [31:0] n27308;
wire     [31:0] n27309;
wire     [31:0] n27310;
wire     [31:0] n27311;
wire     [31:0] n27312;
wire     [31:0] n27313;
wire     [31:0] n27314;
wire     [31:0] n27315;
wire     [31:0] n27316;
wire     [31:0] n27317;
wire     [31:0] n27318;
wire     [31:0] n27319;
wire     [31:0] n27320;
wire     [31:0] n27321;
wire     [31:0] n27322;
wire     [31:0] n27323;
wire     [31:0] n27324;
wire     [31:0] n27325;
wire     [31:0] n27326;
wire     [31:0] n27327;
wire     [31:0] n27328;
wire     [31:0] n27329;
wire     [31:0] n27330;
wire     [31:0] n27331;
wire     [31:0] n27332;
wire     [31:0] n27333;
wire     [31:0] n27334;
wire     [31:0] n27335;
wire     [31:0] n27336;
wire     [31:0] n27337;
wire     [31:0] n27338;
wire     [31:0] n27339;
wire     [31:0] n27340;
wire     [31:0] n27341;
wire     [31:0] n27342;
wire     [31:0] n27343;
wire     [31:0] n27344;
wire     [31:0] n27345;
wire     [31:0] n27346;
wire     [31:0] n27347;
wire     [31:0] n27348;
wire     [31:0] n27349;
wire     [31:0] n27350;
wire     [31:0] n27351;
wire     [31:0] n27352;
wire     [31:0] n27353;
wire     [31:0] n27354;
wire     [31:0] n27355;
wire     [31:0] n27356;
wire     [31:0] n27357;
wire     [31:0] n27358;
wire     [31:0] n27359;
wire     [31:0] n27360;
wire     [31:0] n27361;
wire     [31:0] n27362;
wire     [31:0] n27363;
wire     [31:0] n27364;
wire     [31:0] n27365;
wire     [31:0] n27366;
wire     [31:0] n27367;
wire     [31:0] n27368;
wire     [31:0] n27369;
wire     [31:0] n27370;
wire     [31:0] n27371;
wire     [31:0] n27372;
wire     [31:0] n27373;
wire     [31:0] n27374;
wire     [31:0] n27375;
wire     [31:0] n27376;
wire     [31:0] n27377;
wire     [31:0] n27378;
wire     [31:0] n27379;
wire     [31:0] n27380;
wire     [31:0] n27381;
wire     [31:0] n27382;
wire     [31:0] n27383;
wire     [31:0] n27384;
wire     [31:0] n27385;
wire     [31:0] n27386;
wire     [31:0] n27387;
wire     [31:0] n27388;
wire     [31:0] n27389;
wire     [31:0] n27390;
wire     [31:0] n27391;
wire     [31:0] n27392;
wire     [31:0] n27393;
wire     [31:0] n27394;
wire     [31:0] n27395;
wire     [31:0] n27396;
wire     [31:0] n27397;
wire     [31:0] n27398;
wire     [31:0] n27399;
wire     [31:0] n27400;
wire     [31:0] n27401;
wire     [31:0] n27402;
wire     [31:0] n27403;
wire     [31:0] n27404;
wire     [31:0] n27405;
wire     [31:0] n27406;
wire     [31:0] n27407;
wire     [31:0] n27408;
wire     [31:0] n27409;
wire     [31:0] n27410;
wire     [31:0] n27411;
wire     [31:0] n27412;
wire     [31:0] n27413;
wire     [31:0] n27414;
wire     [31:0] n27415;
wire     [31:0] n27416;
wire     [31:0] n27417;
wire     [31:0] n27418;
wire     [31:0] n27419;
wire     [31:0] n27420;
wire     [31:0] n27421;
wire     [31:0] n27422;
wire     [31:0] n27423;
wire     [31:0] n27424;
wire     [31:0] n27425;
wire     [31:0] n27426;
wire     [31:0] n27427;
wire            n27428;
wire            n27429;
wire            n27430;
wire            n27431;
wire            n27432;
wire            n27433;
wire            n27434;
wire            n27435;
wire            n27436;
wire            n27437;
wire            n27438;
wire            n27439;
wire            n27440;
wire            n27441;
wire            n27442;
wire            n27443;
wire            n27444;
wire            n27445;
wire            n27446;
wire            n27447;
wire            n27448;
wire            n27449;
wire            n27450;
wire            n27451;
wire            n27452;
wire            n27453;
wire            n27454;
wire            n27455;
wire            n27456;
wire            n27457;
wire            n27458;
wire            n27459;
wire            n27460;
wire            n27461;
wire            n27462;
wire            n27463;
wire            n27464;
wire            n27465;
wire            n27466;
wire            n27467;
wire            n27468;
wire            n27469;
wire            n27470;
wire            n27471;
wire            n27472;
wire            n27473;
wire            n27474;
wire            n27475;
wire            n27476;
wire            n27477;
wire            n27478;
wire            n27479;
wire            n27480;
wire            n27481;
wire            n27482;
wire            n27483;
wire            n27484;
wire            n27485;
wire            n27486;
wire            n27487;
wire            n27488;
wire            n27489;
wire            n27490;
wire            n27491;
wire            n27492;
wire            n27493;
wire            n27494;
wire            n27495;
wire            n27496;
wire            n27497;
wire            n27498;
wire            n27499;
wire            n27500;
wire            n27501;
wire            n27502;
wire            n27503;
wire            n27504;
wire            n27505;
wire            n27506;
wire            n27507;
wire            n27508;
wire            n27509;
wire            n27510;
wire            n27511;
wire            n27512;
wire            n27513;
wire            n27514;
wire            n27515;
wire            n27516;
wire            n27517;
wire            n27518;
wire            n27519;
wire            n27520;
wire            n27521;
wire            n27522;
wire            n27523;
wire            n27524;
wire            n27525;
wire            n27526;
wire            n27527;
wire            n27528;
wire            n27529;
wire            n27530;
wire            n27531;
wire            n27532;
wire            n27533;
wire            n27534;
wire            n27535;
wire            n27536;
wire            n27537;
wire            n27538;
wire            n27539;
wire            n27540;
wire            n27541;
wire            n27542;
wire            n27543;
wire            n27544;
wire            n27545;
wire            n27546;
wire            n27547;
wire            n27548;
wire            n27549;
wire            n27550;
wire            n27551;
wire            n27552;
wire            n27553;
wire            n27554;
wire            n27555;
wire            n27556;
wire            n27557;
wire            n27558;
wire            n27559;
wire            n27560;
wire            n27561;
wire            n27562;
wire            n27563;
wire            n27564;
wire            n27565;
wire            n27566;
wire            n27567;
wire            n27568;
wire            n27569;
wire            n27570;
wire            n27571;
wire            n27572;
wire            n27573;
wire            n27574;
wire            n27575;
wire            n27576;
wire            n27577;
wire            n27578;
wire            n27579;
wire            n27580;
wire            n27581;
wire            n27582;
wire            n27583;
wire            n27584;
wire            n27585;
wire            n27586;
wire            n27587;
wire            n27588;
wire            n27589;
wire            n27590;
wire            n27591;
wire            n27592;
wire            n27593;
wire            n27594;
wire            n27595;
wire            n27596;
wire            n27597;
wire            n27598;
wire            n27599;
wire            n27600;
wire            n27601;
wire            n27602;
wire            n27603;
wire            n27604;
wire            n27605;
wire            n27606;
wire            n27607;
wire            n27608;
wire            n27609;
wire            n27610;
wire            n27611;
wire            n27612;
wire            n27613;
wire            n27614;
wire            n27615;
wire            n27616;
wire            n27617;
wire            n27618;
wire            n27619;
wire            n27620;
wire            n27621;
wire            n27622;
wire            n27623;
wire            n27624;
wire            n27625;
wire            n27626;
wire            n27627;
wire            n27628;
wire            n27629;
wire            n27630;
wire            n27631;
wire            n27632;
wire            n27633;
wire            n27634;
wire            n27635;
wire            n27636;
wire            n27637;
wire            n27638;
wire            n27639;
wire            n27640;
wire            n27641;
wire            n27642;
wire            n27643;
wire            n27644;
wire            n27645;
wire            n27646;
wire            n27647;
wire            n27648;
wire            n27649;
wire            n27650;
wire            n27651;
wire            n27652;
wire            n27653;
wire            n27654;
wire            n27655;
wire            n27656;
wire            n27657;
wire            n27658;
wire            n27659;
wire            n27660;
wire            n27661;
wire            n27662;
wire            n27663;
wire            n27664;
wire            n27665;
wire            n27666;
wire            n27667;
wire            n27668;
wire            n27669;
wire            n27670;
wire            n27671;
wire            n27672;
wire            n27673;
wire            n27674;
wire            n27675;
wire            n27676;
wire            n27677;
wire            n27678;
wire            n27679;
wire            n27680;
wire            n27681;
wire            n27682;
wire            n27683;
wire            n27684;
wire            n27685;
wire            n27686;
wire            n27687;
wire            n27688;
wire            n27689;
wire            n27690;
wire            n27691;
wire            n27692;
wire            n27693;
wire            n27694;
wire            n27695;
wire            n27696;
wire            n27697;
wire            n27698;
wire            n27699;
wire            n27700;
wire            n27701;
wire            n27702;
wire            n27703;
wire            n27704;
wire            n27705;
wire            n27706;
wire            n27707;
wire            n27708;
wire            n27709;
wire            n27710;
wire            n27711;
wire            n27712;
wire            n27713;
wire            n27714;
wire            n27715;
wire            n27716;
wire            n27717;
wire            n27718;
wire            n27719;
wire            n27720;
wire            n27721;
wire            n27722;
wire            n27723;
wire            n27724;
wire            n27725;
wire            n27726;
wire            n27727;
wire            n27728;
wire            n27729;
wire            n27730;
wire            n27731;
wire            n27732;
wire            n27733;
wire            n27734;
wire            n27735;
wire            n27736;
wire            n27737;
wire            n27738;
wire            n27739;
wire            n27740;
wire            n27741;
wire            n27742;
wire            n27743;
wire            n27744;
wire            n27745;
wire            n27746;
wire            n27747;
wire            n27748;
wire            n27749;
wire            n27750;
wire            n27751;
wire            n27752;
wire            n27753;
wire            n27754;
wire            n27755;
wire            n27756;
wire            n27757;
wire            n27758;
wire            n27759;
wire            n27760;
wire            n27761;
wire            n27762;
wire            n27763;
wire            n27764;
wire            n27765;
wire            n27766;
wire            n27767;
wire            n27768;
wire            n27769;
wire            n27770;
wire            n27771;
wire            n27772;
wire            n27773;
wire            n27774;
wire            n27775;
wire            n27776;
wire            n27777;
wire            n27778;
wire            n27779;
wire            n27780;
wire            n27781;
wire            n27782;
wire            n27783;
wire            n27784;
wire            n27785;
wire            n27786;
wire            n27787;
wire            n27788;
wire            n27789;
wire            n27790;
wire            n27791;
wire            n27792;
wire            n27793;
wire            n27794;
wire            n27795;
wire            n27796;
wire            n27797;
wire            n27798;
wire            n27799;
wire            n27800;
wire            n27801;
wire            n27802;
wire            n27803;
wire            n27804;
wire            n27805;
wire            n27806;
wire            n27807;
wire            n27808;
wire            n27809;
wire            n27810;
wire            n27811;
wire            n27812;
wire            n27813;
wire            n27814;
wire            n27815;
wire            n27816;
wire            n27817;
wire            n27818;
wire            n27819;
wire            n27820;
wire            n27821;
wire            n27822;
wire            n27823;
wire            n27824;
wire            n27825;
wire            n27826;
wire            n27827;
wire            n27828;
wire            n27829;
wire            n27830;
wire            n27831;
wire            n27832;
wire            n27833;
wire            n27834;
wire            n27835;
wire            n27836;
wire            n27837;
wire            n27838;
wire            n27839;
wire            n27840;
wire            n27841;
wire            n27842;
wire            n27843;
wire            n27844;
wire            n27845;
wire            n27846;
wire            n27847;
wire            n27848;
wire            n27849;
wire            n27850;
wire            n27851;
wire            n27852;
wire            n27853;
wire            n27854;
wire            n27855;
wire            n27856;
wire            n27857;
wire            n27858;
wire            n27859;
wire            n27860;
wire            n27861;
wire            n27862;
wire            n27863;
wire            n27864;
wire            n27865;
wire            n27866;
wire            n27867;
wire            n27868;
wire            n27869;
wire            n27870;
wire            n27871;
wire            n27872;
wire            n27873;
wire            n27874;
wire            n27875;
wire            n27876;
wire            n27877;
wire            n27878;
wire            n27879;
wire            n27880;
wire            n27881;
wire            n27882;
wire            n27883;
wire            n27884;
wire            n27885;
wire            n27886;
wire            n27887;
wire            n27888;
wire            n27889;
wire            n27890;
wire            n27891;
wire            n27892;
wire            n27893;
wire            n27894;
wire            n27895;
wire            n27896;
wire            n27897;
wire            n27898;
wire            n27899;
wire            n27900;
wire            n27901;
wire            n27902;
wire            n27903;
wire            n27904;
wire            n27905;
wire            n27906;
wire            n27907;
wire            n27908;
wire            n27909;
wire            n27910;
wire            n27911;
wire            n27912;
wire            n27913;
wire            n27914;
wire            n27915;
wire            n27916;
wire            n27917;
wire            n27918;
wire            n27919;
wire            n27920;
wire            n27921;
wire            n27922;
wire            n27923;
wire            n27924;
wire            n27925;
wire            n27926;
wire            n27927;
wire            n27928;
wire            n27929;
wire            n27930;
wire            n27931;
wire            n27932;
wire            n27933;
wire            n27934;
wire            n27935;
wire            n27936;
wire            n27937;
wire            n27938;
wire            n27939;
wire     [31:0] n27940;
wire     [31:0] n27941;
wire     [31:0] n27942;
wire     [31:0] n27943;
wire     [31:0] n27944;
wire     [31:0] n27945;
wire     [31:0] n27946;
wire     [31:0] n27947;
wire     [31:0] n27948;
wire     [31:0] n27949;
wire     [31:0] n27950;
wire     [31:0] n27951;
wire     [31:0] n27952;
wire     [31:0] n27953;
wire     [31:0] n27954;
wire     [31:0] n27955;
wire     [31:0] n27956;
wire     [31:0] n27957;
wire     [31:0] n27958;
wire     [31:0] n27959;
wire     [31:0] n27960;
wire     [31:0] n27961;
wire     [31:0] n27962;
wire     [31:0] n27963;
wire     [31:0] n27964;
wire     [31:0] n27965;
wire     [31:0] n27966;
wire     [31:0] n27967;
wire     [31:0] n27968;
wire     [31:0] n27969;
wire     [31:0] n27970;
wire     [31:0] n27971;
wire     [31:0] n27972;
wire     [31:0] n27973;
wire     [31:0] n27974;
wire     [31:0] n27975;
wire     [31:0] n27976;
wire     [31:0] n27977;
wire     [31:0] n27978;
wire     [31:0] n27979;
wire     [31:0] n27980;
wire     [31:0] n27981;
wire     [31:0] n27982;
wire     [31:0] n27983;
wire     [31:0] n27984;
wire     [31:0] n27985;
wire     [31:0] n27986;
wire     [31:0] n27987;
wire     [31:0] n27988;
wire     [31:0] n27989;
wire     [31:0] n27990;
wire     [31:0] n27991;
wire     [31:0] n27992;
wire     [31:0] n27993;
wire     [31:0] n27994;
wire     [31:0] n27995;
wire     [31:0] n27996;
wire     [31:0] n27997;
wire     [31:0] n27998;
wire     [31:0] n27999;
wire     [31:0] n28000;
wire     [31:0] n28001;
wire     [31:0] n28002;
wire     [31:0] n28003;
wire     [31:0] n28004;
wire     [31:0] n28005;
wire     [31:0] n28006;
wire     [31:0] n28007;
wire     [31:0] n28008;
wire     [31:0] n28009;
wire     [31:0] n28010;
wire     [31:0] n28011;
wire     [31:0] n28012;
wire     [31:0] n28013;
wire     [31:0] n28014;
wire     [31:0] n28015;
wire     [31:0] n28016;
wire     [31:0] n28017;
wire     [31:0] n28018;
wire     [31:0] n28019;
wire     [31:0] n28020;
wire     [31:0] n28021;
wire     [31:0] n28022;
wire     [31:0] n28023;
wire     [31:0] n28024;
wire     [31:0] n28025;
wire     [31:0] n28026;
wire     [31:0] n28027;
wire     [31:0] n28028;
wire     [31:0] n28029;
wire     [31:0] n28030;
wire     [31:0] n28031;
wire     [31:0] n28032;
wire     [31:0] n28033;
wire     [31:0] n28034;
wire     [31:0] n28035;
wire     [31:0] n28036;
wire     [31:0] n28037;
wire     [31:0] n28038;
wire     [31:0] n28039;
wire     [31:0] n28040;
wire     [31:0] n28041;
wire     [31:0] n28042;
wire     [31:0] n28043;
wire     [31:0] n28044;
wire     [31:0] n28045;
wire     [31:0] n28046;
wire     [31:0] n28047;
wire     [31:0] n28048;
wire     [31:0] n28049;
wire     [31:0] n28050;
wire     [31:0] n28051;
wire     [31:0] n28052;
wire     [31:0] n28053;
wire     [31:0] n28054;
wire     [31:0] n28055;
wire     [31:0] n28056;
wire     [31:0] n28057;
wire     [31:0] n28058;
wire     [31:0] n28059;
wire     [31:0] n28060;
wire     [31:0] n28061;
wire     [31:0] n28062;
wire     [31:0] n28063;
wire     [31:0] n28064;
wire     [31:0] n28065;
wire     [31:0] n28066;
wire     [31:0] n28067;
wire     [31:0] n28068;
wire     [31:0] n28069;
wire     [31:0] n28070;
wire     [31:0] n28071;
wire     [31:0] n28072;
wire     [31:0] n28073;
wire     [31:0] n28074;
wire     [31:0] n28075;
wire     [31:0] n28076;
wire     [31:0] n28077;
wire     [31:0] n28078;
wire     [31:0] n28079;
wire     [31:0] n28080;
wire     [31:0] n28081;
wire     [31:0] n28082;
wire     [31:0] n28083;
wire     [31:0] n28084;
wire     [31:0] n28085;
wire     [31:0] n28086;
wire     [31:0] n28087;
wire     [31:0] n28088;
wire     [31:0] n28089;
wire     [31:0] n28090;
wire     [31:0] n28091;
wire     [31:0] n28092;
wire     [31:0] n28093;
wire     [31:0] n28094;
wire     [31:0] n28095;
wire     [31:0] n28096;
wire     [31:0] n28097;
wire     [31:0] n28098;
wire     [31:0] n28099;
wire     [31:0] n28100;
wire     [31:0] n28101;
wire     [31:0] n28102;
wire     [31:0] n28103;
wire     [31:0] n28104;
wire     [31:0] n28105;
wire     [31:0] n28106;
wire     [31:0] n28107;
wire     [31:0] n28108;
wire     [31:0] n28109;
wire     [31:0] n28110;
wire     [31:0] n28111;
wire     [31:0] n28112;
wire     [31:0] n28113;
wire     [31:0] n28114;
wire     [31:0] n28115;
wire     [31:0] n28116;
wire     [31:0] n28117;
wire     [31:0] n28118;
wire     [31:0] n28119;
wire     [31:0] n28120;
wire     [31:0] n28121;
wire     [31:0] n28122;
wire     [31:0] n28123;
wire     [31:0] n28124;
wire     [31:0] n28125;
wire     [31:0] n28126;
wire     [31:0] n28127;
wire     [31:0] n28128;
wire     [31:0] n28129;
wire     [31:0] n28130;
wire     [31:0] n28131;
wire     [31:0] n28132;
wire     [31:0] n28133;
wire     [31:0] n28134;
wire     [31:0] n28135;
wire     [31:0] n28136;
wire     [31:0] n28137;
wire     [31:0] n28138;
wire     [31:0] n28139;
wire     [31:0] n28140;
wire     [31:0] n28141;
wire     [31:0] n28142;
wire     [31:0] n28143;
wire     [31:0] n28144;
wire     [31:0] n28145;
wire     [31:0] n28146;
wire     [31:0] n28147;
wire     [31:0] n28148;
wire     [31:0] n28149;
wire     [31:0] n28150;
wire     [31:0] n28151;
wire     [31:0] n28152;
wire     [31:0] n28153;
wire     [31:0] n28154;
wire     [31:0] n28155;
wire     [31:0] n28156;
wire     [31:0] n28157;
wire     [31:0] n28158;
wire     [31:0] n28159;
wire     [31:0] n28160;
wire     [31:0] n28161;
wire     [31:0] n28162;
wire     [31:0] n28163;
wire     [31:0] n28164;
wire     [31:0] n28165;
wire     [31:0] n28166;
wire     [31:0] n28167;
wire     [31:0] n28168;
wire     [31:0] n28169;
wire     [31:0] n28170;
wire     [31:0] n28171;
wire     [31:0] n28172;
wire     [31:0] n28173;
wire     [31:0] n28174;
wire     [31:0] n28175;
wire     [31:0] n28176;
wire     [31:0] n28177;
wire     [31:0] n28178;
wire     [31:0] n28179;
wire     [31:0] n28180;
wire     [31:0] n28181;
wire     [31:0] n28182;
wire     [31:0] n28183;
wire     [31:0] n28184;
wire     [31:0] n28185;
wire     [31:0] n28186;
wire     [31:0] n28187;
wire     [31:0] n28188;
wire     [31:0] n28189;
wire     [31:0] n28190;
wire     [31:0] n28191;
wire     [31:0] n28192;
wire     [31:0] n28193;
wire     [31:0] n28194;
wire     [31:0] n28195;
wire     [31:0] n28196;
wire     [31:0] n28197;
wire     [31:0] n28198;
wire     [31:0] n28199;
wire     [31:0] n28200;
wire     [31:0] n28201;
wire     [31:0] n28202;
wire     [31:0] n28203;
wire     [31:0] n28204;
wire     [31:0] n28205;
wire     [31:0] n28206;
wire     [31:0] n28207;
wire     [31:0] n28208;
wire     [31:0] n28209;
wire     [31:0] n28210;
wire     [31:0] n28211;
wire     [31:0] n28212;
wire     [31:0] n28213;
wire     [31:0] n28214;
wire     [31:0] n28215;
wire     [31:0] n28216;
wire     [31:0] n28217;
wire     [31:0] n28218;
wire     [31:0] n28219;
wire     [31:0] n28220;
wire     [31:0] n28221;
wire     [31:0] n28222;
wire     [31:0] n28223;
wire     [31:0] n28224;
wire     [31:0] n28225;
wire     [31:0] n28226;
wire     [31:0] n28227;
wire     [31:0] n28228;
wire     [31:0] n28229;
wire     [31:0] n28230;
wire     [31:0] n28231;
wire     [31:0] n28232;
wire     [31:0] n28233;
wire     [31:0] n28234;
wire     [31:0] n28235;
wire     [31:0] n28236;
wire     [31:0] n28237;
wire     [31:0] n28238;
wire     [31:0] n28239;
wire     [31:0] n28240;
wire     [31:0] n28241;
wire     [31:0] n28242;
wire     [31:0] n28243;
wire     [31:0] n28244;
wire     [31:0] n28245;
wire     [31:0] n28246;
wire     [31:0] n28247;
wire     [31:0] n28248;
wire     [31:0] n28249;
wire     [31:0] n28250;
wire     [31:0] n28251;
wire     [31:0] n28252;
wire     [31:0] n28253;
wire     [31:0] n28254;
wire     [31:0] n28255;
wire     [31:0] n28256;
wire     [31:0] n28257;
wire     [31:0] n28258;
wire     [31:0] n28259;
wire     [31:0] n28260;
wire     [31:0] n28261;
wire     [31:0] n28262;
wire     [31:0] n28263;
wire     [31:0] n28264;
wire     [31:0] n28265;
wire     [31:0] n28266;
wire     [31:0] n28267;
wire     [31:0] n28268;
wire     [31:0] n28269;
wire     [31:0] n28270;
wire     [31:0] n28271;
wire     [31:0] n28272;
wire     [31:0] n28273;
wire     [31:0] n28274;
wire     [31:0] n28275;
wire     [31:0] n28276;
wire     [31:0] n28277;
wire     [31:0] n28278;
wire     [31:0] n28279;
wire     [31:0] n28280;
wire     [31:0] n28281;
wire     [31:0] n28282;
wire     [31:0] n28283;
wire     [31:0] n28284;
wire     [31:0] n28285;
wire     [31:0] n28286;
wire     [31:0] n28287;
wire     [31:0] n28288;
wire     [31:0] n28289;
wire     [31:0] n28290;
wire     [31:0] n28291;
wire     [31:0] n28292;
wire     [31:0] n28293;
wire     [31:0] n28294;
wire     [31:0] n28295;
wire     [31:0] n28296;
wire     [31:0] n28297;
wire     [31:0] n28298;
wire     [31:0] n28299;
wire     [31:0] n28300;
wire     [31:0] n28301;
wire     [31:0] n28302;
wire     [31:0] n28303;
wire     [31:0] n28304;
wire     [31:0] n28305;
wire     [31:0] n28306;
wire     [31:0] n28307;
wire     [31:0] n28308;
wire     [31:0] n28309;
wire     [31:0] n28310;
wire     [31:0] n28311;
wire     [31:0] n28312;
wire     [31:0] n28313;
wire     [31:0] n28314;
wire     [31:0] n28315;
wire     [31:0] n28316;
wire     [31:0] n28317;
wire     [31:0] n28318;
wire     [31:0] n28319;
wire     [31:0] n28320;
wire     [31:0] n28321;
wire     [31:0] n28322;
wire     [31:0] n28323;
wire     [31:0] n28324;
wire     [31:0] n28325;
wire     [31:0] n28326;
wire     [31:0] n28327;
wire     [31:0] n28328;
wire     [31:0] n28329;
wire     [31:0] n28330;
wire     [31:0] n28331;
wire     [31:0] n28332;
wire     [31:0] n28333;
wire     [31:0] n28334;
wire     [31:0] n28335;
wire     [31:0] n28336;
wire     [31:0] n28337;
wire     [31:0] n28338;
wire     [31:0] n28339;
wire     [31:0] n28340;
wire     [31:0] n28341;
wire     [31:0] n28342;
wire     [31:0] n28343;
wire     [31:0] n28344;
wire     [31:0] n28345;
wire     [31:0] n28346;
wire     [31:0] n28347;
wire     [31:0] n28348;
wire     [31:0] n28349;
wire     [31:0] n28350;
wire     [31:0] n28351;
wire     [31:0] n28352;
wire     [31:0] n28353;
wire     [31:0] n28354;
wire     [31:0] n28355;
wire     [31:0] n28356;
wire     [31:0] n28357;
wire     [31:0] n28358;
wire     [31:0] n28359;
wire     [31:0] n28360;
wire     [31:0] n28361;
wire     [31:0] n28362;
wire     [31:0] n28363;
wire     [31:0] n28364;
wire     [31:0] n28365;
wire     [31:0] n28366;
wire     [31:0] n28367;
wire     [31:0] n28368;
wire     [31:0] n28369;
wire     [31:0] n28370;
wire     [31:0] n28371;
wire     [31:0] n28372;
wire     [31:0] n28373;
wire     [31:0] n28374;
wire     [31:0] n28375;
wire     [31:0] n28376;
wire     [31:0] n28377;
wire     [31:0] n28378;
wire     [31:0] n28379;
wire     [31:0] n28380;
wire     [31:0] n28381;
wire     [31:0] n28382;
wire     [31:0] n28383;
wire     [31:0] n28384;
wire     [31:0] n28385;
wire     [31:0] n28386;
wire     [31:0] n28387;
wire     [31:0] n28388;
wire     [31:0] n28389;
wire     [31:0] n28390;
wire     [31:0] n28391;
wire     [31:0] n28392;
wire     [31:0] n28393;
wire     [31:0] n28394;
wire     [31:0] n28395;
wire     [31:0] n28396;
wire     [31:0] n28397;
wire     [31:0] n28398;
wire     [31:0] n28399;
wire     [31:0] n28400;
wire     [31:0] n28401;
wire     [31:0] n28402;
wire     [31:0] n28403;
wire     [31:0] n28404;
wire     [31:0] n28405;
wire     [31:0] n28406;
wire     [31:0] n28407;
wire     [31:0] n28408;
wire     [31:0] n28409;
wire     [31:0] n28410;
wire     [31:0] n28411;
wire     [31:0] n28412;
wire     [31:0] n28413;
wire     [31:0] n28414;
wire     [31:0] n28415;
wire     [31:0] n28416;
wire     [31:0] n28417;
wire     [31:0] n28418;
wire     [31:0] n28419;
wire     [31:0] n28420;
wire     [31:0] n28421;
wire     [31:0] n28422;
wire     [31:0] n28423;
wire     [31:0] n28424;
wire     [31:0] n28425;
wire     [31:0] n28426;
wire     [31:0] n28427;
wire     [31:0] n28428;
wire     [31:0] n28429;
wire     [31:0] n28430;
wire     [31:0] n28431;
wire     [31:0] n28432;
wire     [31:0] n28433;
wire     [31:0] n28434;
wire     [31:0] n28435;
wire     [31:0] n28436;
wire     [31:0] n28437;
wire     [31:0] n28438;
wire     [31:0] n28439;
wire     [31:0] n28440;
wire     [31:0] n28441;
wire     [31:0] n28442;
wire     [31:0] n28443;
wire     [31:0] n28444;
wire     [31:0] n28445;
wire     [31:0] n28446;
wire     [31:0] n28447;
wire     [31:0] n28448;
wire     [31:0] n28449;
wire     [31:0] n28450;
wire     [31:0] n28451;
wire     [31:0] n28452;
wire     [31:0] n28453;
wire     [31:0] n28454;
wire     [31:0] n28455;
wire     [31:0] n28456;
wire     [31:0] n28457;
wire     [31:0] n28458;
wire     [31:0] n28459;
wire     [31:0] n28460;
wire     [31:0] n28461;
wire            n28462;
wire            n28463;
wire     [31:0] n28464;
wire     [31:0] n28465;
wire     [31:0] n28466;
wire     [31:0] n28467;
wire     [31:0] n28468;
wire     [31:0] n28469;
wire     [31:0] n28470;
wire     [31:0] n28471;
wire     [31:0] n28472;
wire     [31:0] n28473;
wire     [31:0] n28474;
wire     [31:0] n28475;
wire     [31:0] n28476;
wire     [31:0] n28477;
wire     [31:0] n28478;
wire     [31:0] n28479;
wire     [31:0] n28480;
wire     [31:0] n28481;
wire     [31:0] n28482;
wire     [31:0] n28483;
wire     [31:0] n28484;
wire     [31:0] n28485;
wire     [31:0] n28486;
wire     [31:0] n28487;
wire     [31:0] n28488;
wire     [31:0] n28489;
wire     [31:0] n28490;
wire     [31:0] n28491;
wire     [31:0] n28492;
wire     [31:0] n28493;
wire     [31:0] n28494;
wire     [31:0] n28495;
wire     [31:0] n28496;
wire            n28497;
wire            n28498;
wire            n28499;
wire            n28500;
wire            n28501;
wire            n28502;
wire            n28503;
wire            n28504;
wire            n28505;
wire            n28506;
wire            n28507;
wire            n28508;
wire            n28509;
wire            n28510;
wire            n28511;
wire            n28512;
wire            n28513;
wire            n28514;
wire            n28515;
wire            n28516;
wire            n28517;
wire            n28518;
wire            n28519;
wire            n28520;
wire            n28521;
wire            n28522;
wire            n28523;
wire            n28524;
wire            n28525;
wire            n28526;
wire            n28527;
wire            n28528;
wire            n28529;
wire            n28530;
wire            n28531;
wire            n28532;
wire            n28533;
wire            n28534;
wire            n28535;
wire            n28536;
wire            n28537;
wire            n28538;
wire            n28539;
wire            n28540;
wire            n28541;
wire            n28542;
wire            n28543;
wire            n28544;
wire            n28545;
wire            n28546;
wire            n28547;
wire            n28548;
wire            n28549;
wire            n28550;
wire            n28551;
wire            n28552;
wire            n28553;
wire            n28554;
wire            n28555;
wire            n28556;
wire            n28557;
wire            n28558;
wire            n28559;
wire            n28560;
wire            n28561;
wire            n28562;
wire            n28563;
wire            n28564;
wire            n28565;
wire            n28566;
wire            n28567;
wire            n28568;
wire            n28569;
wire            n28570;
wire            n28571;
wire            n28572;
wire            n28573;
wire            n28574;
wire            n28575;
wire            n28576;
wire            n28577;
wire            n28578;
wire            n28579;
wire            n28580;
wire            n28581;
wire            n28582;
wire            n28583;
wire            n28584;
wire            n28585;
wire            n28586;
wire            n28587;
wire            n28588;
wire            n28589;
wire            n28590;
wire            n28591;
wire            n28592;
wire            n28593;
wire            n28594;
wire            n28595;
wire            n28596;
wire            n28597;
wire            n28598;
wire            n28599;
wire            n28600;
wire            n28601;
wire            n28602;
wire            n28603;
wire            n28604;
wire            n28605;
wire            n28606;
wire            n28607;
wire            n28608;
wire            n28609;
wire            n28610;
wire            n28611;
wire            n28612;
wire            n28613;
wire            n28614;
wire            n28615;
wire            n28616;
wire            n28617;
wire            n28618;
wire            n28619;
wire            n28620;
wire            n28621;
wire            n28622;
wire            n28623;
wire            n28624;
wire            n28625;
wire            n28626;
wire            n28627;
wire            n28628;
wire            n28629;
wire            n28630;
wire            n28631;
wire            n28632;
wire            n28633;
wire            n28634;
wire            n28635;
wire            n28636;
wire            n28637;
wire            n28638;
wire            n28639;
wire            n28640;
wire            n28641;
wire            n28642;
wire            n28643;
wire            n28644;
wire            n28645;
wire            n28646;
wire            n28647;
wire            n28648;
wire            n28649;
wire            n28650;
wire            n28651;
wire            n28652;
wire            n28653;
wire            n28654;
wire            n28655;
wire            n28656;
wire            n28657;
wire            n28658;
wire            n28659;
wire            n28660;
wire            n28661;
wire            n28662;
wire            n28663;
wire            n28664;
wire            n28665;
wire            n28666;
wire            n28667;
wire            n28668;
wire            n28669;
wire            n28670;
wire            n28671;
wire            n28672;
wire            n28673;
wire            n28674;
wire            n28675;
wire            n28676;
wire            n28677;
wire            n28678;
wire            n28679;
wire            n28680;
wire            n28681;
wire            n28682;
wire            n28683;
wire            n28684;
wire            n28685;
wire            n28686;
wire            n28687;
wire            n28688;
wire            n28689;
wire            n28690;
wire            n28691;
wire            n28692;
wire            n28693;
wire            n28694;
wire            n28695;
wire            n28696;
wire            n28697;
wire            n28698;
wire            n28699;
wire            n28700;
wire            n28701;
wire            n28702;
wire            n28703;
wire            n28704;
wire            n28705;
wire            n28706;
wire            n28707;
wire            n28708;
wire            n28709;
wire            n28710;
wire            n28711;
wire            n28712;
wire            n28713;
wire            n28714;
wire            n28715;
wire            n28716;
wire            n28717;
wire            n28718;
wire            n28719;
wire            n28720;
wire            n28721;
wire            n28722;
wire            n28723;
wire            n28724;
wire            n28725;
wire            n28726;
wire            n28727;
wire            n28728;
wire            n28729;
wire            n28730;
wire            n28731;
wire            n28732;
wire            n28733;
wire            n28734;
wire            n28735;
wire            n28736;
wire            n28737;
wire            n28738;
wire            n28739;
wire            n28740;
wire            n28741;
wire            n28742;
wire            n28743;
wire            n28744;
wire            n28745;
wire            n28746;
wire            n28747;
wire            n28748;
wire            n28749;
wire            n28750;
wire            n28751;
wire            n28752;
wire            n28753;
wire            n28754;
wire            n28755;
wire            n28756;
wire            n28757;
wire            n28758;
wire            n28759;
wire            n28760;
wire            n28761;
wire            n28762;
wire            n28763;
wire            n28764;
wire            n28765;
wire            n28766;
wire            n28767;
wire            n28768;
wire            n28769;
wire            n28770;
wire            n28771;
wire            n28772;
wire            n28773;
wire            n28774;
wire            n28775;
wire            n28776;
wire            n28777;
wire            n28778;
wire            n28779;
wire            n28780;
wire            n28781;
wire            n28782;
wire            n28783;
wire            n28784;
wire            n28785;
wire            n28786;
wire            n28787;
wire            n28788;
wire            n28789;
wire            n28790;
wire            n28791;
wire            n28792;
wire            n28793;
wire            n28794;
wire            n28795;
wire            n28796;
wire            n28797;
wire            n28798;
wire            n28799;
wire            n28800;
wire            n28801;
wire            n28802;
wire            n28803;
wire            n28804;
wire            n28805;
wire            n28806;
wire            n28807;
wire            n28808;
wire            n28809;
wire            n28810;
wire            n28811;
wire            n28812;
wire            n28813;
wire            n28814;
wire            n28815;
wire            n28816;
wire            n28817;
wire            n28818;
wire            n28819;
wire            n28820;
wire            n28821;
wire            n28822;
wire            n28823;
wire            n28824;
wire            n28825;
wire            n28826;
wire            n28827;
wire            n28828;
wire            n28829;
wire            n28830;
wire            n28831;
wire            n28832;
wire            n28833;
wire            n28834;
wire            n28835;
wire            n28836;
wire            n28837;
wire            n28838;
wire            n28839;
wire            n28840;
wire            n28841;
wire            n28842;
wire            n28843;
wire            n28844;
wire            n28845;
wire            n28846;
wire            n28847;
wire            n28848;
wire            n28849;
wire            n28850;
wire            n28851;
wire            n28852;
wire            n28853;
wire            n28854;
wire            n28855;
wire            n28856;
wire            n28857;
wire            n28858;
wire            n28859;
wire            n28860;
wire            n28861;
wire            n28862;
wire            n28863;
wire            n28864;
wire            n28865;
wire            n28866;
wire            n28867;
wire            n28868;
wire            n28869;
wire            n28870;
wire            n28871;
wire            n28872;
wire            n28873;
wire            n28874;
wire            n28875;
wire            n28876;
wire            n28877;
wire            n28878;
wire            n28879;
wire            n28880;
wire            n28881;
wire            n28882;
wire            n28883;
wire            n28884;
wire            n28885;
wire            n28886;
wire            n28887;
wire            n28888;
wire            n28889;
wire            n28890;
wire            n28891;
wire            n28892;
wire            n28893;
wire            n28894;
wire            n28895;
wire            n28896;
wire            n28897;
wire            n28898;
wire            n28899;
wire            n28900;
wire            n28901;
wire            n28902;
wire            n28903;
wire            n28904;
wire            n28905;
wire            n28906;
wire            n28907;
wire            n28908;
wire            n28909;
wire            n28910;
wire            n28911;
wire            n28912;
wire            n28913;
wire            n28914;
wire            n28915;
wire            n28916;
wire            n28917;
wire            n28918;
wire            n28919;
wire            n28920;
wire            n28921;
wire            n28922;
wire            n28923;
wire            n28924;
wire            n28925;
wire            n28926;
wire            n28927;
wire            n28928;
wire            n28929;
wire            n28930;
wire            n28931;
wire            n28932;
wire            n28933;
wire            n28934;
wire            n28935;
wire            n28936;
wire            n28937;
wire            n28938;
wire            n28939;
wire            n28940;
wire            n28941;
wire            n28942;
wire            n28943;
wire            n28944;
wire            n28945;
wire            n28946;
wire            n28947;
wire            n28948;
wire            n28949;
wire            n28950;
wire            n28951;
wire            n28952;
wire            n28953;
wire            n28954;
wire            n28955;
wire            n28956;
wire            n28957;
wire            n28958;
wire            n28959;
wire            n28960;
wire            n28961;
wire            n28962;
wire            n28963;
wire            n28964;
wire            n28965;
wire            n28966;
wire            n28967;
wire            n28968;
wire            n28969;
wire            n28970;
wire            n28971;
wire            n28972;
wire            n28973;
wire            n28974;
wire            n28975;
wire            n28976;
wire            n28977;
wire            n28978;
wire            n28979;
wire            n28980;
wire            n28981;
wire            n28982;
wire            n28983;
wire            n28984;
wire            n28985;
wire            n28986;
wire            n28987;
wire            n28988;
wire            n28989;
wire            n28990;
wire            n28991;
wire            n28992;
wire            n28993;
wire            n28994;
wire            n28995;
wire            n28996;
wire            n28997;
wire            n28998;
wire            n28999;
wire            n29000;
wire            n29001;
wire            n29002;
wire            n29003;
wire            n29004;
wire            n29005;
wire            n29006;
wire            n29007;
wire            n29008;
wire            n29009;
wire            n29010;
wire            n29011;
wire            n29012;
wire            n29013;
wire            n29014;
wire            n29015;
wire            n29016;
wire            n29017;
wire            n29018;
wire            n29019;
wire            n29020;
wire            n29021;
wire            n29022;
wire            n29023;
wire            n29024;
wire     [31:0] n29025;
wire     [31:0] n29026;
wire     [31:0] n29027;
wire     [31:0] n29028;
wire     [31:0] n29029;
wire     [31:0] n29030;
wire     [31:0] n29031;
wire     [31:0] n29032;
wire     [31:0] n29033;
wire     [31:0] n29034;
wire     [31:0] n29035;
wire     [31:0] n29036;
wire     [31:0] n29037;
wire     [31:0] n29038;
wire     [31:0] n29039;
wire     [31:0] n29040;
wire     [31:0] n29041;
wire     [31:0] n29042;
wire     [31:0] n29043;
wire     [31:0] n29044;
wire     [31:0] n29045;
wire     [31:0] n29046;
wire     [31:0] n29047;
wire     [31:0] n29048;
wire     [31:0] n29049;
wire     [31:0] n29050;
wire     [31:0] n29051;
wire     [31:0] n29052;
wire     [31:0] n29053;
wire     [31:0] n29054;
wire     [31:0] n29055;
wire     [31:0] n29056;
wire     [31:0] n29057;
wire     [31:0] n29058;
wire     [31:0] n29059;
wire     [31:0] n29060;
wire     [31:0] n29061;
wire     [31:0] n29062;
wire     [31:0] n29063;
wire     [31:0] n29064;
wire     [31:0] n29065;
wire     [31:0] n29066;
wire     [31:0] n29067;
wire     [31:0] n29068;
wire     [31:0] n29069;
wire     [31:0] n29070;
wire     [31:0] n29071;
wire     [31:0] n29072;
wire     [31:0] n29073;
wire     [31:0] n29074;
wire     [31:0] n29075;
wire     [31:0] n29076;
wire     [31:0] n29077;
wire     [31:0] n29078;
wire     [31:0] n29079;
wire     [31:0] n29080;
wire     [31:0] n29081;
wire     [31:0] n29082;
wire     [31:0] n29083;
wire     [31:0] n29084;
wire     [31:0] n29085;
wire     [31:0] n29086;
wire     [31:0] n29087;
wire     [31:0] n29088;
wire     [31:0] n29089;
wire     [31:0] n29090;
wire     [31:0] n29091;
wire     [31:0] n29092;
wire     [31:0] n29093;
wire     [31:0] n29094;
wire     [31:0] n29095;
wire     [31:0] n29096;
wire     [31:0] n29097;
wire     [31:0] n29098;
wire     [31:0] n29099;
wire     [31:0] n29100;
wire     [31:0] n29101;
wire     [31:0] n29102;
wire     [31:0] n29103;
wire     [31:0] n29104;
wire     [31:0] n29105;
wire     [31:0] n29106;
wire     [31:0] n29107;
wire     [31:0] n29108;
wire     [31:0] n29109;
wire     [31:0] n29110;
wire     [31:0] n29111;
wire     [31:0] n29112;
wire     [31:0] n29113;
wire     [31:0] n29114;
wire     [31:0] n29115;
wire     [31:0] n29116;
wire     [31:0] n29117;
wire     [31:0] n29118;
wire     [31:0] n29119;
wire     [31:0] n29120;
wire     [31:0] n29121;
wire     [31:0] n29122;
wire     [31:0] n29123;
wire     [31:0] n29124;
wire     [31:0] n29125;
wire     [31:0] n29126;
wire     [31:0] n29127;
wire     [31:0] n29128;
wire     [31:0] n29129;
wire     [31:0] n29130;
wire     [31:0] n29131;
wire     [31:0] n29132;
wire     [31:0] n29133;
wire     [31:0] n29134;
wire     [31:0] n29135;
wire     [31:0] n29136;
wire     [31:0] n29137;
wire     [31:0] n29138;
wire     [31:0] n29139;
wire     [31:0] n29140;
wire     [31:0] n29141;
wire     [31:0] n29142;
wire     [31:0] n29143;
wire     [31:0] n29144;
wire     [31:0] n29145;
wire     [31:0] n29146;
wire     [31:0] n29147;
wire     [31:0] n29148;
wire     [31:0] n29149;
wire     [31:0] n29150;
wire     [31:0] n29151;
wire     [31:0] n29152;
wire     [31:0] n29153;
wire     [31:0] n29154;
wire     [31:0] n29155;
wire     [31:0] n29156;
wire     [31:0] n29157;
wire     [31:0] n29158;
wire     [31:0] n29159;
wire     [31:0] n29160;
wire     [31:0] n29161;
wire     [31:0] n29162;
wire     [31:0] n29163;
wire     [31:0] n29164;
wire     [31:0] n29165;
wire     [31:0] n29166;
wire     [31:0] n29167;
wire     [31:0] n29168;
wire     [31:0] n29169;
wire     [31:0] n29170;
wire     [31:0] n29171;
wire     [31:0] n29172;
wire     [31:0] n29173;
wire     [31:0] n29174;
wire     [31:0] n29175;
wire     [31:0] n29176;
wire     [31:0] n29177;
wire     [31:0] n29178;
wire     [31:0] n29179;
wire     [31:0] n29180;
wire     [31:0] n29181;
wire     [31:0] n29182;
wire     [31:0] n29183;
wire     [31:0] n29184;
wire     [31:0] n29185;
wire     [31:0] n29186;
wire     [31:0] n29187;
wire     [31:0] n29188;
wire     [31:0] n29189;
wire     [31:0] n29190;
wire     [31:0] n29191;
wire     [31:0] n29192;
wire     [31:0] n29193;
wire     [31:0] n29194;
wire     [31:0] n29195;
wire     [31:0] n29196;
wire     [31:0] n29197;
wire     [31:0] n29198;
wire     [31:0] n29199;
wire     [31:0] n29200;
wire     [31:0] n29201;
wire     [31:0] n29202;
wire     [31:0] n29203;
wire     [31:0] n29204;
wire     [31:0] n29205;
wire     [31:0] n29206;
wire     [31:0] n29207;
wire     [31:0] n29208;
wire     [31:0] n29209;
wire     [31:0] n29210;
wire     [31:0] n29211;
wire     [31:0] n29212;
wire     [31:0] n29213;
wire     [31:0] n29214;
wire     [31:0] n29215;
wire     [31:0] n29216;
wire     [31:0] n29217;
wire     [31:0] n29218;
wire     [31:0] n29219;
wire     [31:0] n29220;
wire     [31:0] n29221;
wire     [31:0] n29222;
wire     [31:0] n29223;
wire     [31:0] n29224;
wire     [31:0] n29225;
wire     [31:0] n29226;
wire     [31:0] n29227;
wire     [31:0] n29228;
wire     [31:0] n29229;
wire     [31:0] n29230;
wire     [31:0] n29231;
wire     [31:0] n29232;
wire     [31:0] n29233;
wire     [31:0] n29234;
wire     [31:0] n29235;
wire     [31:0] n29236;
wire     [31:0] n29237;
wire     [31:0] n29238;
wire     [31:0] n29239;
wire     [31:0] n29240;
wire     [31:0] n29241;
wire     [31:0] n29242;
wire     [31:0] n29243;
wire     [31:0] n29244;
wire     [31:0] n29245;
wire     [31:0] n29246;
wire     [31:0] n29247;
wire     [31:0] n29248;
wire     [31:0] n29249;
wire     [31:0] n29250;
wire     [31:0] n29251;
wire     [31:0] n29252;
wire     [31:0] n29253;
wire     [31:0] n29254;
wire     [31:0] n29255;
wire     [31:0] n29256;
wire     [31:0] n29257;
wire     [31:0] n29258;
wire     [31:0] n29259;
wire     [31:0] n29260;
wire     [31:0] n29261;
wire     [31:0] n29262;
wire     [31:0] n29263;
wire     [31:0] n29264;
wire     [31:0] n29265;
wire     [31:0] n29266;
wire     [31:0] n29267;
wire     [31:0] n29268;
wire     [31:0] n29269;
wire     [31:0] n29270;
wire     [31:0] n29271;
wire     [31:0] n29272;
wire     [31:0] n29273;
wire     [31:0] n29274;
wire     [31:0] n29275;
wire     [31:0] n29276;
wire     [31:0] n29277;
wire     [31:0] n29278;
wire     [31:0] n29279;
wire     [31:0] n29280;
wire     [31:0] n29281;
wire     [31:0] n29282;
wire     [31:0] n29283;
wire     [31:0] n29284;
wire     [31:0] n29285;
wire     [31:0] n29286;
wire     [31:0] n29287;
wire     [31:0] n29288;
wire     [31:0] n29289;
wire     [31:0] n29290;
wire     [31:0] n29291;
wire     [31:0] n29292;
wire     [31:0] n29293;
wire     [31:0] n29294;
wire     [31:0] n29295;
wire     [31:0] n29296;
wire     [31:0] n29297;
wire     [31:0] n29298;
wire     [31:0] n29299;
wire     [31:0] n29300;
wire     [31:0] n29301;
wire     [31:0] n29302;
wire     [31:0] n29303;
wire     [31:0] n29304;
wire     [31:0] n29305;
wire     [31:0] n29306;
wire     [31:0] n29307;
wire     [31:0] n29308;
wire     [31:0] n29309;
wire     [31:0] n29310;
wire     [31:0] n29311;
wire     [31:0] n29312;
wire     [31:0] n29313;
wire     [31:0] n29314;
wire     [31:0] n29315;
wire     [31:0] n29316;
wire     [31:0] n29317;
wire     [31:0] n29318;
wire     [31:0] n29319;
wire     [31:0] n29320;
wire     [31:0] n29321;
wire     [31:0] n29322;
wire     [31:0] n29323;
wire     [31:0] n29324;
wire     [31:0] n29325;
wire     [31:0] n29326;
wire     [31:0] n29327;
wire     [31:0] n29328;
wire     [31:0] n29329;
wire     [31:0] n29330;
wire     [31:0] n29331;
wire     [31:0] n29332;
wire     [31:0] n29333;
wire     [31:0] n29334;
wire     [31:0] n29335;
wire     [31:0] n29336;
wire     [31:0] n29337;
wire     [31:0] n29338;
wire     [31:0] n29339;
wire     [31:0] n29340;
wire     [31:0] n29341;
wire     [31:0] n29342;
wire     [31:0] n29343;
wire     [31:0] n29344;
wire     [31:0] n29345;
wire     [31:0] n29346;
wire     [31:0] n29347;
wire     [31:0] n29348;
wire     [31:0] n29349;
wire     [31:0] n29350;
wire     [31:0] n29351;
wire     [31:0] n29352;
wire     [31:0] n29353;
wire     [31:0] n29354;
wire     [31:0] n29355;
wire     [31:0] n29356;
wire     [31:0] n29357;
wire     [31:0] n29358;
wire     [31:0] n29359;
wire     [31:0] n29360;
wire     [31:0] n29361;
wire     [31:0] n29362;
wire     [31:0] n29363;
wire     [31:0] n29364;
wire     [31:0] n29365;
wire     [31:0] n29366;
wire     [31:0] n29367;
wire     [31:0] n29368;
wire     [31:0] n29369;
wire     [31:0] n29370;
wire     [31:0] n29371;
wire     [31:0] n29372;
wire     [31:0] n29373;
wire     [31:0] n29374;
wire     [31:0] n29375;
wire     [31:0] n29376;
wire     [31:0] n29377;
wire     [31:0] n29378;
wire     [31:0] n29379;
wire     [31:0] n29380;
wire     [31:0] n29381;
wire     [31:0] n29382;
wire     [31:0] n29383;
wire     [31:0] n29384;
wire     [31:0] n29385;
wire     [31:0] n29386;
wire     [31:0] n29387;
wire     [31:0] n29388;
wire     [31:0] n29389;
wire     [31:0] n29390;
wire     [31:0] n29391;
wire     [31:0] n29392;
wire     [31:0] n29393;
wire     [31:0] n29394;
wire     [31:0] n29395;
wire     [31:0] n29396;
wire     [31:0] n29397;
wire     [31:0] n29398;
wire     [31:0] n29399;
wire     [31:0] n29400;
wire     [31:0] n29401;
wire     [31:0] n29402;
wire     [31:0] n29403;
wire     [31:0] n29404;
wire     [31:0] n29405;
wire     [31:0] n29406;
wire     [31:0] n29407;
wire     [31:0] n29408;
wire     [31:0] n29409;
wire     [31:0] n29410;
wire     [31:0] n29411;
wire     [31:0] n29412;
wire     [31:0] n29413;
wire     [31:0] n29414;
wire     [31:0] n29415;
wire     [31:0] n29416;
wire     [31:0] n29417;
wire     [31:0] n29418;
wire     [31:0] n29419;
wire     [31:0] n29420;
wire     [31:0] n29421;
wire     [31:0] n29422;
wire     [31:0] n29423;
wire     [31:0] n29424;
wire     [31:0] n29425;
wire     [31:0] n29426;
wire     [31:0] n29427;
wire     [31:0] n29428;
wire     [31:0] n29429;
wire     [31:0] n29430;
wire     [31:0] n29431;
wire     [31:0] n29432;
wire     [31:0] n29433;
wire     [31:0] n29434;
wire     [31:0] n29435;
wire     [31:0] n29436;
wire     [31:0] n29437;
wire     [31:0] n29438;
wire     [31:0] n29439;
wire     [31:0] n29440;
wire     [31:0] n29441;
wire     [31:0] n29442;
wire     [31:0] n29443;
wire     [31:0] n29444;
wire     [31:0] n29445;
wire     [31:0] n29446;
wire     [31:0] n29447;
wire     [31:0] n29448;
wire     [31:0] n29449;
wire     [31:0] n29450;
wire     [31:0] n29451;
wire     [31:0] n29452;
wire     [31:0] n29453;
wire     [31:0] n29454;
wire     [31:0] n29455;
wire     [31:0] n29456;
wire     [31:0] n29457;
wire     [31:0] n29458;
wire     [31:0] n29459;
wire     [31:0] n29460;
wire     [31:0] n29461;
wire     [31:0] n29462;
wire     [31:0] n29463;
wire     [31:0] n29464;
wire     [31:0] n29465;
wire     [31:0] n29466;
wire     [31:0] n29467;
wire     [31:0] n29468;
wire     [31:0] n29469;
wire     [31:0] n29470;
wire     [31:0] n29471;
wire     [31:0] n29472;
wire     [31:0] n29473;
wire     [31:0] n29474;
wire     [31:0] n29475;
wire     [31:0] n29476;
wire     [31:0] n29477;
wire     [31:0] n29478;
wire     [31:0] n29479;
wire     [31:0] n29480;
wire     [31:0] n29481;
wire     [31:0] n29482;
wire     [31:0] n29483;
wire     [31:0] n29484;
wire     [31:0] n29485;
wire     [31:0] n29486;
wire     [31:0] n29487;
wire     [31:0] n29488;
wire     [31:0] n29489;
wire     [31:0] n29490;
wire     [31:0] n29491;
wire     [31:0] n29492;
wire     [31:0] n29493;
wire     [31:0] n29494;
wire     [31:0] n29495;
wire     [31:0] n29496;
wire     [31:0] n29497;
wire     [31:0] n29498;
wire     [31:0] n29499;
wire     [31:0] n29500;
wire     [31:0] n29501;
wire     [31:0] n29502;
wire     [31:0] n29503;
wire     [31:0] n29504;
wire     [31:0] n29505;
wire     [31:0] n29506;
wire     [31:0] n29507;
wire     [31:0] n29508;
wire     [31:0] n29509;
wire     [31:0] n29510;
wire     [31:0] n29511;
wire     [31:0] n29512;
wire     [31:0] n29513;
wire     [31:0] n29514;
wire     [31:0] n29515;
wire     [31:0] n29516;
wire     [31:0] n29517;
wire     [31:0] n29518;
wire     [31:0] n29519;
wire     [31:0] n29520;
wire     [31:0] n29521;
wire     [31:0] n29522;
wire     [31:0] n29523;
wire     [31:0] n29524;
wire     [31:0] n29525;
wire     [31:0] n29526;
wire     [31:0] n29527;
wire     [31:0] n29528;
wire     [31:0] n29529;
wire     [31:0] n29530;
wire     [31:0] n29531;
wire     [31:0] n29532;
wire     [31:0] n29533;
wire     [31:0] n29534;
wire     [31:0] n29535;
wire     [31:0] n29536;
wire     [31:0] n29537;
wire     [31:0] n29538;
wire     [31:0] n29539;
wire     [31:0] n29540;
wire     [31:0] n29541;
wire     [31:0] n29542;
wire     [31:0] n29543;
wire     [31:0] n29544;
wire     [31:0] n29545;
wire     [31:0] n29546;
wire            n29547;
wire            n29548;
wire            n29549;
wire            n29550;
wire            n29551;
wire            n29552;
wire            n29553;
wire            n29554;
wire            n29555;
wire            n29556;
wire            n29557;
wire            n29558;
wire            n29559;
wire            n29560;
wire            n29561;
wire            n29562;
wire            n29563;
wire            n29564;
wire            n29565;
wire            n29566;
wire            n29567;
wire            n29568;
wire            n29569;
wire            n29570;
wire            n29571;
wire            n29572;
wire            n29573;
wire            n29574;
wire            n29575;
wire            n29576;
wire            n29577;
wire            n29578;
wire            n29579;
wire            n29580;
wire            n29581;
wire            n29582;
wire            n29583;
wire            n29584;
wire            n29585;
wire            n29586;
wire            n29587;
wire            n29588;
wire            n29589;
wire            n29590;
wire            n29591;
wire            n29592;
wire            n29593;
wire            n29594;
wire            n29595;
wire            n29596;
wire            n29597;
wire            n29598;
wire            n29599;
wire            n29600;
wire            n29601;
wire            n29602;
wire            n29603;
wire            n29604;
wire            n29605;
wire            n29606;
wire            n29607;
wire            n29608;
wire            n29609;
wire            n29610;
wire            n29611;
wire            n29612;
wire            n29613;
wire            n29614;
wire            n29615;
wire            n29616;
wire            n29617;
wire            n29618;
wire            n29619;
wire            n29620;
wire            n29621;
wire            n29622;
wire            n29623;
wire            n29624;
wire            n29625;
wire            n29626;
wire            n29627;
wire            n29628;
wire            n29629;
wire            n29630;
wire            n29631;
wire            n29632;
wire            n29633;
wire            n29634;
wire            n29635;
wire            n29636;
wire            n29637;
wire            n29638;
wire            n29639;
wire            n29640;
wire            n29641;
wire            n29642;
wire            n29643;
wire            n29644;
wire            n29645;
wire            n29646;
wire            n29647;
wire            n29648;
wire            n29649;
wire            n29650;
wire            n29651;
wire            n29652;
wire            n29653;
wire            n29654;
wire            n29655;
wire            n29656;
wire            n29657;
wire            n29658;
wire            n29659;
wire            n29660;
wire            n29661;
wire            n29662;
wire            n29663;
wire            n29664;
wire            n29665;
wire            n29666;
wire            n29667;
wire            n29668;
wire            n29669;
wire            n29670;
wire            n29671;
wire            n29672;
wire            n29673;
wire            n29674;
wire            n29675;
wire            n29676;
wire            n29677;
wire            n29678;
wire            n29679;
wire            n29680;
wire            n29681;
wire            n29682;
wire            n29683;
wire            n29684;
wire            n29685;
wire            n29686;
wire            n29687;
wire            n29688;
wire            n29689;
wire            n29690;
wire            n29691;
wire            n29692;
wire            n29693;
wire            n29694;
wire            n29695;
wire            n29696;
wire            n29697;
wire            n29698;
wire            n29699;
wire            n29700;
wire            n29701;
wire            n29702;
wire            n29703;
wire            n29704;
wire            n29705;
wire            n29706;
wire            n29707;
wire            n29708;
wire            n29709;
wire            n29710;
wire            n29711;
wire            n29712;
wire            n29713;
wire            n29714;
wire            n29715;
wire            n29716;
wire            n29717;
wire            n29718;
wire            n29719;
wire            n29720;
wire            n29721;
wire            n29722;
wire            n29723;
wire            n29724;
wire            n29725;
wire            n29726;
wire            n29727;
wire            n29728;
wire            n29729;
wire            n29730;
wire            n29731;
wire            n29732;
wire            n29733;
wire            n29734;
wire            n29735;
wire            n29736;
wire            n29737;
wire            n29738;
wire            n29739;
wire            n29740;
wire            n29741;
wire            n29742;
wire            n29743;
wire            n29744;
wire            n29745;
wire            n29746;
wire            n29747;
wire            n29748;
wire            n29749;
wire            n29750;
wire            n29751;
wire            n29752;
wire            n29753;
wire            n29754;
wire            n29755;
wire            n29756;
wire            n29757;
wire            n29758;
wire            n29759;
wire            n29760;
wire            n29761;
wire            n29762;
wire            n29763;
wire            n29764;
wire            n29765;
wire            n29766;
wire            n29767;
wire            n29768;
wire            n29769;
wire            n29770;
wire            n29771;
wire            n29772;
wire            n29773;
wire            n29774;
wire            n29775;
wire            n29776;
wire            n29777;
wire            n29778;
wire            n29779;
wire            n29780;
wire            n29781;
wire            n29782;
wire            n29783;
wire            n29784;
wire            n29785;
wire            n29786;
wire            n29787;
wire            n29788;
wire            n29789;
wire            n29790;
wire            n29791;
wire            n29792;
wire            n29793;
wire            n29794;
wire            n29795;
wire            n29796;
wire            n29797;
wire            n29798;
wire            n29799;
wire            n29800;
wire            n29801;
wire            n29802;
wire            n29803;
wire            n29804;
wire            n29805;
wire            n29806;
wire            n29807;
wire            n29808;
wire            n29809;
wire            n29810;
wire            n29811;
wire            n29812;
wire            n29813;
wire            n29814;
wire            n29815;
wire            n29816;
wire            n29817;
wire            n29818;
wire            n29819;
wire            n29820;
wire            n29821;
wire            n29822;
wire            n29823;
wire            n29824;
wire            n29825;
wire            n29826;
wire            n29827;
wire            n29828;
wire            n29829;
wire            n29830;
wire            n29831;
wire            n29832;
wire            n29833;
wire            n29834;
wire            n29835;
wire            n29836;
wire            n29837;
wire            n29838;
wire            n29839;
wire            n29840;
wire            n29841;
wire            n29842;
wire            n29843;
wire            n29844;
wire            n29845;
wire            n29846;
wire            n29847;
wire            n29848;
wire            n29849;
wire            n29850;
wire            n29851;
wire            n29852;
wire            n29853;
wire            n29854;
wire            n29855;
wire            n29856;
wire            n29857;
wire            n29858;
wire            n29859;
wire            n29860;
wire            n29861;
wire            n29862;
wire            n29863;
wire            n29864;
wire            n29865;
wire            n29866;
wire            n29867;
wire            n29868;
wire            n29869;
wire            n29870;
wire            n29871;
wire            n29872;
wire            n29873;
wire            n29874;
wire            n29875;
wire            n29876;
wire            n29877;
wire            n29878;
wire            n29879;
wire            n29880;
wire            n29881;
wire            n29882;
wire            n29883;
wire            n29884;
wire            n29885;
wire            n29886;
wire            n29887;
wire            n29888;
wire            n29889;
wire            n29890;
wire            n29891;
wire            n29892;
wire            n29893;
wire            n29894;
wire            n29895;
wire            n29896;
wire            n29897;
wire            n29898;
wire            n29899;
wire            n29900;
wire            n29901;
wire            n29902;
wire            n29903;
wire            n29904;
wire            n29905;
wire            n29906;
wire            n29907;
wire            n29908;
wire            n29909;
wire            n29910;
wire            n29911;
wire            n29912;
wire            n29913;
wire            n29914;
wire            n29915;
wire            n29916;
wire            n29917;
wire            n29918;
wire            n29919;
wire            n29920;
wire            n29921;
wire            n29922;
wire            n29923;
wire            n29924;
wire            n29925;
wire            n29926;
wire            n29927;
wire            n29928;
wire            n29929;
wire            n29930;
wire            n29931;
wire            n29932;
wire            n29933;
wire            n29934;
wire            n29935;
wire            n29936;
wire            n29937;
wire            n29938;
wire            n29939;
wire            n29940;
wire            n29941;
wire            n29942;
wire            n29943;
wire            n29944;
wire            n29945;
wire            n29946;
wire            n29947;
wire            n29948;
wire            n29949;
wire            n29950;
wire            n29951;
wire            n29952;
wire            n29953;
wire            n29954;
wire            n29955;
wire            n29956;
wire            n29957;
wire            n29958;
wire            n29959;
wire            n29960;
wire            n29961;
wire            n29962;
wire            n29963;
wire            n29964;
wire            n29965;
wire            n29966;
wire            n29967;
wire            n29968;
wire            n29969;
wire            n29970;
wire            n29971;
wire            n29972;
wire            n29973;
wire            n29974;
wire            n29975;
wire            n29976;
wire            n29977;
wire            n29978;
wire            n29979;
wire            n29980;
wire            n29981;
wire            n29982;
wire            n29983;
wire            n29984;
wire            n29985;
wire            n29986;
wire            n29987;
wire            n29988;
wire            n29989;
wire            n29990;
wire            n29991;
wire            n29992;
wire            n29993;
wire            n29994;
wire            n29995;
wire            n29996;
wire            n29997;
wire            n29998;
wire            n29999;
wire            n30000;
wire            n30001;
wire            n30002;
wire            n30003;
wire            n30004;
wire            n30005;
wire            n30006;
wire            n30007;
wire            n30008;
wire            n30009;
wire            n30010;
wire            n30011;
wire            n30012;
wire            n30013;
wire            n30014;
wire            n30015;
wire            n30016;
wire            n30017;
wire            n30018;
wire            n30019;
wire            n30020;
wire            n30021;
wire            n30022;
wire            n30023;
wire            n30024;
wire            n30025;
wire            n30026;
wire            n30027;
wire            n30028;
wire            n30029;
wire            n30030;
wire            n30031;
wire            n30032;
wire            n30033;
wire            n30034;
wire            n30035;
wire            n30036;
wire            n30037;
wire            n30038;
wire            n30039;
wire            n30040;
wire            n30041;
wire            n30042;
wire            n30043;
wire            n30044;
wire            n30045;
wire            n30046;
wire            n30047;
wire            n30048;
wire            n30049;
wire            n30050;
wire            n30051;
wire            n30052;
wire            n30053;
wire            n30054;
wire            n30055;
wire            n30056;
wire            n30057;
wire            n30058;
wire     [31:0] n30059;
wire     [31:0] n30060;
wire     [31:0] n30061;
wire     [31:0] n30062;
wire     [31:0] n30063;
wire     [31:0] n30064;
wire     [31:0] n30065;
wire     [31:0] n30066;
wire     [31:0] n30067;
wire     [31:0] n30068;
wire     [31:0] n30069;
wire     [31:0] n30070;
wire     [31:0] n30071;
wire     [31:0] n30072;
wire     [31:0] n30073;
wire     [31:0] n30074;
wire     [31:0] n30075;
wire     [31:0] n30076;
wire     [31:0] n30077;
wire     [31:0] n30078;
wire     [31:0] n30079;
wire     [31:0] n30080;
wire     [31:0] n30081;
wire     [31:0] n30082;
wire     [31:0] n30083;
wire     [31:0] n30084;
wire     [31:0] n30085;
wire     [31:0] n30086;
wire     [31:0] n30087;
wire     [31:0] n30088;
wire     [31:0] n30089;
wire     [31:0] n30090;
wire     [31:0] n30091;
wire     [31:0] n30092;
wire     [31:0] n30093;
wire     [31:0] n30094;
wire     [31:0] n30095;
wire     [31:0] n30096;
wire     [31:0] n30097;
wire     [31:0] n30098;
wire     [31:0] n30099;
wire     [31:0] n30100;
wire     [31:0] n30101;
wire     [31:0] n30102;
wire     [31:0] n30103;
wire     [31:0] n30104;
wire     [31:0] n30105;
wire     [31:0] n30106;
wire     [31:0] n30107;
wire     [31:0] n30108;
wire     [31:0] n30109;
wire     [31:0] n30110;
wire     [31:0] n30111;
wire     [31:0] n30112;
wire     [31:0] n30113;
wire     [31:0] n30114;
wire     [31:0] n30115;
wire     [31:0] n30116;
wire     [31:0] n30117;
wire     [31:0] n30118;
wire     [31:0] n30119;
wire     [31:0] n30120;
wire     [31:0] n30121;
wire     [31:0] n30122;
wire     [31:0] n30123;
wire     [31:0] n30124;
wire     [31:0] n30125;
wire     [31:0] n30126;
wire     [31:0] n30127;
wire     [31:0] n30128;
wire     [31:0] n30129;
wire     [31:0] n30130;
wire     [31:0] n30131;
wire     [31:0] n30132;
wire     [31:0] n30133;
wire     [31:0] n30134;
wire     [31:0] n30135;
wire     [31:0] n30136;
wire     [31:0] n30137;
wire     [31:0] n30138;
wire     [31:0] n30139;
wire     [31:0] n30140;
wire     [31:0] n30141;
wire     [31:0] n30142;
wire     [31:0] n30143;
wire     [31:0] n30144;
wire     [31:0] n30145;
wire     [31:0] n30146;
wire     [31:0] n30147;
wire     [31:0] n30148;
wire     [31:0] n30149;
wire     [31:0] n30150;
wire     [31:0] n30151;
wire     [31:0] n30152;
wire     [31:0] n30153;
wire     [31:0] n30154;
wire     [31:0] n30155;
wire     [31:0] n30156;
wire     [31:0] n30157;
wire     [31:0] n30158;
wire     [31:0] n30159;
wire     [31:0] n30160;
wire     [31:0] n30161;
wire     [31:0] n30162;
wire     [31:0] n30163;
wire     [31:0] n30164;
wire     [31:0] n30165;
wire     [31:0] n30166;
wire     [31:0] n30167;
wire     [31:0] n30168;
wire     [31:0] n30169;
wire     [31:0] n30170;
wire     [31:0] n30171;
wire     [31:0] n30172;
wire     [31:0] n30173;
wire     [31:0] n30174;
wire     [31:0] n30175;
wire     [31:0] n30176;
wire     [31:0] n30177;
wire     [31:0] n30178;
wire     [31:0] n30179;
wire     [31:0] n30180;
wire     [31:0] n30181;
wire     [31:0] n30182;
wire     [31:0] n30183;
wire     [31:0] n30184;
wire     [31:0] n30185;
wire     [31:0] n30186;
wire     [31:0] n30187;
wire     [31:0] n30188;
wire     [31:0] n30189;
wire     [31:0] n30190;
wire     [31:0] n30191;
wire     [31:0] n30192;
wire     [31:0] n30193;
wire     [31:0] n30194;
wire     [31:0] n30195;
wire     [31:0] n30196;
wire     [31:0] n30197;
wire     [31:0] n30198;
wire     [31:0] n30199;
wire     [31:0] n30200;
wire     [31:0] n30201;
wire     [31:0] n30202;
wire     [31:0] n30203;
wire     [31:0] n30204;
wire     [31:0] n30205;
wire     [31:0] n30206;
wire     [31:0] n30207;
wire     [31:0] n30208;
wire     [31:0] n30209;
wire     [31:0] n30210;
wire     [31:0] n30211;
wire     [31:0] n30212;
wire     [31:0] n30213;
wire     [31:0] n30214;
wire     [31:0] n30215;
wire     [31:0] n30216;
wire     [31:0] n30217;
wire     [31:0] n30218;
wire     [31:0] n30219;
wire     [31:0] n30220;
wire     [31:0] n30221;
wire     [31:0] n30222;
wire     [31:0] n30223;
wire     [31:0] n30224;
wire     [31:0] n30225;
wire     [31:0] n30226;
wire     [31:0] n30227;
wire     [31:0] n30228;
wire     [31:0] n30229;
wire     [31:0] n30230;
wire     [31:0] n30231;
wire     [31:0] n30232;
wire     [31:0] n30233;
wire     [31:0] n30234;
wire     [31:0] n30235;
wire     [31:0] n30236;
wire     [31:0] n30237;
wire     [31:0] n30238;
wire     [31:0] n30239;
wire     [31:0] n30240;
wire     [31:0] n30241;
wire     [31:0] n30242;
wire     [31:0] n30243;
wire     [31:0] n30244;
wire     [31:0] n30245;
wire     [31:0] n30246;
wire     [31:0] n30247;
wire     [31:0] n30248;
wire     [31:0] n30249;
wire     [31:0] n30250;
wire     [31:0] n30251;
wire     [31:0] n30252;
wire     [31:0] n30253;
wire     [31:0] n30254;
wire     [31:0] n30255;
wire     [31:0] n30256;
wire     [31:0] n30257;
wire     [31:0] n30258;
wire     [31:0] n30259;
wire     [31:0] n30260;
wire     [31:0] n30261;
wire     [31:0] n30262;
wire     [31:0] n30263;
wire     [31:0] n30264;
wire     [31:0] n30265;
wire     [31:0] n30266;
wire     [31:0] n30267;
wire     [31:0] n30268;
wire     [31:0] n30269;
wire     [31:0] n30270;
wire     [31:0] n30271;
wire     [31:0] n30272;
wire     [31:0] n30273;
wire     [31:0] n30274;
wire     [31:0] n30275;
wire     [31:0] n30276;
wire     [31:0] n30277;
wire     [31:0] n30278;
wire     [31:0] n30279;
wire     [31:0] n30280;
wire     [31:0] n30281;
wire     [31:0] n30282;
wire     [31:0] n30283;
wire     [31:0] n30284;
wire     [31:0] n30285;
wire     [31:0] n30286;
wire     [31:0] n30287;
wire     [31:0] n30288;
wire     [31:0] n30289;
wire     [31:0] n30290;
wire     [31:0] n30291;
wire     [31:0] n30292;
wire     [31:0] n30293;
wire     [31:0] n30294;
wire     [31:0] n30295;
wire     [31:0] n30296;
wire     [31:0] n30297;
wire     [31:0] n30298;
wire     [31:0] n30299;
wire     [31:0] n30300;
wire     [31:0] n30301;
wire     [31:0] n30302;
wire     [31:0] n30303;
wire     [31:0] n30304;
wire     [31:0] n30305;
wire     [31:0] n30306;
wire     [31:0] n30307;
wire     [31:0] n30308;
wire     [31:0] n30309;
wire     [31:0] n30310;
wire     [31:0] n30311;
wire     [31:0] n30312;
wire     [31:0] n30313;
wire     [31:0] n30314;
wire     [31:0] n30315;
wire     [31:0] n30316;
wire     [31:0] n30317;
wire     [31:0] n30318;
wire     [31:0] n30319;
wire     [31:0] n30320;
wire     [31:0] n30321;
wire     [31:0] n30322;
wire     [31:0] n30323;
wire     [31:0] n30324;
wire     [31:0] n30325;
wire     [31:0] n30326;
wire     [31:0] n30327;
wire     [31:0] n30328;
wire     [31:0] n30329;
wire     [31:0] n30330;
wire     [31:0] n30331;
wire     [31:0] n30332;
wire     [31:0] n30333;
wire     [31:0] n30334;
wire     [31:0] n30335;
wire     [31:0] n30336;
wire     [31:0] n30337;
wire     [31:0] n30338;
wire     [31:0] n30339;
wire     [31:0] n30340;
wire     [31:0] n30341;
wire     [31:0] n30342;
wire     [31:0] n30343;
wire     [31:0] n30344;
wire     [31:0] n30345;
wire     [31:0] n30346;
wire     [31:0] n30347;
wire     [31:0] n30348;
wire     [31:0] n30349;
wire     [31:0] n30350;
wire     [31:0] n30351;
wire     [31:0] n30352;
wire     [31:0] n30353;
wire     [31:0] n30354;
wire     [31:0] n30355;
wire     [31:0] n30356;
wire     [31:0] n30357;
wire     [31:0] n30358;
wire     [31:0] n30359;
wire     [31:0] n30360;
wire     [31:0] n30361;
wire     [31:0] n30362;
wire     [31:0] n30363;
wire     [31:0] n30364;
wire     [31:0] n30365;
wire     [31:0] n30366;
wire     [31:0] n30367;
wire     [31:0] n30368;
wire     [31:0] n30369;
wire     [31:0] n30370;
wire     [31:0] n30371;
wire     [31:0] n30372;
wire     [31:0] n30373;
wire     [31:0] n30374;
wire     [31:0] n30375;
wire     [31:0] n30376;
wire     [31:0] n30377;
wire     [31:0] n30378;
wire     [31:0] n30379;
wire     [31:0] n30380;
wire     [31:0] n30381;
wire     [31:0] n30382;
wire     [31:0] n30383;
wire     [31:0] n30384;
wire     [31:0] n30385;
wire     [31:0] n30386;
wire     [31:0] n30387;
wire     [31:0] n30388;
wire     [31:0] n30389;
wire     [31:0] n30390;
wire     [31:0] n30391;
wire     [31:0] n30392;
wire     [31:0] n30393;
wire     [31:0] n30394;
wire     [31:0] n30395;
wire     [31:0] n30396;
wire     [31:0] n30397;
wire     [31:0] n30398;
wire     [31:0] n30399;
wire     [31:0] n30400;
wire     [31:0] n30401;
wire     [31:0] n30402;
wire     [31:0] n30403;
wire     [31:0] n30404;
wire     [31:0] n30405;
wire     [31:0] n30406;
wire     [31:0] n30407;
wire     [31:0] n30408;
wire     [31:0] n30409;
wire     [31:0] n30410;
wire     [31:0] n30411;
wire     [31:0] n30412;
wire     [31:0] n30413;
wire     [31:0] n30414;
wire     [31:0] n30415;
wire     [31:0] n30416;
wire     [31:0] n30417;
wire     [31:0] n30418;
wire     [31:0] n30419;
wire     [31:0] n30420;
wire     [31:0] n30421;
wire     [31:0] n30422;
wire     [31:0] n30423;
wire     [31:0] n30424;
wire     [31:0] n30425;
wire     [31:0] n30426;
wire     [31:0] n30427;
wire     [31:0] n30428;
wire     [31:0] n30429;
wire     [31:0] n30430;
wire     [31:0] n30431;
wire     [31:0] n30432;
wire     [31:0] n30433;
wire     [31:0] n30434;
wire     [31:0] n30435;
wire     [31:0] n30436;
wire     [31:0] n30437;
wire     [31:0] n30438;
wire     [31:0] n30439;
wire     [31:0] n30440;
wire     [31:0] n30441;
wire     [31:0] n30442;
wire     [31:0] n30443;
wire     [31:0] n30444;
wire     [31:0] n30445;
wire     [31:0] n30446;
wire     [31:0] n30447;
wire     [31:0] n30448;
wire     [31:0] n30449;
wire     [31:0] n30450;
wire     [31:0] n30451;
wire     [31:0] n30452;
wire     [31:0] n30453;
wire     [31:0] n30454;
wire     [31:0] n30455;
wire     [31:0] n30456;
wire     [31:0] n30457;
wire     [31:0] n30458;
wire     [31:0] n30459;
wire     [31:0] n30460;
wire     [31:0] n30461;
wire     [31:0] n30462;
wire     [31:0] n30463;
wire     [31:0] n30464;
wire     [31:0] n30465;
wire     [31:0] n30466;
wire     [31:0] n30467;
wire     [31:0] n30468;
wire     [31:0] n30469;
wire     [31:0] n30470;
wire     [31:0] n30471;
wire     [31:0] n30472;
wire     [31:0] n30473;
wire     [31:0] n30474;
wire     [31:0] n30475;
wire     [31:0] n30476;
wire     [31:0] n30477;
wire     [31:0] n30478;
wire     [31:0] n30479;
wire     [31:0] n30480;
wire     [31:0] n30481;
wire     [31:0] n30482;
wire     [31:0] n30483;
wire     [31:0] n30484;
wire     [31:0] n30485;
wire     [31:0] n30486;
wire     [31:0] n30487;
wire     [31:0] n30488;
wire     [31:0] n30489;
wire     [31:0] n30490;
wire     [31:0] n30491;
wire     [31:0] n30492;
wire     [31:0] n30493;
wire     [31:0] n30494;
wire     [31:0] n30495;
wire     [31:0] n30496;
wire     [31:0] n30497;
wire     [31:0] n30498;
wire     [31:0] n30499;
wire     [31:0] n30500;
wire     [31:0] n30501;
wire     [31:0] n30502;
wire     [31:0] n30503;
wire     [31:0] n30504;
wire     [31:0] n30505;
wire     [31:0] n30506;
wire     [31:0] n30507;
wire     [31:0] n30508;
wire     [31:0] n30509;
wire     [31:0] n30510;
wire     [31:0] n30511;
wire     [31:0] n30512;
wire     [31:0] n30513;
wire     [31:0] n30514;
wire     [31:0] n30515;
wire     [31:0] n30516;
wire     [31:0] n30517;
wire     [31:0] n30518;
wire     [31:0] n30519;
wire     [31:0] n30520;
wire     [31:0] n30521;
wire     [31:0] n30522;
wire     [31:0] n30523;
wire     [31:0] n30524;
wire     [31:0] n30525;
wire     [31:0] n30526;
wire     [31:0] n30527;
wire     [31:0] n30528;
wire     [31:0] n30529;
wire     [31:0] n30530;
wire     [31:0] n30531;
wire     [31:0] n30532;
wire     [31:0] n30533;
wire     [31:0] n30534;
wire     [31:0] n30535;
wire     [31:0] n30536;
wire     [31:0] n30537;
wire     [31:0] n30538;
wire     [31:0] n30539;
wire     [31:0] n30540;
wire     [31:0] n30541;
wire     [31:0] n30542;
wire     [31:0] n30543;
wire     [31:0] n30544;
wire     [31:0] n30545;
wire     [31:0] n30546;
wire     [31:0] n30547;
wire     [31:0] n30548;
wire     [31:0] n30549;
wire     [31:0] n30550;
wire     [31:0] n30551;
wire     [31:0] n30552;
wire     [31:0] n30553;
wire     [31:0] n30554;
wire     [31:0] n30555;
wire     [31:0] n30556;
wire     [31:0] n30557;
wire     [31:0] n30558;
wire     [31:0] n30559;
wire     [31:0] n30560;
wire     [31:0] n30561;
wire     [31:0] n30562;
wire     [31:0] n30563;
wire     [31:0] n30564;
wire     [31:0] n30565;
wire     [31:0] n30566;
wire     [31:0] n30567;
wire     [31:0] n30568;
wire     [31:0] n30569;
wire     [31:0] n30570;
wire     [31:0] n30571;
wire     [31:0] n30572;
wire     [31:0] n30573;
wire     [31:0] n30574;
wire     [31:0] n30575;
wire     [31:0] n30576;
wire     [31:0] n30577;
wire     [31:0] n30578;
wire     [31:0] n30579;
wire     [31:0] n30580;
wire            n30581;
wire            n30582;
wire     [31:0] n30583;
wire     [31:0] n30584;
wire     [31:0] n30585;
wire     [31:0] n30586;
wire     [31:0] n30587;
wire     [31:0] n30588;
wire     [31:0] n30589;
wire     [31:0] n30590;
wire     [31:0] n30591;
wire     [31:0] n30592;
wire     [31:0] n30593;
wire     [31:0] n30594;
wire     [31:0] n30595;
wire     [31:0] n30596;
wire     [31:0] n30597;
wire     [31:0] n30598;
wire     [31:0] n30599;
wire     [31:0] n30600;
wire     [31:0] n30601;
wire     [31:0] n30602;
wire     [31:0] n30603;
wire     [31:0] n30604;
wire     [31:0] n30605;
wire     [31:0] n30606;
wire     [31:0] n30607;
wire     [31:0] n30608;
wire     [31:0] n30609;
wire     [31:0] n30610;
wire     [31:0] n30611;
wire     [31:0] n30612;
wire     [31:0] n30613;
wire     [31:0] n30614;
wire     [31:0] n30615;
wire            n30616;
wire            n30617;
wire            n30618;
wire            n30619;
wire            n30620;
wire            n30621;
wire            n30622;
wire            n30623;
wire            n30624;
wire            n30625;
wire            n30626;
wire            n30627;
wire            n30628;
wire            n30629;
wire            n30630;
wire            n30631;
wire            n30632;
wire            n30633;
wire            n30634;
wire            n30635;
wire            n30636;
wire            n30637;
wire            n30638;
wire            n30639;
wire            n30640;
wire            n30641;
wire            n30642;
wire            n30643;
wire            n30644;
wire            n30645;
wire            n30646;
wire            n30647;
wire            n30648;
wire            n30649;
wire            n30650;
wire            n30651;
wire            n30652;
wire            n30653;
wire            n30654;
wire            n30655;
wire            n30656;
wire            n30657;
wire            n30658;
wire            n30659;
wire            n30660;
wire            n30661;
wire            n30662;
wire            n30663;
wire            n30664;
wire            n30665;
wire            n30666;
wire            n30667;
wire            n30668;
wire            n30669;
wire            n30670;
wire            n30671;
wire            n30672;
wire            n30673;
wire            n30674;
wire            n30675;
wire            n30676;
wire            n30677;
wire            n30678;
wire            n30679;
wire            n30680;
wire            n30681;
wire            n30682;
wire            n30683;
wire            n30684;
wire            n30685;
wire            n30686;
wire            n30687;
wire            n30688;
wire            n30689;
wire            n30690;
wire            n30691;
wire            n30692;
wire            n30693;
wire            n30694;
wire            n30695;
wire            n30696;
wire            n30697;
wire            n30698;
wire            n30699;
wire            n30700;
wire            n30701;
wire            n30702;
wire            n30703;
wire            n30704;
wire            n30705;
wire            n30706;
wire            n30707;
wire            n30708;
wire            n30709;
wire            n30710;
wire            n30711;
wire            n30712;
wire            n30713;
wire            n30714;
wire            n30715;
wire            n30716;
wire            n30717;
wire            n30718;
wire            n30719;
wire            n30720;
wire            n30721;
wire            n30722;
wire            n30723;
wire            n30724;
wire            n30725;
wire            n30726;
wire            n30727;
wire            n30728;
wire            n30729;
wire            n30730;
wire            n30731;
wire            n30732;
wire            n30733;
wire            n30734;
wire            n30735;
wire            n30736;
wire            n30737;
wire            n30738;
wire            n30739;
wire            n30740;
wire            n30741;
wire            n30742;
wire            n30743;
wire            n30744;
wire            n30745;
wire            n30746;
wire            n30747;
wire            n30748;
wire            n30749;
wire            n30750;
wire            n30751;
wire            n30752;
wire            n30753;
wire            n30754;
wire            n30755;
wire            n30756;
wire            n30757;
wire            n30758;
wire            n30759;
wire            n30760;
wire            n30761;
wire            n30762;
wire            n30763;
wire            n30764;
wire            n30765;
wire            n30766;
wire            n30767;
wire            n30768;
wire            n30769;
wire            n30770;
wire            n30771;
wire            n30772;
wire            n30773;
wire            n30774;
wire            n30775;
wire            n30776;
wire            n30777;
wire            n30778;
wire            n30779;
wire            n30780;
wire            n30781;
wire            n30782;
wire            n30783;
wire            n30784;
wire            n30785;
wire            n30786;
wire            n30787;
wire            n30788;
wire            n30789;
wire            n30790;
wire            n30791;
wire            n30792;
wire            n30793;
wire            n30794;
wire            n30795;
wire            n30796;
wire            n30797;
wire            n30798;
wire            n30799;
wire            n30800;
wire            n30801;
wire            n30802;
wire            n30803;
wire            n30804;
wire            n30805;
wire            n30806;
wire            n30807;
wire            n30808;
wire            n30809;
wire            n30810;
wire            n30811;
wire            n30812;
wire            n30813;
wire            n30814;
wire            n30815;
wire            n30816;
wire            n30817;
wire            n30818;
wire            n30819;
wire            n30820;
wire            n30821;
wire            n30822;
wire            n30823;
wire            n30824;
wire            n30825;
wire            n30826;
wire            n30827;
wire            n30828;
wire            n30829;
wire            n30830;
wire            n30831;
wire            n30832;
wire            n30833;
wire            n30834;
wire            n30835;
wire            n30836;
wire            n30837;
wire            n30838;
wire            n30839;
wire            n30840;
wire            n30841;
wire            n30842;
wire            n30843;
wire            n30844;
wire            n30845;
wire            n30846;
wire            n30847;
wire            n30848;
wire            n30849;
wire            n30850;
wire            n30851;
wire            n30852;
wire            n30853;
wire            n30854;
wire            n30855;
wire            n30856;
wire            n30857;
wire            n30858;
wire            n30859;
wire            n30860;
wire            n30861;
wire            n30862;
wire            n30863;
wire            n30864;
wire            n30865;
wire            n30866;
wire            n30867;
wire            n30868;
wire            n30869;
wire            n30870;
wire            n30871;
wire            n30872;
wire            n30873;
wire            n30874;
wire            n30875;
wire            n30876;
wire            n30877;
wire            n30878;
wire            n30879;
wire            n30880;
wire            n30881;
wire            n30882;
wire            n30883;
wire            n30884;
wire            n30885;
wire            n30886;
wire            n30887;
wire            n30888;
wire            n30889;
wire            n30890;
wire            n30891;
wire            n30892;
wire            n30893;
wire            n30894;
wire            n30895;
wire            n30896;
wire            n30897;
wire            n30898;
wire            n30899;
wire            n30900;
wire            n30901;
wire            n30902;
wire            n30903;
wire            n30904;
wire            n30905;
wire            n30906;
wire            n30907;
wire            n30908;
wire            n30909;
wire            n30910;
wire            n30911;
wire            n30912;
wire            n30913;
wire            n30914;
wire            n30915;
wire            n30916;
wire            n30917;
wire            n30918;
wire            n30919;
wire            n30920;
wire            n30921;
wire            n30922;
wire            n30923;
wire            n30924;
wire            n30925;
wire            n30926;
wire            n30927;
wire            n30928;
wire            n30929;
wire            n30930;
wire            n30931;
wire            n30932;
wire            n30933;
wire            n30934;
wire            n30935;
wire            n30936;
wire            n30937;
wire            n30938;
wire            n30939;
wire            n30940;
wire            n30941;
wire            n30942;
wire            n30943;
wire            n30944;
wire            n30945;
wire            n30946;
wire            n30947;
wire            n30948;
wire            n30949;
wire            n30950;
wire            n30951;
wire            n30952;
wire            n30953;
wire            n30954;
wire            n30955;
wire            n30956;
wire            n30957;
wire            n30958;
wire            n30959;
wire            n30960;
wire            n30961;
wire            n30962;
wire            n30963;
wire            n30964;
wire            n30965;
wire            n30966;
wire            n30967;
wire            n30968;
wire            n30969;
wire            n30970;
wire            n30971;
wire            n30972;
wire            n30973;
wire            n30974;
wire            n30975;
wire            n30976;
wire            n30977;
wire            n30978;
wire            n30979;
wire            n30980;
wire            n30981;
wire            n30982;
wire            n30983;
wire            n30984;
wire            n30985;
wire            n30986;
wire            n30987;
wire            n30988;
wire            n30989;
wire            n30990;
wire            n30991;
wire            n30992;
wire            n30993;
wire            n30994;
wire            n30995;
wire            n30996;
wire            n30997;
wire            n30998;
wire            n30999;
wire            n31000;
wire            n31001;
wire            n31002;
wire            n31003;
wire            n31004;
wire            n31005;
wire            n31006;
wire            n31007;
wire            n31008;
wire            n31009;
wire            n31010;
wire            n31011;
wire            n31012;
wire            n31013;
wire            n31014;
wire            n31015;
wire            n31016;
wire            n31017;
wire            n31018;
wire            n31019;
wire            n31020;
wire            n31021;
wire            n31022;
wire            n31023;
wire            n31024;
wire            n31025;
wire            n31026;
wire            n31027;
wire            n31028;
wire            n31029;
wire            n31030;
wire            n31031;
wire            n31032;
wire            n31033;
wire            n31034;
wire            n31035;
wire            n31036;
wire            n31037;
wire            n31038;
wire            n31039;
wire            n31040;
wire            n31041;
wire            n31042;
wire            n31043;
wire            n31044;
wire            n31045;
wire            n31046;
wire            n31047;
wire            n31048;
wire            n31049;
wire            n31050;
wire            n31051;
wire            n31052;
wire            n31053;
wire            n31054;
wire            n31055;
wire            n31056;
wire            n31057;
wire            n31058;
wire            n31059;
wire            n31060;
wire            n31061;
wire            n31062;
wire            n31063;
wire            n31064;
wire            n31065;
wire            n31066;
wire            n31067;
wire            n31068;
wire            n31069;
wire            n31070;
wire            n31071;
wire            n31072;
wire            n31073;
wire            n31074;
wire            n31075;
wire            n31076;
wire            n31077;
wire            n31078;
wire            n31079;
wire            n31080;
wire            n31081;
wire            n31082;
wire            n31083;
wire            n31084;
wire            n31085;
wire            n31086;
wire            n31087;
wire            n31088;
wire            n31089;
wire            n31090;
wire            n31091;
wire            n31092;
wire            n31093;
wire            n31094;
wire            n31095;
wire            n31096;
wire            n31097;
wire            n31098;
wire            n31099;
wire            n31100;
wire            n31101;
wire            n31102;
wire            n31103;
wire            n31104;
wire            n31105;
wire            n31106;
wire            n31107;
wire            n31108;
wire            n31109;
wire            n31110;
wire            n31111;
wire            n31112;
wire            n31113;
wire            n31114;
wire            n31115;
wire            n31116;
wire            n31117;
wire            n31118;
wire            n31119;
wire            n31120;
wire            n31121;
wire            n31122;
wire            n31123;
wire            n31124;
wire            n31125;
wire            n31126;
wire            n31127;
wire            n31128;
wire            n31129;
wire            n31130;
wire            n31131;
wire            n31132;
wire            n31133;
wire            n31134;
wire            n31135;
wire            n31136;
wire            n31137;
wire            n31138;
wire            n31139;
wire            n31140;
wire            n31141;
wire            n31142;
wire            n31143;
wire     [31:0] n31144;
wire     [31:0] n31145;
wire     [31:0] n31146;
wire     [31:0] n31147;
wire     [31:0] n31148;
wire     [31:0] n31149;
wire     [31:0] n31150;
wire     [31:0] n31151;
wire     [31:0] n31152;
wire     [31:0] n31153;
wire     [31:0] n31154;
wire     [31:0] n31155;
wire     [31:0] n31156;
wire     [31:0] n31157;
wire     [31:0] n31158;
wire     [31:0] n31159;
wire     [31:0] n31160;
wire     [31:0] n31161;
wire     [31:0] n31162;
wire     [31:0] n31163;
wire     [31:0] n31164;
wire     [31:0] n31165;
wire     [31:0] n31166;
wire     [31:0] n31167;
wire     [31:0] n31168;
wire     [31:0] n31169;
wire     [31:0] n31170;
wire     [31:0] n31171;
wire     [31:0] n31172;
wire     [31:0] n31173;
wire     [31:0] n31174;
wire     [31:0] n31175;
wire     [31:0] n31176;
wire     [31:0] n31177;
wire     [31:0] n31178;
wire     [31:0] n31179;
wire     [31:0] n31180;
wire     [31:0] n31181;
wire     [31:0] n31182;
wire     [31:0] n31183;
wire     [31:0] n31184;
wire     [31:0] n31185;
wire     [31:0] n31186;
wire     [31:0] n31187;
wire     [31:0] n31188;
wire     [31:0] n31189;
wire     [31:0] n31190;
wire     [31:0] n31191;
wire     [31:0] n31192;
wire     [31:0] n31193;
wire     [31:0] n31194;
wire     [31:0] n31195;
wire     [31:0] n31196;
wire     [31:0] n31197;
wire     [31:0] n31198;
wire     [31:0] n31199;
wire     [31:0] n31200;
wire     [31:0] n31201;
wire     [31:0] n31202;
wire     [31:0] n31203;
wire     [31:0] n31204;
wire     [31:0] n31205;
wire     [31:0] n31206;
wire     [31:0] n31207;
wire     [31:0] n31208;
wire     [31:0] n31209;
wire     [31:0] n31210;
wire     [31:0] n31211;
wire     [31:0] n31212;
wire     [31:0] n31213;
wire     [31:0] n31214;
wire     [31:0] n31215;
wire     [31:0] n31216;
wire     [31:0] n31217;
wire     [31:0] n31218;
wire     [31:0] n31219;
wire     [31:0] n31220;
wire     [31:0] n31221;
wire     [31:0] n31222;
wire     [31:0] n31223;
wire     [31:0] n31224;
wire     [31:0] n31225;
wire     [31:0] n31226;
wire     [31:0] n31227;
wire     [31:0] n31228;
wire     [31:0] n31229;
wire     [31:0] n31230;
wire     [31:0] n31231;
wire     [31:0] n31232;
wire     [31:0] n31233;
wire     [31:0] n31234;
wire     [31:0] n31235;
wire     [31:0] n31236;
wire     [31:0] n31237;
wire     [31:0] n31238;
wire     [31:0] n31239;
wire     [31:0] n31240;
wire     [31:0] n31241;
wire     [31:0] n31242;
wire     [31:0] n31243;
wire     [31:0] n31244;
wire     [31:0] n31245;
wire     [31:0] n31246;
wire     [31:0] n31247;
wire     [31:0] n31248;
wire     [31:0] n31249;
wire     [31:0] n31250;
wire     [31:0] n31251;
wire     [31:0] n31252;
wire     [31:0] n31253;
wire     [31:0] n31254;
wire     [31:0] n31255;
wire     [31:0] n31256;
wire     [31:0] n31257;
wire     [31:0] n31258;
wire     [31:0] n31259;
wire     [31:0] n31260;
wire     [31:0] n31261;
wire     [31:0] n31262;
wire     [31:0] n31263;
wire     [31:0] n31264;
wire     [31:0] n31265;
wire     [31:0] n31266;
wire     [31:0] n31267;
wire     [31:0] n31268;
wire     [31:0] n31269;
wire     [31:0] n31270;
wire     [31:0] n31271;
wire     [31:0] n31272;
wire     [31:0] n31273;
wire     [31:0] n31274;
wire     [31:0] n31275;
wire     [31:0] n31276;
wire     [31:0] n31277;
wire     [31:0] n31278;
wire     [31:0] n31279;
wire     [31:0] n31280;
wire     [31:0] n31281;
wire     [31:0] n31282;
wire     [31:0] n31283;
wire     [31:0] n31284;
wire     [31:0] n31285;
wire     [31:0] n31286;
wire     [31:0] n31287;
wire     [31:0] n31288;
wire     [31:0] n31289;
wire     [31:0] n31290;
wire     [31:0] n31291;
wire     [31:0] n31292;
wire     [31:0] n31293;
wire     [31:0] n31294;
wire     [31:0] n31295;
wire     [31:0] n31296;
wire     [31:0] n31297;
wire     [31:0] n31298;
wire     [31:0] n31299;
wire     [31:0] n31300;
wire     [31:0] n31301;
wire     [31:0] n31302;
wire     [31:0] n31303;
wire     [31:0] n31304;
wire     [31:0] n31305;
wire     [31:0] n31306;
wire     [31:0] n31307;
wire     [31:0] n31308;
wire     [31:0] n31309;
wire     [31:0] n31310;
wire     [31:0] n31311;
wire     [31:0] n31312;
wire     [31:0] n31313;
wire     [31:0] n31314;
wire     [31:0] n31315;
wire     [31:0] n31316;
wire     [31:0] n31317;
wire     [31:0] n31318;
wire     [31:0] n31319;
wire     [31:0] n31320;
wire     [31:0] n31321;
wire     [31:0] n31322;
wire     [31:0] n31323;
wire     [31:0] n31324;
wire     [31:0] n31325;
wire     [31:0] n31326;
wire     [31:0] n31327;
wire     [31:0] n31328;
wire     [31:0] n31329;
wire     [31:0] n31330;
wire     [31:0] n31331;
wire     [31:0] n31332;
wire     [31:0] n31333;
wire     [31:0] n31334;
wire     [31:0] n31335;
wire     [31:0] n31336;
wire     [31:0] n31337;
wire     [31:0] n31338;
wire     [31:0] n31339;
wire     [31:0] n31340;
wire     [31:0] n31341;
wire     [31:0] n31342;
wire     [31:0] n31343;
wire     [31:0] n31344;
wire     [31:0] n31345;
wire     [31:0] n31346;
wire     [31:0] n31347;
wire     [31:0] n31348;
wire     [31:0] n31349;
wire     [31:0] n31350;
wire     [31:0] n31351;
wire     [31:0] n31352;
wire     [31:0] n31353;
wire     [31:0] n31354;
wire     [31:0] n31355;
wire     [31:0] n31356;
wire     [31:0] n31357;
wire     [31:0] n31358;
wire     [31:0] n31359;
wire     [31:0] n31360;
wire     [31:0] n31361;
wire     [31:0] n31362;
wire     [31:0] n31363;
wire     [31:0] n31364;
wire     [31:0] n31365;
wire     [31:0] n31366;
wire     [31:0] n31367;
wire     [31:0] n31368;
wire     [31:0] n31369;
wire     [31:0] n31370;
wire     [31:0] n31371;
wire     [31:0] n31372;
wire     [31:0] n31373;
wire     [31:0] n31374;
wire     [31:0] n31375;
wire     [31:0] n31376;
wire     [31:0] n31377;
wire     [31:0] n31378;
wire     [31:0] n31379;
wire     [31:0] n31380;
wire     [31:0] n31381;
wire     [31:0] n31382;
wire     [31:0] n31383;
wire     [31:0] n31384;
wire     [31:0] n31385;
wire     [31:0] n31386;
wire     [31:0] n31387;
wire     [31:0] n31388;
wire     [31:0] n31389;
wire     [31:0] n31390;
wire     [31:0] n31391;
wire     [31:0] n31392;
wire     [31:0] n31393;
wire     [31:0] n31394;
wire     [31:0] n31395;
wire     [31:0] n31396;
wire     [31:0] n31397;
wire     [31:0] n31398;
wire     [31:0] n31399;
wire     [31:0] n31400;
wire     [31:0] n31401;
wire     [31:0] n31402;
wire     [31:0] n31403;
wire     [31:0] n31404;
wire     [31:0] n31405;
wire     [31:0] n31406;
wire     [31:0] n31407;
wire     [31:0] n31408;
wire     [31:0] n31409;
wire     [31:0] n31410;
wire     [31:0] n31411;
wire     [31:0] n31412;
wire     [31:0] n31413;
wire     [31:0] n31414;
wire     [31:0] n31415;
wire     [31:0] n31416;
wire     [31:0] n31417;
wire     [31:0] n31418;
wire     [31:0] n31419;
wire     [31:0] n31420;
wire     [31:0] n31421;
wire     [31:0] n31422;
wire     [31:0] n31423;
wire     [31:0] n31424;
wire     [31:0] n31425;
wire     [31:0] n31426;
wire     [31:0] n31427;
wire     [31:0] n31428;
wire     [31:0] n31429;
wire     [31:0] n31430;
wire     [31:0] n31431;
wire     [31:0] n31432;
wire     [31:0] n31433;
wire     [31:0] n31434;
wire     [31:0] n31435;
wire     [31:0] n31436;
wire     [31:0] n31437;
wire     [31:0] n31438;
wire     [31:0] n31439;
wire     [31:0] n31440;
wire     [31:0] n31441;
wire     [31:0] n31442;
wire     [31:0] n31443;
wire     [31:0] n31444;
wire     [31:0] n31445;
wire     [31:0] n31446;
wire     [31:0] n31447;
wire     [31:0] n31448;
wire     [31:0] n31449;
wire     [31:0] n31450;
wire     [31:0] n31451;
wire     [31:0] n31452;
wire     [31:0] n31453;
wire     [31:0] n31454;
wire     [31:0] n31455;
wire     [31:0] n31456;
wire     [31:0] n31457;
wire     [31:0] n31458;
wire     [31:0] n31459;
wire     [31:0] n31460;
wire     [31:0] n31461;
wire     [31:0] n31462;
wire     [31:0] n31463;
wire     [31:0] n31464;
wire     [31:0] n31465;
wire     [31:0] n31466;
wire     [31:0] n31467;
wire     [31:0] n31468;
wire     [31:0] n31469;
wire     [31:0] n31470;
wire     [31:0] n31471;
wire     [31:0] n31472;
wire     [31:0] n31473;
wire     [31:0] n31474;
wire     [31:0] n31475;
wire     [31:0] n31476;
wire     [31:0] n31477;
wire     [31:0] n31478;
wire     [31:0] n31479;
wire     [31:0] n31480;
wire     [31:0] n31481;
wire     [31:0] n31482;
wire     [31:0] n31483;
wire     [31:0] n31484;
wire     [31:0] n31485;
wire     [31:0] n31486;
wire     [31:0] n31487;
wire     [31:0] n31488;
wire     [31:0] n31489;
wire     [31:0] n31490;
wire     [31:0] n31491;
wire     [31:0] n31492;
wire     [31:0] n31493;
wire     [31:0] n31494;
wire     [31:0] n31495;
wire     [31:0] n31496;
wire     [31:0] n31497;
wire     [31:0] n31498;
wire     [31:0] n31499;
wire     [31:0] n31500;
wire     [31:0] n31501;
wire     [31:0] n31502;
wire     [31:0] n31503;
wire     [31:0] n31504;
wire     [31:0] n31505;
wire     [31:0] n31506;
wire     [31:0] n31507;
wire     [31:0] n31508;
wire     [31:0] n31509;
wire     [31:0] n31510;
wire     [31:0] n31511;
wire     [31:0] n31512;
wire     [31:0] n31513;
wire     [31:0] n31514;
wire     [31:0] n31515;
wire     [31:0] n31516;
wire     [31:0] n31517;
wire     [31:0] n31518;
wire     [31:0] n31519;
wire     [31:0] n31520;
wire     [31:0] n31521;
wire     [31:0] n31522;
wire     [31:0] n31523;
wire     [31:0] n31524;
wire     [31:0] n31525;
wire     [31:0] n31526;
wire     [31:0] n31527;
wire     [31:0] n31528;
wire     [31:0] n31529;
wire     [31:0] n31530;
wire     [31:0] n31531;
wire     [31:0] n31532;
wire     [31:0] n31533;
wire     [31:0] n31534;
wire     [31:0] n31535;
wire     [31:0] n31536;
wire     [31:0] n31537;
wire     [31:0] n31538;
wire     [31:0] n31539;
wire     [31:0] n31540;
wire     [31:0] n31541;
wire     [31:0] n31542;
wire     [31:0] n31543;
wire     [31:0] n31544;
wire     [31:0] n31545;
wire     [31:0] n31546;
wire     [31:0] n31547;
wire     [31:0] n31548;
wire     [31:0] n31549;
wire     [31:0] n31550;
wire     [31:0] n31551;
wire     [31:0] n31552;
wire     [31:0] n31553;
wire     [31:0] n31554;
wire     [31:0] n31555;
wire     [31:0] n31556;
wire     [31:0] n31557;
wire     [31:0] n31558;
wire     [31:0] n31559;
wire     [31:0] n31560;
wire     [31:0] n31561;
wire     [31:0] n31562;
wire     [31:0] n31563;
wire     [31:0] n31564;
wire     [31:0] n31565;
wire     [31:0] n31566;
wire     [31:0] n31567;
wire     [31:0] n31568;
wire     [31:0] n31569;
wire     [31:0] n31570;
wire     [31:0] n31571;
wire     [31:0] n31572;
wire     [31:0] n31573;
wire     [31:0] n31574;
wire     [31:0] n31575;
wire     [31:0] n31576;
wire     [31:0] n31577;
wire     [31:0] n31578;
wire     [31:0] n31579;
wire     [31:0] n31580;
wire     [31:0] n31581;
wire     [31:0] n31582;
wire     [31:0] n31583;
wire     [31:0] n31584;
wire     [31:0] n31585;
wire     [31:0] n31586;
wire     [31:0] n31587;
wire     [31:0] n31588;
wire     [31:0] n31589;
wire     [31:0] n31590;
wire     [31:0] n31591;
wire     [31:0] n31592;
wire     [31:0] n31593;
wire     [31:0] n31594;
wire     [31:0] n31595;
wire     [31:0] n31596;
wire     [31:0] n31597;
wire     [31:0] n31598;
wire     [31:0] n31599;
wire     [31:0] n31600;
wire     [31:0] n31601;
wire     [31:0] n31602;
wire     [31:0] n31603;
wire     [31:0] n31604;
wire     [31:0] n31605;
wire     [31:0] n31606;
wire     [31:0] n31607;
wire     [31:0] n31608;
wire     [31:0] n31609;
wire     [31:0] n31610;
wire     [31:0] n31611;
wire     [31:0] n31612;
wire     [31:0] n31613;
wire     [31:0] n31614;
wire     [31:0] n31615;
wire     [31:0] n31616;
wire     [31:0] n31617;
wire     [31:0] n31618;
wire     [31:0] n31619;
wire     [31:0] n31620;
wire     [31:0] n31621;
wire     [31:0] n31622;
wire     [31:0] n31623;
wire     [31:0] n31624;
wire     [31:0] n31625;
wire     [31:0] n31626;
wire     [31:0] n31627;
wire     [31:0] n31628;
wire     [31:0] n31629;
wire     [31:0] n31630;
wire     [31:0] n31631;
wire     [31:0] n31632;
wire     [31:0] n31633;
wire     [31:0] n31634;
wire     [31:0] n31635;
wire     [31:0] n31636;
wire     [31:0] n31637;
wire     [31:0] n31638;
wire     [31:0] n31639;
wire     [31:0] n31640;
wire     [31:0] n31641;
wire     [31:0] n31642;
wire     [31:0] n31643;
wire     [31:0] n31644;
wire     [31:0] n31645;
wire     [31:0] n31646;
wire     [31:0] n31647;
wire     [31:0] n31648;
wire     [31:0] n31649;
wire     [31:0] n31650;
wire     [31:0] n31651;
wire     [31:0] n31652;
wire     [31:0] n31653;
wire     [31:0] n31654;
wire     [31:0] n31655;
wire     [31:0] n31656;
wire     [31:0] n31657;
wire     [31:0] n31658;
wire     [31:0] n31659;
wire     [31:0] n31660;
wire     [31:0] n31661;
wire     [31:0] n31662;
wire     [31:0] n31663;
wire     [31:0] n31664;
wire     [31:0] n31665;
wire            n31666;
wire            n31667;
wire            n31668;
wire            n31669;
wire            n31670;
wire            n31671;
wire            n31672;
wire            n31673;
wire            n31674;
wire            n31675;
wire            n31676;
wire            n31677;
wire            n31678;
wire            n31679;
wire            n31680;
wire            n31681;
wire            n31682;
wire            n31683;
wire            n31684;
wire            n31685;
wire            n31686;
wire            n31687;
wire            n31688;
wire            n31689;
wire            n31690;
wire            n31691;
wire            n31692;
wire            n31693;
wire            n31694;
wire            n31695;
wire            n31696;
wire            n31697;
wire            n31698;
wire            n31699;
wire            n31700;
wire            n31701;
wire            n31702;
wire            n31703;
wire            n31704;
wire            n31705;
wire            n31706;
wire            n31707;
wire            n31708;
wire            n31709;
wire            n31710;
wire            n31711;
wire            n31712;
wire            n31713;
wire            n31714;
wire            n31715;
wire            n31716;
wire            n31717;
wire            n31718;
wire            n31719;
wire            n31720;
wire            n31721;
wire            n31722;
wire            n31723;
wire            n31724;
wire            n31725;
wire            n31726;
wire            n31727;
wire            n31728;
wire            n31729;
wire            n31730;
wire            n31731;
wire            n31732;
wire            n31733;
wire            n31734;
wire            n31735;
wire            n31736;
wire            n31737;
wire            n31738;
wire            n31739;
wire            n31740;
wire            n31741;
wire            n31742;
wire            n31743;
wire            n31744;
wire            n31745;
wire            n31746;
wire            n31747;
wire            n31748;
wire            n31749;
wire            n31750;
wire            n31751;
wire            n31752;
wire            n31753;
wire            n31754;
wire            n31755;
wire            n31756;
wire            n31757;
wire            n31758;
wire            n31759;
wire            n31760;
wire            n31761;
wire            n31762;
wire            n31763;
wire            n31764;
wire            n31765;
wire            n31766;
wire            n31767;
wire            n31768;
wire            n31769;
wire            n31770;
wire            n31771;
wire            n31772;
wire            n31773;
wire            n31774;
wire            n31775;
wire            n31776;
wire            n31777;
wire            n31778;
wire            n31779;
wire            n31780;
wire            n31781;
wire            n31782;
wire            n31783;
wire            n31784;
wire            n31785;
wire            n31786;
wire            n31787;
wire            n31788;
wire            n31789;
wire            n31790;
wire            n31791;
wire            n31792;
wire            n31793;
wire            n31794;
wire            n31795;
wire            n31796;
wire            n31797;
wire            n31798;
wire            n31799;
wire            n31800;
wire            n31801;
wire            n31802;
wire            n31803;
wire            n31804;
wire            n31805;
wire            n31806;
wire            n31807;
wire            n31808;
wire            n31809;
wire            n31810;
wire            n31811;
wire            n31812;
wire            n31813;
wire            n31814;
wire            n31815;
wire            n31816;
wire            n31817;
wire            n31818;
wire            n31819;
wire            n31820;
wire            n31821;
wire            n31822;
wire            n31823;
wire            n31824;
wire            n31825;
wire            n31826;
wire            n31827;
wire            n31828;
wire            n31829;
wire            n31830;
wire            n31831;
wire            n31832;
wire            n31833;
wire            n31834;
wire            n31835;
wire            n31836;
wire            n31837;
wire            n31838;
wire            n31839;
wire            n31840;
wire            n31841;
wire            n31842;
wire            n31843;
wire            n31844;
wire            n31845;
wire            n31846;
wire            n31847;
wire            n31848;
wire            n31849;
wire            n31850;
wire            n31851;
wire            n31852;
wire            n31853;
wire            n31854;
wire            n31855;
wire            n31856;
wire            n31857;
wire            n31858;
wire            n31859;
wire            n31860;
wire            n31861;
wire            n31862;
wire            n31863;
wire            n31864;
wire            n31865;
wire            n31866;
wire            n31867;
wire            n31868;
wire            n31869;
wire            n31870;
wire            n31871;
wire            n31872;
wire            n31873;
wire            n31874;
wire            n31875;
wire            n31876;
wire            n31877;
wire            n31878;
wire            n31879;
wire            n31880;
wire            n31881;
wire            n31882;
wire            n31883;
wire            n31884;
wire            n31885;
wire            n31886;
wire            n31887;
wire            n31888;
wire            n31889;
wire            n31890;
wire            n31891;
wire            n31892;
wire            n31893;
wire            n31894;
wire            n31895;
wire            n31896;
wire            n31897;
wire            n31898;
wire            n31899;
wire            n31900;
wire            n31901;
wire            n31902;
wire            n31903;
wire            n31904;
wire            n31905;
wire            n31906;
wire            n31907;
wire            n31908;
wire            n31909;
wire            n31910;
wire            n31911;
wire            n31912;
wire            n31913;
wire            n31914;
wire            n31915;
wire            n31916;
wire            n31917;
wire            n31918;
wire            n31919;
wire            n31920;
wire            n31921;
wire            n31922;
wire            n31923;
wire            n31924;
wire            n31925;
wire            n31926;
wire            n31927;
wire            n31928;
wire            n31929;
wire            n31930;
wire            n31931;
wire            n31932;
wire            n31933;
wire            n31934;
wire            n31935;
wire            n31936;
wire            n31937;
wire            n31938;
wire            n31939;
wire            n31940;
wire            n31941;
wire            n31942;
wire            n31943;
wire            n31944;
wire            n31945;
wire            n31946;
wire            n31947;
wire            n31948;
wire            n31949;
wire            n31950;
wire            n31951;
wire            n31952;
wire            n31953;
wire            n31954;
wire            n31955;
wire            n31956;
wire            n31957;
wire            n31958;
wire            n31959;
wire            n31960;
wire            n31961;
wire            n31962;
wire            n31963;
wire            n31964;
wire            n31965;
wire            n31966;
wire            n31967;
wire            n31968;
wire            n31969;
wire            n31970;
wire            n31971;
wire            n31972;
wire            n31973;
wire            n31974;
wire            n31975;
wire            n31976;
wire            n31977;
wire            n31978;
wire            n31979;
wire            n31980;
wire            n31981;
wire            n31982;
wire            n31983;
wire            n31984;
wire            n31985;
wire            n31986;
wire            n31987;
wire            n31988;
wire            n31989;
wire            n31990;
wire            n31991;
wire            n31992;
wire            n31993;
wire            n31994;
wire            n31995;
wire            n31996;
wire            n31997;
wire            n31998;
wire            n31999;
wire            n32000;
wire            n32001;
wire            n32002;
wire            n32003;
wire            n32004;
wire            n32005;
wire            n32006;
wire            n32007;
wire            n32008;
wire            n32009;
wire            n32010;
wire            n32011;
wire            n32012;
wire            n32013;
wire            n32014;
wire            n32015;
wire            n32016;
wire            n32017;
wire            n32018;
wire            n32019;
wire            n32020;
wire            n32021;
wire            n32022;
wire            n32023;
wire            n32024;
wire            n32025;
wire            n32026;
wire            n32027;
wire            n32028;
wire            n32029;
wire            n32030;
wire            n32031;
wire            n32032;
wire            n32033;
wire            n32034;
wire            n32035;
wire            n32036;
wire            n32037;
wire            n32038;
wire            n32039;
wire            n32040;
wire            n32041;
wire            n32042;
wire            n32043;
wire            n32044;
wire            n32045;
wire            n32046;
wire            n32047;
wire            n32048;
wire            n32049;
wire            n32050;
wire            n32051;
wire            n32052;
wire            n32053;
wire            n32054;
wire            n32055;
wire            n32056;
wire            n32057;
wire            n32058;
wire            n32059;
wire            n32060;
wire            n32061;
wire            n32062;
wire            n32063;
wire            n32064;
wire            n32065;
wire            n32066;
wire            n32067;
wire            n32068;
wire            n32069;
wire            n32070;
wire            n32071;
wire            n32072;
wire            n32073;
wire            n32074;
wire            n32075;
wire            n32076;
wire            n32077;
wire            n32078;
wire            n32079;
wire            n32080;
wire            n32081;
wire            n32082;
wire            n32083;
wire            n32084;
wire            n32085;
wire            n32086;
wire            n32087;
wire            n32088;
wire            n32089;
wire            n32090;
wire            n32091;
wire            n32092;
wire            n32093;
wire            n32094;
wire            n32095;
wire            n32096;
wire            n32097;
wire            n32098;
wire            n32099;
wire            n32100;
wire            n32101;
wire            n32102;
wire            n32103;
wire            n32104;
wire            n32105;
wire            n32106;
wire            n32107;
wire            n32108;
wire            n32109;
wire            n32110;
wire            n32111;
wire            n32112;
wire            n32113;
wire            n32114;
wire            n32115;
wire            n32116;
wire            n32117;
wire            n32118;
wire            n32119;
wire            n32120;
wire            n32121;
wire            n32122;
wire            n32123;
wire            n32124;
wire            n32125;
wire            n32126;
wire            n32127;
wire            n32128;
wire            n32129;
wire            n32130;
wire            n32131;
wire            n32132;
wire            n32133;
wire            n32134;
wire            n32135;
wire            n32136;
wire            n32137;
wire            n32138;
wire            n32139;
wire            n32140;
wire            n32141;
wire            n32142;
wire            n32143;
wire            n32144;
wire            n32145;
wire            n32146;
wire            n32147;
wire            n32148;
wire            n32149;
wire            n32150;
wire            n32151;
wire            n32152;
wire            n32153;
wire            n32154;
wire            n32155;
wire            n32156;
wire            n32157;
wire            n32158;
wire            n32159;
wire            n32160;
wire            n32161;
wire            n32162;
wire            n32163;
wire            n32164;
wire            n32165;
wire            n32166;
wire            n32167;
wire            n32168;
wire            n32169;
wire            n32170;
wire            n32171;
wire            n32172;
wire            n32173;
wire            n32174;
wire            n32175;
wire            n32176;
wire            n32177;
wire     [31:0] n32178;
wire     [31:0] n32179;
wire     [31:0] n32180;
wire     [31:0] n32181;
wire     [31:0] n32182;
wire     [31:0] n32183;
wire     [31:0] n32184;
wire     [31:0] n32185;
wire     [31:0] n32186;
wire     [31:0] n32187;
wire     [31:0] n32188;
wire     [31:0] n32189;
wire     [31:0] n32190;
wire     [31:0] n32191;
wire     [31:0] n32192;
wire     [31:0] n32193;
wire     [31:0] n32194;
wire     [31:0] n32195;
wire     [31:0] n32196;
wire     [31:0] n32197;
wire     [31:0] n32198;
wire     [31:0] n32199;
wire     [31:0] n32200;
wire     [31:0] n32201;
wire     [31:0] n32202;
wire     [31:0] n32203;
wire     [31:0] n32204;
wire     [31:0] n32205;
wire     [31:0] n32206;
wire     [31:0] n32207;
wire     [31:0] n32208;
wire     [31:0] n32209;
wire     [31:0] n32210;
wire     [31:0] n32211;
wire     [31:0] n32212;
wire     [31:0] n32213;
wire     [31:0] n32214;
wire     [31:0] n32215;
wire     [31:0] n32216;
wire     [31:0] n32217;
wire     [31:0] n32218;
wire     [31:0] n32219;
wire     [31:0] n32220;
wire     [31:0] n32221;
wire     [31:0] n32222;
wire     [31:0] n32223;
wire     [31:0] n32224;
wire     [31:0] n32225;
wire     [31:0] n32226;
wire     [31:0] n32227;
wire     [31:0] n32228;
wire     [31:0] n32229;
wire     [31:0] n32230;
wire     [31:0] n32231;
wire     [31:0] n32232;
wire     [31:0] n32233;
wire     [31:0] n32234;
wire     [31:0] n32235;
wire     [31:0] n32236;
wire     [31:0] n32237;
wire     [31:0] n32238;
wire     [31:0] n32239;
wire     [31:0] n32240;
wire     [31:0] n32241;
wire     [31:0] n32242;
wire     [31:0] n32243;
wire     [31:0] n32244;
wire     [31:0] n32245;
wire     [31:0] n32246;
wire     [31:0] n32247;
wire     [31:0] n32248;
wire     [31:0] n32249;
wire     [31:0] n32250;
wire     [31:0] n32251;
wire     [31:0] n32252;
wire     [31:0] n32253;
wire     [31:0] n32254;
wire     [31:0] n32255;
wire     [31:0] n32256;
wire     [31:0] n32257;
wire     [31:0] n32258;
wire     [31:0] n32259;
wire     [31:0] n32260;
wire     [31:0] n32261;
wire     [31:0] n32262;
wire     [31:0] n32263;
wire     [31:0] n32264;
wire     [31:0] n32265;
wire     [31:0] n32266;
wire     [31:0] n32267;
wire     [31:0] n32268;
wire     [31:0] n32269;
wire     [31:0] n32270;
wire     [31:0] n32271;
wire     [31:0] n32272;
wire     [31:0] n32273;
wire     [31:0] n32274;
wire     [31:0] n32275;
wire     [31:0] n32276;
wire     [31:0] n32277;
wire     [31:0] n32278;
wire     [31:0] n32279;
wire     [31:0] n32280;
wire     [31:0] n32281;
wire     [31:0] n32282;
wire     [31:0] n32283;
wire     [31:0] n32284;
wire     [31:0] n32285;
wire     [31:0] n32286;
wire     [31:0] n32287;
wire     [31:0] n32288;
wire     [31:0] n32289;
wire     [31:0] n32290;
wire     [31:0] n32291;
wire     [31:0] n32292;
wire     [31:0] n32293;
wire     [31:0] n32294;
wire     [31:0] n32295;
wire     [31:0] n32296;
wire     [31:0] n32297;
wire     [31:0] n32298;
wire     [31:0] n32299;
wire     [31:0] n32300;
wire     [31:0] n32301;
wire     [31:0] n32302;
wire     [31:0] n32303;
wire     [31:0] n32304;
wire     [31:0] n32305;
wire     [31:0] n32306;
wire     [31:0] n32307;
wire     [31:0] n32308;
wire     [31:0] n32309;
wire     [31:0] n32310;
wire     [31:0] n32311;
wire     [31:0] n32312;
wire     [31:0] n32313;
wire     [31:0] n32314;
wire     [31:0] n32315;
wire     [31:0] n32316;
wire     [31:0] n32317;
wire     [31:0] n32318;
wire     [31:0] n32319;
wire     [31:0] n32320;
wire     [31:0] n32321;
wire     [31:0] n32322;
wire     [31:0] n32323;
wire     [31:0] n32324;
wire     [31:0] n32325;
wire     [31:0] n32326;
wire     [31:0] n32327;
wire     [31:0] n32328;
wire     [31:0] n32329;
wire     [31:0] n32330;
wire     [31:0] n32331;
wire     [31:0] n32332;
wire     [31:0] n32333;
wire     [31:0] n32334;
wire     [31:0] n32335;
wire     [31:0] n32336;
wire     [31:0] n32337;
wire     [31:0] n32338;
wire     [31:0] n32339;
wire     [31:0] n32340;
wire     [31:0] n32341;
wire     [31:0] n32342;
wire     [31:0] n32343;
wire     [31:0] n32344;
wire     [31:0] n32345;
wire     [31:0] n32346;
wire     [31:0] n32347;
wire     [31:0] n32348;
wire     [31:0] n32349;
wire     [31:0] n32350;
wire     [31:0] n32351;
wire     [31:0] n32352;
wire     [31:0] n32353;
wire     [31:0] n32354;
wire     [31:0] n32355;
wire     [31:0] n32356;
wire     [31:0] n32357;
wire     [31:0] n32358;
wire     [31:0] n32359;
wire     [31:0] n32360;
wire     [31:0] n32361;
wire     [31:0] n32362;
wire     [31:0] n32363;
wire     [31:0] n32364;
wire     [31:0] n32365;
wire     [31:0] n32366;
wire     [31:0] n32367;
wire     [31:0] n32368;
wire     [31:0] n32369;
wire     [31:0] n32370;
wire     [31:0] n32371;
wire     [31:0] n32372;
wire     [31:0] n32373;
wire     [31:0] n32374;
wire     [31:0] n32375;
wire     [31:0] n32376;
wire     [31:0] n32377;
wire     [31:0] n32378;
wire     [31:0] n32379;
wire     [31:0] n32380;
wire     [31:0] n32381;
wire     [31:0] n32382;
wire     [31:0] n32383;
wire     [31:0] n32384;
wire     [31:0] n32385;
wire     [31:0] n32386;
wire     [31:0] n32387;
wire     [31:0] n32388;
wire     [31:0] n32389;
wire     [31:0] n32390;
wire     [31:0] n32391;
wire     [31:0] n32392;
wire     [31:0] n32393;
wire     [31:0] n32394;
wire     [31:0] n32395;
wire     [31:0] n32396;
wire     [31:0] n32397;
wire     [31:0] n32398;
wire     [31:0] n32399;
wire     [31:0] n32400;
wire     [31:0] n32401;
wire     [31:0] n32402;
wire     [31:0] n32403;
wire     [31:0] n32404;
wire     [31:0] n32405;
wire     [31:0] n32406;
wire     [31:0] n32407;
wire     [31:0] n32408;
wire     [31:0] n32409;
wire     [31:0] n32410;
wire     [31:0] n32411;
wire     [31:0] n32412;
wire     [31:0] n32413;
wire     [31:0] n32414;
wire     [31:0] n32415;
wire     [31:0] n32416;
wire     [31:0] n32417;
wire     [31:0] n32418;
wire     [31:0] n32419;
wire     [31:0] n32420;
wire     [31:0] n32421;
wire     [31:0] n32422;
wire     [31:0] n32423;
wire     [31:0] n32424;
wire     [31:0] n32425;
wire     [31:0] n32426;
wire     [31:0] n32427;
wire     [31:0] n32428;
wire     [31:0] n32429;
wire     [31:0] n32430;
wire     [31:0] n32431;
wire     [31:0] n32432;
wire     [31:0] n32433;
wire     [31:0] n32434;
wire     [31:0] n32435;
wire     [31:0] n32436;
wire     [31:0] n32437;
wire     [31:0] n32438;
wire     [31:0] n32439;
wire     [31:0] n32440;
wire     [31:0] n32441;
wire     [31:0] n32442;
wire     [31:0] n32443;
wire     [31:0] n32444;
wire     [31:0] n32445;
wire     [31:0] n32446;
wire     [31:0] n32447;
wire     [31:0] n32448;
wire     [31:0] n32449;
wire     [31:0] n32450;
wire     [31:0] n32451;
wire     [31:0] n32452;
wire     [31:0] n32453;
wire     [31:0] n32454;
wire     [31:0] n32455;
wire     [31:0] n32456;
wire     [31:0] n32457;
wire     [31:0] n32458;
wire     [31:0] n32459;
wire     [31:0] n32460;
wire     [31:0] n32461;
wire     [31:0] n32462;
wire     [31:0] n32463;
wire     [31:0] n32464;
wire     [31:0] n32465;
wire     [31:0] n32466;
wire     [31:0] n32467;
wire     [31:0] n32468;
wire     [31:0] n32469;
wire     [31:0] n32470;
wire     [31:0] n32471;
wire     [31:0] n32472;
wire     [31:0] n32473;
wire     [31:0] n32474;
wire     [31:0] n32475;
wire     [31:0] n32476;
wire     [31:0] n32477;
wire     [31:0] n32478;
wire     [31:0] n32479;
wire     [31:0] n32480;
wire     [31:0] n32481;
wire     [31:0] n32482;
wire     [31:0] n32483;
wire     [31:0] n32484;
wire     [31:0] n32485;
wire     [31:0] n32486;
wire     [31:0] n32487;
wire     [31:0] n32488;
wire     [31:0] n32489;
wire     [31:0] n32490;
wire     [31:0] n32491;
wire     [31:0] n32492;
wire     [31:0] n32493;
wire     [31:0] n32494;
wire     [31:0] n32495;
wire     [31:0] n32496;
wire     [31:0] n32497;
wire     [31:0] n32498;
wire     [31:0] n32499;
wire     [31:0] n32500;
wire     [31:0] n32501;
wire     [31:0] n32502;
wire     [31:0] n32503;
wire     [31:0] n32504;
wire     [31:0] n32505;
wire     [31:0] n32506;
wire     [31:0] n32507;
wire     [31:0] n32508;
wire     [31:0] n32509;
wire     [31:0] n32510;
wire     [31:0] n32511;
wire     [31:0] n32512;
wire     [31:0] n32513;
wire     [31:0] n32514;
wire     [31:0] n32515;
wire     [31:0] n32516;
wire     [31:0] n32517;
wire     [31:0] n32518;
wire     [31:0] n32519;
wire     [31:0] n32520;
wire     [31:0] n32521;
wire     [31:0] n32522;
wire     [31:0] n32523;
wire     [31:0] n32524;
wire     [31:0] n32525;
wire     [31:0] n32526;
wire     [31:0] n32527;
wire     [31:0] n32528;
wire     [31:0] n32529;
wire     [31:0] n32530;
wire     [31:0] n32531;
wire     [31:0] n32532;
wire     [31:0] n32533;
wire     [31:0] n32534;
wire     [31:0] n32535;
wire     [31:0] n32536;
wire     [31:0] n32537;
wire     [31:0] n32538;
wire     [31:0] n32539;
wire     [31:0] n32540;
wire     [31:0] n32541;
wire     [31:0] n32542;
wire     [31:0] n32543;
wire     [31:0] n32544;
wire     [31:0] n32545;
wire     [31:0] n32546;
wire     [31:0] n32547;
wire     [31:0] n32548;
wire     [31:0] n32549;
wire     [31:0] n32550;
wire     [31:0] n32551;
wire     [31:0] n32552;
wire     [31:0] n32553;
wire     [31:0] n32554;
wire     [31:0] n32555;
wire     [31:0] n32556;
wire     [31:0] n32557;
wire     [31:0] n32558;
wire     [31:0] n32559;
wire     [31:0] n32560;
wire     [31:0] n32561;
wire     [31:0] n32562;
wire     [31:0] n32563;
wire     [31:0] n32564;
wire     [31:0] n32565;
wire     [31:0] n32566;
wire     [31:0] n32567;
wire     [31:0] n32568;
wire     [31:0] n32569;
wire     [31:0] n32570;
wire     [31:0] n32571;
wire     [31:0] n32572;
wire     [31:0] n32573;
wire     [31:0] n32574;
wire     [31:0] n32575;
wire     [31:0] n32576;
wire     [31:0] n32577;
wire     [31:0] n32578;
wire     [31:0] n32579;
wire     [31:0] n32580;
wire     [31:0] n32581;
wire     [31:0] n32582;
wire     [31:0] n32583;
wire     [31:0] n32584;
wire     [31:0] n32585;
wire     [31:0] n32586;
wire     [31:0] n32587;
wire     [31:0] n32588;
wire     [31:0] n32589;
wire     [31:0] n32590;
wire     [31:0] n32591;
wire     [31:0] n32592;
wire     [31:0] n32593;
wire     [31:0] n32594;
wire     [31:0] n32595;
wire     [31:0] n32596;
wire     [31:0] n32597;
wire     [31:0] n32598;
wire     [31:0] n32599;
wire     [31:0] n32600;
wire     [31:0] n32601;
wire     [31:0] n32602;
wire     [31:0] n32603;
wire     [31:0] n32604;
wire     [31:0] n32605;
wire     [31:0] n32606;
wire     [31:0] n32607;
wire     [31:0] n32608;
wire     [31:0] n32609;
wire     [31:0] n32610;
wire     [31:0] n32611;
wire     [31:0] n32612;
wire     [31:0] n32613;
wire     [31:0] n32614;
wire     [31:0] n32615;
wire     [31:0] n32616;
wire     [31:0] n32617;
wire     [31:0] n32618;
wire     [31:0] n32619;
wire     [31:0] n32620;
wire     [31:0] n32621;
wire     [31:0] n32622;
wire     [31:0] n32623;
wire     [31:0] n32624;
wire     [31:0] n32625;
wire     [31:0] n32626;
wire     [31:0] n32627;
wire     [31:0] n32628;
wire     [31:0] n32629;
wire     [31:0] n32630;
wire     [31:0] n32631;
wire     [31:0] n32632;
wire     [31:0] n32633;
wire     [31:0] n32634;
wire     [31:0] n32635;
wire     [31:0] n32636;
wire     [31:0] n32637;
wire     [31:0] n32638;
wire     [31:0] n32639;
wire     [31:0] n32640;
wire     [31:0] n32641;
wire     [31:0] n32642;
wire     [31:0] n32643;
wire     [31:0] n32644;
wire     [31:0] n32645;
wire     [31:0] n32646;
wire     [31:0] n32647;
wire     [31:0] n32648;
wire     [31:0] n32649;
wire     [31:0] n32650;
wire     [31:0] n32651;
wire     [31:0] n32652;
wire     [31:0] n32653;
wire     [31:0] n32654;
wire     [31:0] n32655;
wire     [31:0] n32656;
wire     [31:0] n32657;
wire     [31:0] n32658;
wire     [31:0] n32659;
wire     [31:0] n32660;
wire     [31:0] n32661;
wire     [31:0] n32662;
wire     [31:0] n32663;
wire     [31:0] n32664;
wire     [31:0] n32665;
wire     [31:0] n32666;
wire     [31:0] n32667;
wire     [31:0] n32668;
wire     [31:0] n32669;
wire     [31:0] n32670;
wire     [31:0] n32671;
wire     [31:0] n32672;
wire     [31:0] n32673;
wire     [31:0] n32674;
wire     [31:0] n32675;
wire     [31:0] n32676;
wire     [31:0] n32677;
wire     [31:0] n32678;
wire     [31:0] n32679;
wire     [31:0] n32680;
wire     [31:0] n32681;
wire     [31:0] n32682;
wire     [31:0] n32683;
wire     [31:0] n32684;
wire     [31:0] n32685;
wire     [31:0] n32686;
wire     [31:0] n32687;
wire     [31:0] n32688;
wire     [31:0] n32689;
wire     [31:0] n32690;
wire     [31:0] n32691;
wire     [31:0] n32692;
wire     [31:0] n32693;
wire     [31:0] n32694;
wire     [31:0] n32695;
wire     [31:0] n32696;
wire     [31:0] n32697;
wire     [31:0] n32698;
wire     [31:0] n32699;
wire            n32700;
wire            n32701;
wire     [31:0] n32702;
wire     [31:0] n32703;
wire     [31:0] n32704;
wire     [31:0] n32705;
wire     [31:0] n32706;
wire     [31:0] n32707;
wire     [31:0] n32708;
wire     [31:0] n32709;
wire     [31:0] n32710;
wire     [31:0] n32711;
wire     [31:0] n32712;
wire     [31:0] n32713;
wire     [31:0] n32714;
wire     [31:0] n32715;
wire     [31:0] n32716;
wire     [31:0] n32717;
wire     [31:0] n32718;
wire     [31:0] n32719;
wire     [31:0] n32720;
wire     [31:0] n32721;
wire     [31:0] n32722;
wire     [31:0] n32723;
wire     [31:0] n32724;
wire     [31:0] n32725;
wire     [31:0] n32726;
wire     [31:0] n32727;
wire     [31:0] n32728;
wire     [31:0] n32729;
wire     [31:0] n32730;
wire     [31:0] n32731;
wire     [31:0] n32732;
wire     [31:0] n32733;
wire     [31:0] n32734;
wire            n32735;
wire            n32736;
wire            n32737;
wire            n32738;
wire            n32739;
wire            n32740;
wire            n32741;
wire            n32742;
wire            n32743;
wire            n32744;
wire            n32745;
wire            n32746;
wire            n32747;
wire            n32748;
wire            n32749;
wire            n32750;
wire            n32751;
wire            n32752;
wire            n32753;
wire            n32754;
wire            n32755;
wire            n32756;
wire            n32757;
wire            n32758;
wire            n32759;
wire            n32760;
wire            n32761;
wire            n32762;
wire            n32763;
wire            n32764;
wire            n32765;
wire            n32766;
wire            n32767;
wire            n32768;
wire            n32769;
wire            n32770;
wire            n32771;
wire            n32772;
wire            n32773;
wire            n32774;
wire            n32775;
wire            n32776;
wire            n32777;
wire            n32778;
wire            n32779;
wire            n32780;
wire            n32781;
wire            n32782;
wire            n32783;
wire            n32784;
wire            n32785;
wire            n32786;
wire            n32787;
wire            n32788;
wire            n32789;
wire            n32790;
wire            n32791;
wire            n32792;
wire            n32793;
wire            n32794;
wire            n32795;
wire            n32796;
wire            n32797;
wire            n32798;
wire            n32799;
wire            n32800;
wire            n32801;
wire            n32802;
wire            n32803;
wire            n32804;
wire            n32805;
wire            n32806;
wire            n32807;
wire            n32808;
wire            n32809;
wire            n32810;
wire            n32811;
wire            n32812;
wire            n32813;
wire            n32814;
wire            n32815;
wire            n32816;
wire            n32817;
wire            n32818;
wire            n32819;
wire            n32820;
wire            n32821;
wire            n32822;
wire            n32823;
wire            n32824;
wire            n32825;
wire            n32826;
wire            n32827;
wire            n32828;
wire            n32829;
wire            n32830;
wire            n32831;
wire            n32832;
wire            n32833;
wire            n32834;
wire            n32835;
wire            n32836;
wire            n32837;
wire            n32838;
wire            n32839;
wire            n32840;
wire            n32841;
wire            n32842;
wire            n32843;
wire            n32844;
wire            n32845;
wire            n32846;
wire            n32847;
wire            n32848;
wire            n32849;
wire            n32850;
wire            n32851;
wire            n32852;
wire            n32853;
wire            n32854;
wire            n32855;
wire            n32856;
wire            n32857;
wire            n32858;
wire            n32859;
wire            n32860;
wire            n32861;
wire            n32862;
wire            n32863;
wire            n32864;
wire            n32865;
wire            n32866;
wire            n32867;
wire            n32868;
wire            n32869;
wire            n32870;
wire            n32871;
wire            n32872;
wire            n32873;
wire            n32874;
wire            n32875;
wire            n32876;
wire            n32877;
wire            n32878;
wire            n32879;
wire            n32880;
wire            n32881;
wire            n32882;
wire            n32883;
wire            n32884;
wire            n32885;
wire            n32886;
wire            n32887;
wire            n32888;
wire            n32889;
wire            n32890;
wire            n32891;
wire            n32892;
wire            n32893;
wire            n32894;
wire            n32895;
wire            n32896;
wire            n32897;
wire            n32898;
wire            n32899;
wire            n32900;
wire            n32901;
wire            n32902;
wire            n32903;
wire            n32904;
wire            n32905;
wire            n32906;
wire            n32907;
wire            n32908;
wire            n32909;
wire            n32910;
wire            n32911;
wire            n32912;
wire            n32913;
wire            n32914;
wire            n32915;
wire            n32916;
wire            n32917;
wire            n32918;
wire            n32919;
wire            n32920;
wire            n32921;
wire            n32922;
wire            n32923;
wire            n32924;
wire            n32925;
wire            n32926;
wire            n32927;
wire            n32928;
wire            n32929;
wire            n32930;
wire            n32931;
wire            n32932;
wire            n32933;
wire            n32934;
wire            n32935;
wire            n32936;
wire            n32937;
wire            n32938;
wire            n32939;
wire            n32940;
wire            n32941;
wire            n32942;
wire            n32943;
wire            n32944;
wire            n32945;
wire            n32946;
wire            n32947;
wire            n32948;
wire            n32949;
wire            n32950;
wire            n32951;
wire            n32952;
wire            n32953;
wire            n32954;
wire            n32955;
wire            n32956;
wire            n32957;
wire            n32958;
wire            n32959;
wire            n32960;
wire            n32961;
wire            n32962;
wire            n32963;
wire            n32964;
wire            n32965;
wire            n32966;
wire            n32967;
wire            n32968;
wire            n32969;
wire            n32970;
wire            n32971;
wire            n32972;
wire            n32973;
wire            n32974;
wire            n32975;
wire            n32976;
wire            n32977;
wire            n32978;
wire            n32979;
wire            n32980;
wire            n32981;
wire            n32982;
wire            n32983;
wire            n32984;
wire            n32985;
wire            n32986;
wire            n32987;
wire            n32988;
wire            n32989;
wire            n32990;
wire            n32991;
wire            n32992;
wire            n32993;
wire            n32994;
wire            n32995;
wire            n32996;
wire            n32997;
wire            n32998;
wire            n32999;
wire            n33000;
wire            n33001;
wire            n33002;
wire            n33003;
wire            n33004;
wire            n33005;
wire            n33006;
wire            n33007;
wire            n33008;
wire            n33009;
wire            n33010;
wire            n33011;
wire            n33012;
wire            n33013;
wire            n33014;
wire            n33015;
wire            n33016;
wire            n33017;
wire            n33018;
wire            n33019;
wire            n33020;
wire            n33021;
wire            n33022;
wire            n33023;
wire            n33024;
wire            n33025;
wire            n33026;
wire            n33027;
wire            n33028;
wire            n33029;
wire            n33030;
wire            n33031;
wire            n33032;
wire            n33033;
wire            n33034;
wire            n33035;
wire            n33036;
wire            n33037;
wire            n33038;
wire            n33039;
wire            n33040;
wire            n33041;
wire            n33042;
wire            n33043;
wire            n33044;
wire            n33045;
wire            n33046;
wire            n33047;
wire            n33048;
wire            n33049;
wire            n33050;
wire            n33051;
wire            n33052;
wire            n33053;
wire            n33054;
wire            n33055;
wire            n33056;
wire            n33057;
wire            n33058;
wire            n33059;
wire            n33060;
wire            n33061;
wire            n33062;
wire            n33063;
wire            n33064;
wire            n33065;
wire            n33066;
wire            n33067;
wire            n33068;
wire            n33069;
wire            n33070;
wire            n33071;
wire            n33072;
wire            n33073;
wire            n33074;
wire            n33075;
wire            n33076;
wire            n33077;
wire            n33078;
wire            n33079;
wire            n33080;
wire            n33081;
wire            n33082;
wire            n33083;
wire            n33084;
wire            n33085;
wire            n33086;
wire            n33087;
wire            n33088;
wire            n33089;
wire            n33090;
wire            n33091;
wire            n33092;
wire            n33093;
wire            n33094;
wire            n33095;
wire            n33096;
wire            n33097;
wire            n33098;
wire            n33099;
wire            n33100;
wire            n33101;
wire            n33102;
wire            n33103;
wire            n33104;
wire            n33105;
wire            n33106;
wire            n33107;
wire            n33108;
wire            n33109;
wire            n33110;
wire            n33111;
wire            n33112;
wire            n33113;
wire            n33114;
wire            n33115;
wire            n33116;
wire            n33117;
wire            n33118;
wire            n33119;
wire            n33120;
wire            n33121;
wire            n33122;
wire            n33123;
wire            n33124;
wire            n33125;
wire            n33126;
wire            n33127;
wire            n33128;
wire            n33129;
wire            n33130;
wire            n33131;
wire            n33132;
wire            n33133;
wire            n33134;
wire            n33135;
wire            n33136;
wire            n33137;
wire            n33138;
wire            n33139;
wire            n33140;
wire            n33141;
wire            n33142;
wire            n33143;
wire            n33144;
wire            n33145;
wire            n33146;
wire            n33147;
wire            n33148;
wire            n33149;
wire            n33150;
wire            n33151;
wire            n33152;
wire            n33153;
wire            n33154;
wire            n33155;
wire            n33156;
wire            n33157;
wire            n33158;
wire            n33159;
wire            n33160;
wire            n33161;
wire            n33162;
wire            n33163;
wire            n33164;
wire            n33165;
wire            n33166;
wire            n33167;
wire            n33168;
wire            n33169;
wire            n33170;
wire            n33171;
wire            n33172;
wire            n33173;
wire            n33174;
wire            n33175;
wire            n33176;
wire            n33177;
wire            n33178;
wire            n33179;
wire            n33180;
wire            n33181;
wire            n33182;
wire            n33183;
wire            n33184;
wire            n33185;
wire            n33186;
wire            n33187;
wire            n33188;
wire            n33189;
wire            n33190;
wire            n33191;
wire            n33192;
wire            n33193;
wire            n33194;
wire            n33195;
wire            n33196;
wire            n33197;
wire            n33198;
wire            n33199;
wire            n33200;
wire            n33201;
wire            n33202;
wire            n33203;
wire            n33204;
wire            n33205;
wire            n33206;
wire            n33207;
wire            n33208;
wire            n33209;
wire            n33210;
wire            n33211;
wire            n33212;
wire            n33213;
wire            n33214;
wire            n33215;
wire            n33216;
wire            n33217;
wire            n33218;
wire            n33219;
wire            n33220;
wire            n33221;
wire            n33222;
wire            n33223;
wire            n33224;
wire            n33225;
wire            n33226;
wire            n33227;
wire            n33228;
wire            n33229;
wire            n33230;
wire            n33231;
wire            n33232;
wire            n33233;
wire            n33234;
wire            n33235;
wire            n33236;
wire            n33237;
wire            n33238;
wire            n33239;
wire            n33240;
wire            n33241;
wire            n33242;
wire            n33243;
wire            n33244;
wire            n33245;
wire            n33246;
wire            n33247;
wire            n33248;
wire            n33249;
wire            n33250;
wire            n33251;
wire            n33252;
wire            n33253;
wire            n33254;
wire            n33255;
wire            n33256;
wire            n33257;
wire            n33258;
wire            n33259;
wire            n33260;
wire            n33261;
wire            n33262;
wire     [31:0] n33263;
wire     [31:0] n33264;
wire     [31:0] n33265;
wire     [31:0] n33266;
wire     [31:0] n33267;
wire     [31:0] n33268;
wire     [31:0] n33269;
wire     [31:0] n33270;
wire     [31:0] n33271;
wire     [31:0] n33272;
wire     [31:0] n33273;
wire     [31:0] n33274;
wire     [31:0] n33275;
wire     [31:0] n33276;
wire     [31:0] n33277;
wire     [31:0] n33278;
wire     [31:0] n33279;
wire     [31:0] n33280;
wire     [31:0] n33281;
wire     [31:0] n33282;
wire     [31:0] n33283;
wire     [31:0] n33284;
wire     [31:0] n33285;
wire     [31:0] n33286;
wire     [31:0] n33287;
wire     [31:0] n33288;
wire     [31:0] n33289;
wire     [31:0] n33290;
wire     [31:0] n33291;
wire     [31:0] n33292;
wire     [31:0] n33293;
wire     [31:0] n33294;
wire     [31:0] n33295;
wire     [31:0] n33296;
wire     [31:0] n33297;
wire     [31:0] n33298;
wire     [31:0] n33299;
wire     [31:0] n33300;
wire     [31:0] n33301;
wire     [31:0] n33302;
wire     [31:0] n33303;
wire     [31:0] n33304;
wire     [31:0] n33305;
wire     [31:0] n33306;
wire     [31:0] n33307;
wire     [31:0] n33308;
wire     [31:0] n33309;
wire     [31:0] n33310;
wire     [31:0] n33311;
wire     [31:0] n33312;
wire     [31:0] n33313;
wire     [31:0] n33314;
wire     [31:0] n33315;
wire     [31:0] n33316;
wire     [31:0] n33317;
wire     [31:0] n33318;
wire     [31:0] n33319;
wire     [31:0] n33320;
wire     [31:0] n33321;
wire     [31:0] n33322;
wire     [31:0] n33323;
wire     [31:0] n33324;
wire     [31:0] n33325;
wire     [31:0] n33326;
wire     [31:0] n33327;
wire     [31:0] n33328;
wire     [31:0] n33329;
wire     [31:0] n33330;
wire     [31:0] n33331;
wire     [31:0] n33332;
wire     [31:0] n33333;
wire     [31:0] n33334;
wire     [31:0] n33335;
wire     [31:0] n33336;
wire     [31:0] n33337;
wire     [31:0] n33338;
wire     [31:0] n33339;
wire     [31:0] n33340;
wire     [31:0] n33341;
wire     [31:0] n33342;
wire     [31:0] n33343;
wire     [31:0] n33344;
wire     [31:0] n33345;
wire     [31:0] n33346;
wire     [31:0] n33347;
wire     [31:0] n33348;
wire     [31:0] n33349;
wire     [31:0] n33350;
wire     [31:0] n33351;
wire     [31:0] n33352;
wire     [31:0] n33353;
wire     [31:0] n33354;
wire     [31:0] n33355;
wire     [31:0] n33356;
wire     [31:0] n33357;
wire     [31:0] n33358;
wire     [31:0] n33359;
wire     [31:0] n33360;
wire     [31:0] n33361;
wire     [31:0] n33362;
wire     [31:0] n33363;
wire     [31:0] n33364;
wire     [31:0] n33365;
wire     [31:0] n33366;
wire     [31:0] n33367;
wire     [31:0] n33368;
wire     [31:0] n33369;
wire     [31:0] n33370;
wire     [31:0] n33371;
wire     [31:0] n33372;
wire     [31:0] n33373;
wire     [31:0] n33374;
wire     [31:0] n33375;
wire     [31:0] n33376;
wire     [31:0] n33377;
wire     [31:0] n33378;
wire     [31:0] n33379;
wire     [31:0] n33380;
wire     [31:0] n33381;
wire     [31:0] n33382;
wire     [31:0] n33383;
wire     [31:0] n33384;
wire     [31:0] n33385;
wire     [31:0] n33386;
wire     [31:0] n33387;
wire     [31:0] n33388;
wire     [31:0] n33389;
wire     [31:0] n33390;
wire     [31:0] n33391;
wire     [31:0] n33392;
wire     [31:0] n33393;
wire     [31:0] n33394;
wire     [31:0] n33395;
wire     [31:0] n33396;
wire     [31:0] n33397;
wire     [31:0] n33398;
wire     [31:0] n33399;
wire     [31:0] n33400;
wire     [31:0] n33401;
wire     [31:0] n33402;
wire     [31:0] n33403;
wire     [31:0] n33404;
wire     [31:0] n33405;
wire     [31:0] n33406;
wire     [31:0] n33407;
wire     [31:0] n33408;
wire     [31:0] n33409;
wire     [31:0] n33410;
wire     [31:0] n33411;
wire     [31:0] n33412;
wire     [31:0] n33413;
wire     [31:0] n33414;
wire     [31:0] n33415;
wire     [31:0] n33416;
wire     [31:0] n33417;
wire     [31:0] n33418;
wire     [31:0] n33419;
wire     [31:0] n33420;
wire     [31:0] n33421;
wire     [31:0] n33422;
wire     [31:0] n33423;
wire     [31:0] n33424;
wire     [31:0] n33425;
wire     [31:0] n33426;
wire     [31:0] n33427;
wire     [31:0] n33428;
wire     [31:0] n33429;
wire     [31:0] n33430;
wire     [31:0] n33431;
wire     [31:0] n33432;
wire     [31:0] n33433;
wire     [31:0] n33434;
wire     [31:0] n33435;
wire     [31:0] n33436;
wire     [31:0] n33437;
wire     [31:0] n33438;
wire     [31:0] n33439;
wire     [31:0] n33440;
wire     [31:0] n33441;
wire     [31:0] n33442;
wire     [31:0] n33443;
wire     [31:0] n33444;
wire     [31:0] n33445;
wire     [31:0] n33446;
wire     [31:0] n33447;
wire     [31:0] n33448;
wire     [31:0] n33449;
wire     [31:0] n33450;
wire     [31:0] n33451;
wire     [31:0] n33452;
wire     [31:0] n33453;
wire     [31:0] n33454;
wire     [31:0] n33455;
wire     [31:0] n33456;
wire     [31:0] n33457;
wire     [31:0] n33458;
wire     [31:0] n33459;
wire     [31:0] n33460;
wire     [31:0] n33461;
wire     [31:0] n33462;
wire     [31:0] n33463;
wire     [31:0] n33464;
wire     [31:0] n33465;
wire     [31:0] n33466;
wire     [31:0] n33467;
wire     [31:0] n33468;
wire     [31:0] n33469;
wire     [31:0] n33470;
wire     [31:0] n33471;
wire     [31:0] n33472;
wire     [31:0] n33473;
wire     [31:0] n33474;
wire     [31:0] n33475;
wire     [31:0] n33476;
wire     [31:0] n33477;
wire     [31:0] n33478;
wire     [31:0] n33479;
wire     [31:0] n33480;
wire     [31:0] n33481;
wire     [31:0] n33482;
wire     [31:0] n33483;
wire     [31:0] n33484;
wire     [31:0] n33485;
wire     [31:0] n33486;
wire     [31:0] n33487;
wire     [31:0] n33488;
wire     [31:0] n33489;
wire     [31:0] n33490;
wire     [31:0] n33491;
wire     [31:0] n33492;
wire     [31:0] n33493;
wire     [31:0] n33494;
wire     [31:0] n33495;
wire     [31:0] n33496;
wire     [31:0] n33497;
wire     [31:0] n33498;
wire     [31:0] n33499;
wire     [31:0] n33500;
wire     [31:0] n33501;
wire     [31:0] n33502;
wire     [31:0] n33503;
wire     [31:0] n33504;
wire     [31:0] n33505;
wire     [31:0] n33506;
wire     [31:0] n33507;
wire     [31:0] n33508;
wire     [31:0] n33509;
wire     [31:0] n33510;
wire     [31:0] n33511;
wire     [31:0] n33512;
wire     [31:0] n33513;
wire     [31:0] n33514;
wire     [31:0] n33515;
wire     [31:0] n33516;
wire     [31:0] n33517;
wire     [31:0] n33518;
wire     [31:0] n33519;
wire     [31:0] n33520;
wire     [31:0] n33521;
wire     [31:0] n33522;
wire     [31:0] n33523;
wire     [31:0] n33524;
wire     [31:0] n33525;
wire     [31:0] n33526;
wire     [31:0] n33527;
wire     [31:0] n33528;
wire     [31:0] n33529;
wire     [31:0] n33530;
wire     [31:0] n33531;
wire     [31:0] n33532;
wire     [31:0] n33533;
wire     [31:0] n33534;
wire     [31:0] n33535;
wire     [31:0] n33536;
wire     [31:0] n33537;
wire     [31:0] n33538;
wire     [31:0] n33539;
wire     [31:0] n33540;
wire     [31:0] n33541;
wire     [31:0] n33542;
wire     [31:0] n33543;
wire     [31:0] n33544;
wire     [31:0] n33545;
wire     [31:0] n33546;
wire     [31:0] n33547;
wire     [31:0] n33548;
wire     [31:0] n33549;
wire     [31:0] n33550;
wire     [31:0] n33551;
wire     [31:0] n33552;
wire     [31:0] n33553;
wire     [31:0] n33554;
wire     [31:0] n33555;
wire     [31:0] n33556;
wire     [31:0] n33557;
wire     [31:0] n33558;
wire     [31:0] n33559;
wire     [31:0] n33560;
wire     [31:0] n33561;
wire     [31:0] n33562;
wire     [31:0] n33563;
wire     [31:0] n33564;
wire     [31:0] n33565;
wire     [31:0] n33566;
wire     [31:0] n33567;
wire     [31:0] n33568;
wire     [31:0] n33569;
wire     [31:0] n33570;
wire     [31:0] n33571;
wire     [31:0] n33572;
wire     [31:0] n33573;
wire     [31:0] n33574;
wire     [31:0] n33575;
wire     [31:0] n33576;
wire     [31:0] n33577;
wire     [31:0] n33578;
wire     [31:0] n33579;
wire     [31:0] n33580;
wire     [31:0] n33581;
wire     [31:0] n33582;
wire     [31:0] n33583;
wire     [31:0] n33584;
wire     [31:0] n33585;
wire     [31:0] n33586;
wire     [31:0] n33587;
wire     [31:0] n33588;
wire     [31:0] n33589;
wire     [31:0] n33590;
wire     [31:0] n33591;
wire     [31:0] n33592;
wire     [31:0] n33593;
wire     [31:0] n33594;
wire     [31:0] n33595;
wire     [31:0] n33596;
wire     [31:0] n33597;
wire     [31:0] n33598;
wire     [31:0] n33599;
wire     [31:0] n33600;
wire     [31:0] n33601;
wire     [31:0] n33602;
wire     [31:0] n33603;
wire     [31:0] n33604;
wire     [31:0] n33605;
wire     [31:0] n33606;
wire     [31:0] n33607;
wire     [31:0] n33608;
wire     [31:0] n33609;
wire     [31:0] n33610;
wire     [31:0] n33611;
wire     [31:0] n33612;
wire     [31:0] n33613;
wire     [31:0] n33614;
wire     [31:0] n33615;
wire     [31:0] n33616;
wire     [31:0] n33617;
wire     [31:0] n33618;
wire     [31:0] n33619;
wire     [31:0] n33620;
wire     [31:0] n33621;
wire     [31:0] n33622;
wire     [31:0] n33623;
wire     [31:0] n33624;
wire     [31:0] n33625;
wire     [31:0] n33626;
wire     [31:0] n33627;
wire     [31:0] n33628;
wire     [31:0] n33629;
wire     [31:0] n33630;
wire     [31:0] n33631;
wire     [31:0] n33632;
wire     [31:0] n33633;
wire     [31:0] n33634;
wire     [31:0] n33635;
wire     [31:0] n33636;
wire     [31:0] n33637;
wire     [31:0] n33638;
wire     [31:0] n33639;
wire     [31:0] n33640;
wire     [31:0] n33641;
wire     [31:0] n33642;
wire     [31:0] n33643;
wire     [31:0] n33644;
wire     [31:0] n33645;
wire     [31:0] n33646;
wire     [31:0] n33647;
wire     [31:0] n33648;
wire     [31:0] n33649;
wire     [31:0] n33650;
wire     [31:0] n33651;
wire     [31:0] n33652;
wire     [31:0] n33653;
wire     [31:0] n33654;
wire     [31:0] n33655;
wire     [31:0] n33656;
wire     [31:0] n33657;
wire     [31:0] n33658;
wire     [31:0] n33659;
wire     [31:0] n33660;
wire     [31:0] n33661;
wire     [31:0] n33662;
wire     [31:0] n33663;
wire     [31:0] n33664;
wire     [31:0] n33665;
wire     [31:0] n33666;
wire     [31:0] n33667;
wire     [31:0] n33668;
wire     [31:0] n33669;
wire     [31:0] n33670;
wire     [31:0] n33671;
wire     [31:0] n33672;
wire     [31:0] n33673;
wire     [31:0] n33674;
wire     [31:0] n33675;
wire     [31:0] n33676;
wire     [31:0] n33677;
wire     [31:0] n33678;
wire     [31:0] n33679;
wire     [31:0] n33680;
wire     [31:0] n33681;
wire     [31:0] n33682;
wire     [31:0] n33683;
wire     [31:0] n33684;
wire     [31:0] n33685;
wire     [31:0] n33686;
wire     [31:0] n33687;
wire     [31:0] n33688;
wire     [31:0] n33689;
wire     [31:0] n33690;
wire     [31:0] n33691;
wire     [31:0] n33692;
wire     [31:0] n33693;
wire     [31:0] n33694;
wire     [31:0] n33695;
wire     [31:0] n33696;
wire     [31:0] n33697;
wire     [31:0] n33698;
wire     [31:0] n33699;
wire     [31:0] n33700;
wire     [31:0] n33701;
wire     [31:0] n33702;
wire     [31:0] n33703;
wire     [31:0] n33704;
wire     [31:0] n33705;
wire     [31:0] n33706;
wire     [31:0] n33707;
wire     [31:0] n33708;
wire     [31:0] n33709;
wire     [31:0] n33710;
wire     [31:0] n33711;
wire     [31:0] n33712;
wire     [31:0] n33713;
wire     [31:0] n33714;
wire     [31:0] n33715;
wire     [31:0] n33716;
wire     [31:0] n33717;
wire     [31:0] n33718;
wire     [31:0] n33719;
wire     [31:0] n33720;
wire     [31:0] n33721;
wire     [31:0] n33722;
wire     [31:0] n33723;
wire     [31:0] n33724;
wire     [31:0] n33725;
wire     [31:0] n33726;
wire     [31:0] n33727;
wire     [31:0] n33728;
wire     [31:0] n33729;
wire     [31:0] n33730;
wire     [31:0] n33731;
wire     [31:0] n33732;
wire     [31:0] n33733;
wire     [31:0] n33734;
wire     [31:0] n33735;
wire     [31:0] n33736;
wire     [31:0] n33737;
wire     [31:0] n33738;
wire     [31:0] n33739;
wire     [31:0] n33740;
wire     [31:0] n33741;
wire     [31:0] n33742;
wire     [31:0] n33743;
wire     [31:0] n33744;
wire     [31:0] n33745;
wire     [31:0] n33746;
wire     [31:0] n33747;
wire     [31:0] n33748;
wire     [31:0] n33749;
wire     [31:0] n33750;
wire     [31:0] n33751;
wire     [31:0] n33752;
wire     [31:0] n33753;
wire     [31:0] n33754;
wire     [31:0] n33755;
wire     [31:0] n33756;
wire     [31:0] n33757;
wire     [31:0] n33758;
wire     [31:0] n33759;
wire     [31:0] n33760;
wire     [31:0] n33761;
wire     [31:0] n33762;
wire     [31:0] n33763;
wire     [31:0] n33764;
wire     [31:0] n33765;
wire     [31:0] n33766;
wire     [31:0] n33767;
wire     [31:0] n33768;
wire     [31:0] n33769;
wire     [31:0] n33770;
wire     [31:0] n33771;
wire     [31:0] n33772;
wire     [31:0] n33773;
wire     [31:0] n33774;
wire     [31:0] n33775;
wire     [31:0] n33776;
wire     [31:0] n33777;
wire     [31:0] n33778;
wire     [31:0] n33779;
wire     [31:0] n33780;
wire     [31:0] n33781;
wire     [31:0] n33782;
wire     [31:0] n33783;
wire     [31:0] n33784;
wire            n33785;
wire            n33786;
wire            n33787;
wire            n33788;
wire            n33789;
wire            n33790;
wire            n33791;
wire            n33792;
wire            n33793;
wire            n33794;
wire            n33795;
wire            n33796;
wire            n33797;
wire            n33798;
wire            n33799;
wire            n33800;
wire            n33801;
wire            n33802;
wire            n33803;
wire            n33804;
wire            n33805;
wire            n33806;
wire            n33807;
wire            n33808;
wire            n33809;
wire            n33810;
wire            n33811;
wire            n33812;
wire            n33813;
wire            n33814;
wire            n33815;
wire            n33816;
wire            n33817;
wire            n33818;
wire            n33819;
wire            n33820;
wire            n33821;
wire            n33822;
wire            n33823;
wire            n33824;
wire            n33825;
wire            n33826;
wire            n33827;
wire            n33828;
wire            n33829;
wire            n33830;
wire            n33831;
wire            n33832;
wire            n33833;
wire            n33834;
wire            n33835;
wire            n33836;
wire            n33837;
wire            n33838;
wire            n33839;
wire            n33840;
wire            n33841;
wire            n33842;
wire            n33843;
wire            n33844;
wire            n33845;
wire            n33846;
wire            n33847;
wire            n33848;
wire            n33849;
wire            n33850;
wire            n33851;
wire            n33852;
wire            n33853;
wire            n33854;
wire            n33855;
wire            n33856;
wire            n33857;
wire            n33858;
wire            n33859;
wire            n33860;
wire            n33861;
wire            n33862;
wire            n33863;
wire            n33864;
wire            n33865;
wire            n33866;
wire            n33867;
wire            n33868;
wire            n33869;
wire            n33870;
wire            n33871;
wire            n33872;
wire            n33873;
wire            n33874;
wire            n33875;
wire            n33876;
wire            n33877;
wire            n33878;
wire            n33879;
wire            n33880;
wire            n33881;
wire            n33882;
wire            n33883;
wire            n33884;
wire            n33885;
wire            n33886;
wire            n33887;
wire            n33888;
wire            n33889;
wire            n33890;
wire            n33891;
wire            n33892;
wire            n33893;
wire            n33894;
wire            n33895;
wire            n33896;
wire            n33897;
wire            n33898;
wire            n33899;
wire            n33900;
wire            n33901;
wire            n33902;
wire            n33903;
wire            n33904;
wire            n33905;
wire            n33906;
wire            n33907;
wire            n33908;
wire            n33909;
wire            n33910;
wire            n33911;
wire            n33912;
wire            n33913;
wire            n33914;
wire            n33915;
wire            n33916;
wire            n33917;
wire            n33918;
wire            n33919;
wire            n33920;
wire            n33921;
wire            n33922;
wire            n33923;
wire            n33924;
wire            n33925;
wire            n33926;
wire            n33927;
wire            n33928;
wire            n33929;
wire            n33930;
wire            n33931;
wire            n33932;
wire            n33933;
wire            n33934;
wire            n33935;
wire            n33936;
wire            n33937;
wire            n33938;
wire            n33939;
wire            n33940;
wire            n33941;
wire            n33942;
wire            n33943;
wire            n33944;
wire            n33945;
wire            n33946;
wire            n33947;
wire            n33948;
wire            n33949;
wire            n33950;
wire            n33951;
wire            n33952;
wire            n33953;
wire            n33954;
wire            n33955;
wire            n33956;
wire            n33957;
wire            n33958;
wire            n33959;
wire            n33960;
wire            n33961;
wire            n33962;
wire            n33963;
wire            n33964;
wire            n33965;
wire            n33966;
wire            n33967;
wire            n33968;
wire            n33969;
wire            n33970;
wire            n33971;
wire            n33972;
wire            n33973;
wire            n33974;
wire            n33975;
wire            n33976;
wire            n33977;
wire            n33978;
wire            n33979;
wire            n33980;
wire            n33981;
wire            n33982;
wire            n33983;
wire            n33984;
wire            n33985;
wire            n33986;
wire            n33987;
wire            n33988;
wire            n33989;
wire            n33990;
wire            n33991;
wire            n33992;
wire            n33993;
wire            n33994;
wire            n33995;
wire            n33996;
wire            n33997;
wire            n33998;
wire            n33999;
wire            n34000;
wire            n34001;
wire            n34002;
wire            n34003;
wire            n34004;
wire            n34005;
wire            n34006;
wire            n34007;
wire            n34008;
wire            n34009;
wire            n34010;
wire            n34011;
wire            n34012;
wire            n34013;
wire            n34014;
wire            n34015;
wire            n34016;
wire            n34017;
wire            n34018;
wire            n34019;
wire            n34020;
wire            n34021;
wire            n34022;
wire            n34023;
wire            n34024;
wire            n34025;
wire            n34026;
wire            n34027;
wire            n34028;
wire            n34029;
wire            n34030;
wire            n34031;
wire            n34032;
wire            n34033;
wire            n34034;
wire            n34035;
wire            n34036;
wire            n34037;
wire            n34038;
wire            n34039;
wire            n34040;
wire            n34041;
wire            n34042;
wire            n34043;
wire            n34044;
wire            n34045;
wire            n34046;
wire            n34047;
wire            n34048;
wire            n34049;
wire            n34050;
wire            n34051;
wire            n34052;
wire            n34053;
wire            n34054;
wire            n34055;
wire            n34056;
wire            n34057;
wire            n34058;
wire            n34059;
wire            n34060;
wire            n34061;
wire            n34062;
wire            n34063;
wire            n34064;
wire            n34065;
wire            n34066;
wire            n34067;
wire            n34068;
wire            n34069;
wire            n34070;
wire            n34071;
wire            n34072;
wire            n34073;
wire            n34074;
wire            n34075;
wire            n34076;
wire            n34077;
wire            n34078;
wire            n34079;
wire            n34080;
wire            n34081;
wire            n34082;
wire            n34083;
wire            n34084;
wire            n34085;
wire            n34086;
wire            n34087;
wire            n34088;
wire            n34089;
wire            n34090;
wire            n34091;
wire            n34092;
wire            n34093;
wire            n34094;
wire            n34095;
wire            n34096;
wire            n34097;
wire            n34098;
wire            n34099;
wire            n34100;
wire            n34101;
wire            n34102;
wire            n34103;
wire            n34104;
wire            n34105;
wire            n34106;
wire            n34107;
wire            n34108;
wire            n34109;
wire            n34110;
wire            n34111;
wire            n34112;
wire            n34113;
wire            n34114;
wire            n34115;
wire            n34116;
wire            n34117;
wire            n34118;
wire            n34119;
wire            n34120;
wire            n34121;
wire            n34122;
wire            n34123;
wire            n34124;
wire            n34125;
wire            n34126;
wire            n34127;
wire            n34128;
wire            n34129;
wire            n34130;
wire            n34131;
wire            n34132;
wire            n34133;
wire            n34134;
wire            n34135;
wire            n34136;
wire            n34137;
wire            n34138;
wire            n34139;
wire            n34140;
wire            n34141;
wire            n34142;
wire            n34143;
wire            n34144;
wire            n34145;
wire            n34146;
wire            n34147;
wire            n34148;
wire            n34149;
wire            n34150;
wire            n34151;
wire            n34152;
wire            n34153;
wire            n34154;
wire            n34155;
wire            n34156;
wire            n34157;
wire            n34158;
wire            n34159;
wire            n34160;
wire            n34161;
wire            n34162;
wire            n34163;
wire            n34164;
wire            n34165;
wire            n34166;
wire            n34167;
wire            n34168;
wire            n34169;
wire            n34170;
wire            n34171;
wire            n34172;
wire            n34173;
wire            n34174;
wire            n34175;
wire            n34176;
wire            n34177;
wire            n34178;
wire            n34179;
wire            n34180;
wire            n34181;
wire            n34182;
wire            n34183;
wire            n34184;
wire            n34185;
wire            n34186;
wire            n34187;
wire            n34188;
wire            n34189;
wire            n34190;
wire            n34191;
wire            n34192;
wire            n34193;
wire            n34194;
wire            n34195;
wire            n34196;
wire            n34197;
wire            n34198;
wire            n34199;
wire            n34200;
wire            n34201;
wire            n34202;
wire            n34203;
wire            n34204;
wire            n34205;
wire            n34206;
wire            n34207;
wire            n34208;
wire            n34209;
wire            n34210;
wire            n34211;
wire            n34212;
wire            n34213;
wire            n34214;
wire            n34215;
wire            n34216;
wire            n34217;
wire            n34218;
wire            n34219;
wire            n34220;
wire            n34221;
wire            n34222;
wire            n34223;
wire            n34224;
wire            n34225;
wire            n34226;
wire            n34227;
wire            n34228;
wire            n34229;
wire            n34230;
wire            n34231;
wire            n34232;
wire            n34233;
wire            n34234;
wire            n34235;
wire            n34236;
wire            n34237;
wire            n34238;
wire            n34239;
wire            n34240;
wire            n34241;
wire            n34242;
wire            n34243;
wire            n34244;
wire            n34245;
wire            n34246;
wire            n34247;
wire            n34248;
wire            n34249;
wire            n34250;
wire            n34251;
wire            n34252;
wire            n34253;
wire            n34254;
wire            n34255;
wire            n34256;
wire            n34257;
wire            n34258;
wire            n34259;
wire            n34260;
wire            n34261;
wire            n34262;
wire            n34263;
wire            n34264;
wire            n34265;
wire            n34266;
wire            n34267;
wire            n34268;
wire            n34269;
wire            n34270;
wire            n34271;
wire            n34272;
wire            n34273;
wire            n34274;
wire            n34275;
wire            n34276;
wire            n34277;
wire            n34278;
wire            n34279;
wire            n34280;
wire            n34281;
wire            n34282;
wire            n34283;
wire            n34284;
wire            n34285;
wire            n34286;
wire            n34287;
wire            n34288;
wire            n34289;
wire            n34290;
wire            n34291;
wire            n34292;
wire            n34293;
wire            n34294;
wire            n34295;
wire            n34296;
wire     [31:0] n34297;
wire     [31:0] n34298;
wire     [31:0] n34299;
wire     [31:0] n34300;
wire     [31:0] n34301;
wire     [31:0] n34302;
wire     [31:0] n34303;
wire     [31:0] n34304;
wire     [31:0] n34305;
wire     [31:0] n34306;
wire     [31:0] n34307;
wire     [31:0] n34308;
wire     [31:0] n34309;
wire     [31:0] n34310;
wire     [31:0] n34311;
wire     [31:0] n34312;
wire     [31:0] n34313;
wire     [31:0] n34314;
wire     [31:0] n34315;
wire     [31:0] n34316;
wire     [31:0] n34317;
wire     [31:0] n34318;
wire     [31:0] n34319;
wire     [31:0] n34320;
wire     [31:0] n34321;
wire     [31:0] n34322;
wire     [31:0] n34323;
wire     [31:0] n34324;
wire     [31:0] n34325;
wire     [31:0] n34326;
wire     [31:0] n34327;
wire     [31:0] n34328;
wire     [31:0] n34329;
wire     [31:0] n34330;
wire     [31:0] n34331;
wire     [31:0] n34332;
wire     [31:0] n34333;
wire     [31:0] n34334;
wire     [31:0] n34335;
wire     [31:0] n34336;
wire     [31:0] n34337;
wire     [31:0] n34338;
wire     [31:0] n34339;
wire     [31:0] n34340;
wire     [31:0] n34341;
wire     [31:0] n34342;
wire     [31:0] n34343;
wire     [31:0] n34344;
wire     [31:0] n34345;
wire     [31:0] n34346;
wire     [31:0] n34347;
wire     [31:0] n34348;
wire     [31:0] n34349;
wire     [31:0] n34350;
wire     [31:0] n34351;
wire     [31:0] n34352;
wire     [31:0] n34353;
wire     [31:0] n34354;
wire     [31:0] n34355;
wire     [31:0] n34356;
wire     [31:0] n34357;
wire     [31:0] n34358;
wire     [31:0] n34359;
wire     [31:0] n34360;
wire     [31:0] n34361;
wire     [31:0] n34362;
wire     [31:0] n34363;
wire     [31:0] n34364;
wire     [31:0] n34365;
wire     [31:0] n34366;
wire     [31:0] n34367;
wire     [31:0] n34368;
wire     [31:0] n34369;
wire     [31:0] n34370;
wire     [31:0] n34371;
wire     [31:0] n34372;
wire     [31:0] n34373;
wire     [31:0] n34374;
wire     [31:0] n34375;
wire     [31:0] n34376;
wire     [31:0] n34377;
wire     [31:0] n34378;
wire     [31:0] n34379;
wire     [31:0] n34380;
wire     [31:0] n34381;
wire     [31:0] n34382;
wire     [31:0] n34383;
wire     [31:0] n34384;
wire     [31:0] n34385;
wire     [31:0] n34386;
wire     [31:0] n34387;
wire     [31:0] n34388;
wire     [31:0] n34389;
wire     [31:0] n34390;
wire     [31:0] n34391;
wire     [31:0] n34392;
wire     [31:0] n34393;
wire     [31:0] n34394;
wire     [31:0] n34395;
wire     [31:0] n34396;
wire     [31:0] n34397;
wire     [31:0] n34398;
wire     [31:0] n34399;
wire     [31:0] n34400;
wire     [31:0] n34401;
wire     [31:0] n34402;
wire     [31:0] n34403;
wire     [31:0] n34404;
wire     [31:0] n34405;
wire     [31:0] n34406;
wire     [31:0] n34407;
wire     [31:0] n34408;
wire     [31:0] n34409;
wire     [31:0] n34410;
wire     [31:0] n34411;
wire     [31:0] n34412;
wire     [31:0] n34413;
wire     [31:0] n34414;
wire     [31:0] n34415;
wire     [31:0] n34416;
wire     [31:0] n34417;
wire     [31:0] n34418;
wire     [31:0] n34419;
wire     [31:0] n34420;
wire     [31:0] n34421;
wire     [31:0] n34422;
wire     [31:0] n34423;
wire     [31:0] n34424;
wire     [31:0] n34425;
wire     [31:0] n34426;
wire     [31:0] n34427;
wire     [31:0] n34428;
wire     [31:0] n34429;
wire     [31:0] n34430;
wire     [31:0] n34431;
wire     [31:0] n34432;
wire     [31:0] n34433;
wire     [31:0] n34434;
wire     [31:0] n34435;
wire     [31:0] n34436;
wire     [31:0] n34437;
wire     [31:0] n34438;
wire     [31:0] n34439;
wire     [31:0] n34440;
wire     [31:0] n34441;
wire     [31:0] n34442;
wire     [31:0] n34443;
wire     [31:0] n34444;
wire     [31:0] n34445;
wire     [31:0] n34446;
wire     [31:0] n34447;
wire     [31:0] n34448;
wire     [31:0] n34449;
wire     [31:0] n34450;
wire     [31:0] n34451;
wire     [31:0] n34452;
wire     [31:0] n34453;
wire     [31:0] n34454;
wire     [31:0] n34455;
wire     [31:0] n34456;
wire     [31:0] n34457;
wire     [31:0] n34458;
wire     [31:0] n34459;
wire     [31:0] n34460;
wire     [31:0] n34461;
wire     [31:0] n34462;
wire     [31:0] n34463;
wire     [31:0] n34464;
wire     [31:0] n34465;
wire     [31:0] n34466;
wire     [31:0] n34467;
wire     [31:0] n34468;
wire     [31:0] n34469;
wire     [31:0] n34470;
wire     [31:0] n34471;
wire     [31:0] n34472;
wire     [31:0] n34473;
wire     [31:0] n34474;
wire     [31:0] n34475;
wire     [31:0] n34476;
wire     [31:0] n34477;
wire     [31:0] n34478;
wire     [31:0] n34479;
wire     [31:0] n34480;
wire     [31:0] n34481;
wire     [31:0] n34482;
wire     [31:0] n34483;
wire     [31:0] n34484;
wire     [31:0] n34485;
wire     [31:0] n34486;
wire     [31:0] n34487;
wire     [31:0] n34488;
wire     [31:0] n34489;
wire     [31:0] n34490;
wire     [31:0] n34491;
wire     [31:0] n34492;
wire     [31:0] n34493;
wire     [31:0] n34494;
wire     [31:0] n34495;
wire     [31:0] n34496;
wire     [31:0] n34497;
wire     [31:0] n34498;
wire     [31:0] n34499;
wire     [31:0] n34500;
wire     [31:0] n34501;
wire     [31:0] n34502;
wire     [31:0] n34503;
wire     [31:0] n34504;
wire     [31:0] n34505;
wire     [31:0] n34506;
wire     [31:0] n34507;
wire     [31:0] n34508;
wire     [31:0] n34509;
wire     [31:0] n34510;
wire     [31:0] n34511;
wire     [31:0] n34512;
wire     [31:0] n34513;
wire     [31:0] n34514;
wire     [31:0] n34515;
wire     [31:0] n34516;
wire     [31:0] n34517;
wire     [31:0] n34518;
wire     [31:0] n34519;
wire     [31:0] n34520;
wire     [31:0] n34521;
wire     [31:0] n34522;
wire     [31:0] n34523;
wire     [31:0] n34524;
wire     [31:0] n34525;
wire     [31:0] n34526;
wire     [31:0] n34527;
wire     [31:0] n34528;
wire     [31:0] n34529;
wire     [31:0] n34530;
wire     [31:0] n34531;
wire     [31:0] n34532;
wire     [31:0] n34533;
wire     [31:0] n34534;
wire     [31:0] n34535;
wire     [31:0] n34536;
wire     [31:0] n34537;
wire     [31:0] n34538;
wire     [31:0] n34539;
wire     [31:0] n34540;
wire     [31:0] n34541;
wire     [31:0] n34542;
wire     [31:0] n34543;
wire     [31:0] n34544;
wire     [31:0] n34545;
wire     [31:0] n34546;
wire     [31:0] n34547;
wire     [31:0] n34548;
wire     [31:0] n34549;
wire     [31:0] n34550;
wire     [31:0] n34551;
wire     [31:0] n34552;
wire     [31:0] n34553;
wire     [31:0] n34554;
wire     [31:0] n34555;
wire     [31:0] n34556;
wire     [31:0] n34557;
wire     [31:0] n34558;
wire     [31:0] n34559;
wire     [31:0] n34560;
wire     [31:0] n34561;
wire     [31:0] n34562;
wire     [31:0] n34563;
wire     [31:0] n34564;
wire     [31:0] n34565;
wire     [31:0] n34566;
wire     [31:0] n34567;
wire     [31:0] n34568;
wire     [31:0] n34569;
wire     [31:0] n34570;
wire     [31:0] n34571;
wire     [31:0] n34572;
wire     [31:0] n34573;
wire     [31:0] n34574;
wire     [31:0] n34575;
wire     [31:0] n34576;
wire     [31:0] n34577;
wire     [31:0] n34578;
wire     [31:0] n34579;
wire     [31:0] n34580;
wire     [31:0] n34581;
wire     [31:0] n34582;
wire     [31:0] n34583;
wire     [31:0] n34584;
wire     [31:0] n34585;
wire     [31:0] n34586;
wire     [31:0] n34587;
wire     [31:0] n34588;
wire     [31:0] n34589;
wire     [31:0] n34590;
wire     [31:0] n34591;
wire     [31:0] n34592;
wire     [31:0] n34593;
wire     [31:0] n34594;
wire     [31:0] n34595;
wire     [31:0] n34596;
wire     [31:0] n34597;
wire     [31:0] n34598;
wire     [31:0] n34599;
wire     [31:0] n34600;
wire     [31:0] n34601;
wire     [31:0] n34602;
wire     [31:0] n34603;
wire     [31:0] n34604;
wire     [31:0] n34605;
wire     [31:0] n34606;
wire     [31:0] n34607;
wire     [31:0] n34608;
wire     [31:0] n34609;
wire     [31:0] n34610;
wire     [31:0] n34611;
wire     [31:0] n34612;
wire     [31:0] n34613;
wire     [31:0] n34614;
wire     [31:0] n34615;
wire     [31:0] n34616;
wire     [31:0] n34617;
wire     [31:0] n34618;
wire     [31:0] n34619;
wire     [31:0] n34620;
wire     [31:0] n34621;
wire     [31:0] n34622;
wire     [31:0] n34623;
wire     [31:0] n34624;
wire     [31:0] n34625;
wire     [31:0] n34626;
wire     [31:0] n34627;
wire     [31:0] n34628;
wire     [31:0] n34629;
wire     [31:0] n34630;
wire     [31:0] n34631;
wire     [31:0] n34632;
wire     [31:0] n34633;
wire     [31:0] n34634;
wire     [31:0] n34635;
wire     [31:0] n34636;
wire     [31:0] n34637;
wire     [31:0] n34638;
wire     [31:0] n34639;
wire     [31:0] n34640;
wire     [31:0] n34641;
wire     [31:0] n34642;
wire     [31:0] n34643;
wire     [31:0] n34644;
wire     [31:0] n34645;
wire     [31:0] n34646;
wire     [31:0] n34647;
wire     [31:0] n34648;
wire     [31:0] n34649;
wire     [31:0] n34650;
wire     [31:0] n34651;
wire     [31:0] n34652;
wire     [31:0] n34653;
wire     [31:0] n34654;
wire     [31:0] n34655;
wire     [31:0] n34656;
wire     [31:0] n34657;
wire     [31:0] n34658;
wire     [31:0] n34659;
wire     [31:0] n34660;
wire     [31:0] n34661;
wire     [31:0] n34662;
wire     [31:0] n34663;
wire     [31:0] n34664;
wire     [31:0] n34665;
wire     [31:0] n34666;
wire     [31:0] n34667;
wire     [31:0] n34668;
wire     [31:0] n34669;
wire     [31:0] n34670;
wire     [31:0] n34671;
wire     [31:0] n34672;
wire     [31:0] n34673;
wire     [31:0] n34674;
wire     [31:0] n34675;
wire     [31:0] n34676;
wire     [31:0] n34677;
wire     [31:0] n34678;
wire     [31:0] n34679;
wire     [31:0] n34680;
wire     [31:0] n34681;
wire     [31:0] n34682;
wire     [31:0] n34683;
wire     [31:0] n34684;
wire     [31:0] n34685;
wire     [31:0] n34686;
wire     [31:0] n34687;
wire     [31:0] n34688;
wire     [31:0] n34689;
wire     [31:0] n34690;
wire     [31:0] n34691;
wire     [31:0] n34692;
wire     [31:0] n34693;
wire     [31:0] n34694;
wire     [31:0] n34695;
wire     [31:0] n34696;
wire     [31:0] n34697;
wire     [31:0] n34698;
wire     [31:0] n34699;
wire     [31:0] n34700;
wire     [31:0] n34701;
wire     [31:0] n34702;
wire     [31:0] n34703;
wire     [31:0] n34704;
wire     [31:0] n34705;
wire     [31:0] n34706;
wire     [31:0] n34707;
wire     [31:0] n34708;
wire     [31:0] n34709;
wire     [31:0] n34710;
wire     [31:0] n34711;
wire     [31:0] n34712;
wire     [31:0] n34713;
wire     [31:0] n34714;
wire     [31:0] n34715;
wire     [31:0] n34716;
wire     [31:0] n34717;
wire     [31:0] n34718;
wire     [31:0] n34719;
wire     [31:0] n34720;
wire     [31:0] n34721;
wire     [31:0] n34722;
wire     [31:0] n34723;
wire     [31:0] n34724;
wire     [31:0] n34725;
wire     [31:0] n34726;
wire     [31:0] n34727;
wire     [31:0] n34728;
wire     [31:0] n34729;
wire     [31:0] n34730;
wire     [31:0] n34731;
wire     [31:0] n34732;
wire     [31:0] n34733;
wire     [31:0] n34734;
wire     [31:0] n34735;
wire     [31:0] n34736;
wire     [31:0] n34737;
wire     [31:0] n34738;
wire     [31:0] n34739;
wire     [31:0] n34740;
wire     [31:0] n34741;
wire     [31:0] n34742;
wire     [31:0] n34743;
wire     [31:0] n34744;
wire     [31:0] n34745;
wire     [31:0] n34746;
wire     [31:0] n34747;
wire     [31:0] n34748;
wire     [31:0] n34749;
wire     [31:0] n34750;
wire     [31:0] n34751;
wire     [31:0] n34752;
wire     [31:0] n34753;
wire     [31:0] n34754;
wire     [31:0] n34755;
wire     [31:0] n34756;
wire     [31:0] n34757;
wire     [31:0] n34758;
wire     [31:0] n34759;
wire     [31:0] n34760;
wire     [31:0] n34761;
wire     [31:0] n34762;
wire     [31:0] n34763;
wire     [31:0] n34764;
wire     [31:0] n34765;
wire     [31:0] n34766;
wire     [31:0] n34767;
wire     [31:0] n34768;
wire     [31:0] n34769;
wire     [31:0] n34770;
wire     [31:0] n34771;
wire     [31:0] n34772;
wire     [31:0] n34773;
wire     [31:0] n34774;
wire     [31:0] n34775;
wire     [31:0] n34776;
wire     [31:0] n34777;
wire     [31:0] n34778;
wire     [31:0] n34779;
wire     [31:0] n34780;
wire     [31:0] n34781;
wire     [31:0] n34782;
wire     [31:0] n34783;
wire     [31:0] n34784;
wire     [31:0] n34785;
wire     [31:0] n34786;
wire     [31:0] n34787;
wire     [31:0] n34788;
wire     [31:0] n34789;
wire     [31:0] n34790;
wire     [31:0] n34791;
wire     [31:0] n34792;
wire     [31:0] n34793;
wire     [31:0] n34794;
wire     [31:0] n34795;
wire     [31:0] n34796;
wire     [31:0] n34797;
wire     [31:0] n34798;
wire     [31:0] n34799;
wire     [31:0] n34800;
wire     [31:0] n34801;
wire     [31:0] n34802;
wire     [31:0] n34803;
wire     [31:0] n34804;
wire     [31:0] n34805;
wire     [31:0] n34806;
wire     [31:0] n34807;
wire     [31:0] n34808;
wire     [31:0] n34809;
wire     [31:0] n34810;
wire     [31:0] n34811;
wire     [31:0] n34812;
wire     [31:0] n34813;
wire     [31:0] n34814;
wire     [31:0] n34815;
wire     [31:0] n34816;
wire     [31:0] n34817;
wire     [31:0] n34818;
wire            n34819;
wire            n34820;
wire     [31:0] n34821;
wire     [31:0] n34822;
wire     [31:0] n34823;
wire     [31:0] n34824;
wire     [31:0] n34825;
wire     [31:0] n34826;
wire     [31:0] n34827;
wire     [31:0] n34828;
wire     [31:0] n34829;
wire     [31:0] n34830;
wire     [31:0] n34831;
wire     [31:0] n34832;
wire     [31:0] n34833;
wire     [31:0] n34834;
wire     [31:0] n34835;
wire     [31:0] n34836;
wire     [31:0] n34837;
wire     [31:0] n34838;
wire     [31:0] n34839;
wire     [31:0] n34840;
wire     [31:0] n34841;
wire     [31:0] n34842;
wire     [31:0] n34843;
wire     [31:0] n34844;
wire     [31:0] n34845;
wire     [31:0] n34846;
wire     [31:0] n34847;
wire     [31:0] n34848;
wire     [31:0] n34849;
wire     [31:0] n34850;
wire     [31:0] n34851;
wire     [31:0] n34852;
wire     [31:0] n34853;
wire     [31:0] n34854;
wire     [31:0] n34855;
wire     [31:0] n34856;
wire     [31:0] n34857;
wire     [31:0] n34858;
wire     [31:0] n34859;
wire     [31:0] n34860;
wire     [31:0] n34861;
wire     [31:0] n34862;
wire     [31:0] n34863;
wire     [31:0] n34864;
wire     [31:0] n34865;
wire     [31:0] n34866;
wire     [31:0] n34867;
wire     [31:0] n34868;
wire     [31:0] n34869;
wire     [31:0] n34870;
wire     [31:0] n34871;
wire     [31:0] n34872;
wire     [31:0] n34873;
wire     [31:0] n34874;
wire     [31:0] n34875;
wire     [31:0] n34876;
wire     [31:0] n34877;
wire     [31:0] n34878;
wire     [31:0] n34879;
wire     [31:0] n34880;
wire     [31:0] n34881;
wire     [31:0] n34882;
wire     [31:0] n34883;
wire     [31:0] n34884;
wire     [31:0] n34885;
wire     [31:0] n34886;
wire     [31:0] n34887;
wire     [31:0] n34888;
wire     [31:0] n34889;
wire     [31:0] n34890;
wire     [31:0] n34891;
wire     [31:0] n34892;
wire     [31:0] n34893;
wire     [31:0] n34894;
wire     [31:0] n34895;
wire     [31:0] n34896;
wire     [31:0] n34897;
wire     [31:0] n34898;
wire     [31:0] n34899;
wire     [31:0] n34900;
wire     [31:0] n34901;
wire     [31:0] n34902;
wire     [31:0] n34903;
wire     [31:0] n34904;
wire     [31:0] n34905;
wire     [31:0] n34906;
wire     [31:0] n34907;
wire     [31:0] n34908;
wire     [31:0] n34909;
wire     [31:0] n34910;
wire     [31:0] n34911;
wire     [31:0] n34912;
wire     [31:0] n34913;
wire     [31:0] n34914;
wire     [31:0] n34915;
wire     [31:0] n34916;
wire     [31:0] n34917;
wire     [31:0] n34918;
wire     [31:0] n34919;
wire     [31:0] n34920;
wire     [31:0] n34921;
wire     [31:0] n34922;
wire     [31:0] n34923;
wire     [31:0] n34924;
wire     [31:0] n34925;
wire     [31:0] n34926;
wire     [31:0] n34927;
wire     [31:0] n34928;
wire     [31:0] n34929;
wire     [31:0] n34930;
wire     [31:0] n34931;
wire     [31:0] n34932;
wire     [31:0] n34933;
wire     [31:0] n34934;
wire     [31:0] n34935;
wire     [31:0] n34936;
wire     [31:0] n34937;
wire     [31:0] n34938;
wire     [31:0] n34939;
wire     [31:0] n34940;
wire     [31:0] n34941;
wire     [31:0] n34942;
wire     [31:0] n34943;
wire     [31:0] n34944;
wire     [31:0] n34945;
wire     [31:0] n34946;
wire     [31:0] n34947;
wire     [31:0] n34948;
wire     [31:0] n34949;
wire     [31:0] n34950;
wire     [31:0] n34951;
wire     [31:0] n34952;
wire     [31:0] n34953;
wire     [31:0] n34954;
wire     [31:0] n34955;
wire     [31:0] n34956;
wire     [31:0] n34957;
wire     [31:0] n34958;
wire     [31:0] n34959;
wire     [31:0] n34960;
wire     [31:0] n34961;
wire     [31:0] n34962;
wire     [31:0] n34963;
wire     [31:0] n34964;
wire     [31:0] n34965;
wire     [31:0] n34966;
wire     [31:0] n34967;
wire     [31:0] n34968;
wire     [31:0] n34969;
wire     [31:0] n34970;
wire     [31:0] n34971;
wire     [31:0] n34972;
wire     [31:0] n34973;
wire     [31:0] n34974;
wire     [31:0] n34975;
wire     [31:0] n34976;
wire     [31:0] n34977;
wire     [31:0] n34978;
wire     [31:0] n34979;
wire     [31:0] n34980;
wire     [31:0] n34981;
wire     [31:0] n34982;
wire     [31:0] n34983;
wire     [31:0] n34984;
wire     [31:0] n34985;
wire     [31:0] n34986;
wire     [31:0] n34987;
wire     [31:0] n34988;
wire     [31:0] n34989;
wire     [31:0] n34990;
wire     [31:0] n34991;
wire     [31:0] n34992;
wire     [31:0] n34993;
wire     [31:0] n34994;
wire     [31:0] n34995;
wire     [31:0] n34996;
wire     [31:0] n34997;
wire     [31:0] n34998;
wire     [31:0] n34999;
wire     [31:0] n35000;
wire     [31:0] n35001;
wire     [31:0] n35002;
wire     [31:0] n35003;
wire     [31:0] n35004;
wire     [31:0] n35005;
wire     [31:0] n35006;
wire     [31:0] n35007;
wire     [31:0] n35008;
wire     [31:0] n35009;
wire     [31:0] n35010;
wire     [31:0] n35011;
wire     [31:0] n35012;
wire     [31:0] n35013;
wire     [31:0] n35014;
wire     [31:0] n35015;
wire     [31:0] n35016;
wire     [31:0] n35017;
wire     [31:0] n35018;
wire     [31:0] n35019;
wire     [31:0] n35020;
wire     [31:0] n35021;
wire     [31:0] n35022;
wire     [31:0] n35023;
wire     [31:0] n35024;
wire     [31:0] n35025;
wire     [31:0] n35026;
wire     [31:0] n35027;
wire     [31:0] n35028;
wire     [31:0] n35029;
wire     [31:0] n35030;
wire     [31:0] n35031;
wire     [31:0] n35032;
wire     [31:0] n35033;
wire     [31:0] n35034;
wire     [31:0] n35035;
wire     [31:0] n35036;
wire     [31:0] n35037;
wire     [31:0] n35038;
wire     [31:0] n35039;
wire     [31:0] n35040;
wire     [31:0] n35041;
wire     [31:0] n35042;
wire     [31:0] n35043;
wire     [31:0] n35044;
wire     [31:0] n35045;
wire     [31:0] n35046;
wire     [31:0] n35047;
wire     [31:0] n35048;
wire     [31:0] n35049;
wire     [31:0] n35050;
wire     [31:0] n35051;
wire     [31:0] n35052;
wire     [31:0] n35053;
wire     [31:0] n35054;
wire     [31:0] n35055;
wire     [31:0] n35056;
wire     [31:0] n35057;
wire     [31:0] n35058;
wire     [31:0] n35059;
wire     [31:0] n35060;
wire     [31:0] n35061;
wire     [31:0] n35062;
wire     [31:0] n35063;
wire     [31:0] n35064;
wire     [31:0] n35065;
wire     [31:0] n35066;
wire     [31:0] n35067;
wire     [31:0] n35068;
wire     [31:0] n35069;
wire     [31:0] n35070;
wire     [31:0] n35071;
wire     [31:0] n35072;
wire     [31:0] n35073;
wire     [31:0] n35074;
wire     [31:0] n35075;
wire     [31:0] n35076;
wire     [31:0] n35077;
wire     [31:0] n35078;
wire     [31:0] n35079;
wire     [31:0] n35080;
wire     [31:0] n35081;
wire     [31:0] n35082;
wire     [31:0] n35083;
wire     [31:0] n35084;
wire     [31:0] n35085;
wire     [31:0] n35086;
wire     [31:0] n35087;
wire     [31:0] n35088;
wire     [31:0] n35089;
wire     [31:0] n35090;
wire     [31:0] n35091;
wire     [31:0] n35092;
wire     [31:0] n35093;
wire     [31:0] n35094;
wire     [31:0] n35095;
wire     [31:0] n35096;
wire     [31:0] n35097;
wire     [31:0] n35098;
wire     [31:0] n35099;
wire     [31:0] n35100;
wire     [31:0] n35101;
wire     [31:0] n35102;
wire     [31:0] n35103;
wire     [31:0] n35104;
wire     [31:0] n35105;
wire     [31:0] n35106;
wire     [31:0] n35107;
wire     [31:0] n35108;
wire     [31:0] n35109;
wire     [31:0] n35110;
wire     [31:0] n35111;
wire     [31:0] n35112;
wire     [31:0] n35113;
wire     [31:0] n35114;
wire     [31:0] n35115;
wire     [31:0] n35116;
wire     [31:0] n35117;
wire     [31:0] n35118;
wire     [31:0] n35119;
wire     [31:0] n35120;
wire     [31:0] n35121;
wire     [31:0] n35122;
wire     [31:0] n35123;
wire     [31:0] n35124;
wire     [31:0] n35125;
wire     [31:0] n35126;
wire     [31:0] n35127;
wire     [31:0] n35128;
wire     [31:0] n35129;
wire     [31:0] n35130;
wire     [31:0] n35131;
wire     [31:0] n35132;
wire     [31:0] n35133;
wire     [31:0] n35134;
wire     [31:0] n35135;
wire     [31:0] n35136;
wire     [31:0] n35137;
wire     [31:0] n35138;
wire     [31:0] n35139;
wire     [31:0] n35140;
wire     [31:0] n35141;
wire     [31:0] n35142;
wire     [31:0] n35143;
wire     [31:0] n35144;
wire     [31:0] n35145;
wire     [31:0] n35146;
wire     [31:0] n35147;
wire     [31:0] n35148;
wire     [31:0] n35149;
wire     [31:0] n35150;
wire     [31:0] n35151;
wire     [31:0] n35152;
wire     [31:0] n35153;
wire     [31:0] n35154;
wire     [31:0] n35155;
wire     [31:0] n35156;
wire     [31:0] n35157;
wire     [31:0] n35158;
wire     [31:0] n35159;
wire     [31:0] n35160;
wire     [31:0] n35161;
wire     [31:0] n35162;
wire     [31:0] n35163;
wire     [31:0] n35164;
wire     [31:0] n35165;
wire     [31:0] n35166;
wire     [31:0] n35167;
wire     [31:0] n35168;
wire     [31:0] n35169;
wire     [31:0] n35170;
wire     [31:0] n35171;
wire     [31:0] n35172;
wire     [31:0] n35173;
wire     [31:0] n35174;
wire     [31:0] n35175;
wire     [31:0] n35176;
wire     [31:0] n35177;
wire     [31:0] n35178;
wire     [31:0] n35179;
wire     [31:0] n35180;
wire     [31:0] n35181;
wire     [31:0] n35182;
wire     [31:0] n35183;
wire     [31:0] n35184;
wire     [31:0] n35185;
wire     [31:0] n35186;
wire     [31:0] n35187;
wire     [31:0] n35188;
wire     [31:0] n35189;
wire     [31:0] n35190;
wire     [31:0] n35191;
wire     [31:0] n35192;
wire     [31:0] n35193;
wire     [31:0] n35194;
wire     [31:0] n35195;
wire     [31:0] n35196;
wire     [31:0] n35197;
wire     [31:0] n35198;
wire     [31:0] n35199;
wire     [31:0] n35200;
wire     [31:0] n35201;
wire     [31:0] n35202;
wire     [31:0] n35203;
wire     [31:0] n35204;
wire     [31:0] n35205;
wire     [31:0] n35206;
wire     [31:0] n35207;
wire     [31:0] n35208;
wire     [31:0] n35209;
wire     [31:0] n35210;
wire     [31:0] n35211;
wire     [31:0] n35212;
wire     [31:0] n35213;
wire     [31:0] n35214;
wire     [31:0] n35215;
wire     [31:0] n35216;
wire     [31:0] n35217;
wire     [31:0] n35218;
wire     [31:0] n35219;
wire     [31:0] n35220;
wire     [31:0] n35221;
wire     [31:0] n35222;
wire     [31:0] n35223;
wire     [31:0] n35224;
wire     [31:0] n35225;
wire     [31:0] n35226;
wire     [31:0] n35227;
wire     [31:0] n35228;
wire     [31:0] n35229;
wire     [31:0] n35230;
wire     [31:0] n35231;
wire     [31:0] n35232;
wire     [31:0] n35233;
wire     [31:0] n35234;
wire     [31:0] n35235;
wire     [31:0] n35236;
wire     [31:0] n35237;
wire     [31:0] n35238;
wire     [31:0] n35239;
wire     [31:0] n35240;
wire     [31:0] n35241;
wire     [31:0] n35242;
wire     [31:0] n35243;
wire     [31:0] n35244;
wire     [31:0] n35245;
wire     [31:0] n35246;
wire     [31:0] n35247;
wire     [31:0] n35248;
wire     [31:0] n35249;
wire     [31:0] n35250;
wire     [31:0] n35251;
wire     [31:0] n35252;
wire     [31:0] n35253;
wire     [31:0] n35254;
wire     [31:0] n35255;
wire     [31:0] n35256;
wire     [31:0] n35257;
wire     [31:0] n35258;
wire     [31:0] n35259;
wire     [31:0] n35260;
wire     [31:0] n35261;
wire     [31:0] n35262;
wire     [31:0] n35263;
wire     [31:0] n35264;
wire     [31:0] n35265;
wire     [31:0] n35266;
wire     [31:0] n35267;
wire     [31:0] n35268;
wire     [31:0] n35269;
wire     [31:0] n35270;
wire     [31:0] n35271;
wire     [31:0] n35272;
wire     [31:0] n35273;
wire     [31:0] n35274;
wire     [31:0] n35275;
wire     [31:0] n35276;
wire     [31:0] n35277;
wire     [31:0] n35278;
wire     [31:0] n35279;
wire     [31:0] n35280;
wire     [31:0] n35281;
wire     [31:0] n35282;
wire     [31:0] n35283;
wire     [31:0] n35284;
wire     [31:0] n35285;
wire     [31:0] n35286;
wire     [31:0] n35287;
wire     [31:0] n35288;
wire     [31:0] n35289;
wire     [31:0] n35290;
wire     [31:0] n35291;
wire     [31:0] n35292;
wire     [31:0] n35293;
wire     [31:0] n35294;
wire     [31:0] n35295;
wire     [31:0] n35296;
wire     [31:0] n35297;
wire     [31:0] n35298;
wire     [31:0] n35299;
wire     [31:0] n35300;
wire     [31:0] n35301;
wire     [31:0] n35302;
wire     [31:0] n35303;
wire     [31:0] n35304;
wire     [31:0] n35305;
wire     [31:0] n35306;
wire     [31:0] n35307;
wire     [31:0] n35308;
wire     [31:0] n35309;
wire     [31:0] n35310;
wire     [31:0] n35311;
wire     [31:0] n35312;
wire     [31:0] n35313;
wire     [31:0] n35314;
wire     [31:0] n35315;
wire     [31:0] n35316;
wire     [31:0] n35317;
wire     [31:0] n35318;
wire     [31:0] n35319;
wire     [31:0] n35320;
wire     [31:0] n35321;
wire     [31:0] n35322;
wire     [31:0] n35323;
wire     [31:0] n35324;
wire     [31:0] n35325;
wire     [31:0] n35326;
wire     [31:0] n35327;
wire     [31:0] n35328;
wire     [31:0] n35329;
wire     [31:0] n35330;
wire     [31:0] n35331;
wire     [31:0] n35332;
wire     [31:0] n35333;
wire     [31:0] n35334;
wire     [31:0] n35335;
wire     [31:0] n35336;
wire     [31:0] n35337;
wire     [31:0] n35338;
wire     [31:0] n35339;
wire     [31:0] n35340;
wire     [31:0] n35341;
wire     [31:0] n35342;
wire     [31:0] n35343;
wire     [31:0] n35344;
wire     [31:0] n35345;
wire     [31:0] n35346;
wire     [31:0] n35347;
wire     [31:0] n35348;
wire     [31:0] n35349;
wire     [31:0] n35350;
wire     [31:0] n35351;
wire     [31:0] n35352;
wire     [31:0] n35353;
wire     [31:0] n35354;
wire     [31:0] n35355;
wire     [31:0] n35356;
wire     [31:0] n35357;
wire     [31:0] n35358;
wire     [31:0] n35359;
wire     [31:0] n35360;
wire     [31:0] n35361;
wire     [31:0] n35362;
wire     [31:0] n35363;
wire     [31:0] n35364;
wire     [31:0] n35365;
wire     [31:0] n35366;
wire     [31:0] n35367;
wire     [31:0] n35368;
wire     [31:0] n35369;
wire     [31:0] n35370;
wire     [31:0] n35371;
wire     [31:0] n35372;
wire     [31:0] n35373;
wire     [31:0] n35374;
wire     [31:0] n35375;
wire     [31:0] n35376;
wire     [31:0] n35377;
wire     [31:0] n35378;
wire     [31:0] n35379;
wire     [31:0] n35380;
wire     [31:0] n35381;
wire     [31:0] n35382;
wire     [31:0] n35383;
wire     [31:0] n35384;
wire     [31:0] n35385;
wire     [31:0] n35386;
wire     [31:0] n35387;
wire     [31:0] n35388;
wire     [31:0] n35389;
wire     [31:0] n35390;
wire     [31:0] n35391;
wire     [31:0] n35392;
wire     [31:0] n35393;
wire     [31:0] n35394;
wire     [31:0] n35395;
wire     [31:0] n35396;
wire     [31:0] n35397;
wire     [31:0] n35398;
wire     [31:0] n35399;
wire     [31:0] n35400;
wire     [31:0] n35401;
wire     [31:0] n35402;
wire     [31:0] n35403;
wire     [31:0] n35404;
wire     [31:0] n35405;
wire     [31:0] n35406;
wire     [31:0] n35407;
wire     [31:0] n35408;
wire     [31:0] n35409;
wire     [31:0] n35410;
wire     [31:0] n35411;
wire     [31:0] n35412;
wire     [31:0] n35413;
wire     [31:0] n35414;
wire     [31:0] n35415;
wire     [31:0] n35416;
wire     [31:0] n35417;
wire     [31:0] n35418;
wire     [31:0] n35419;
wire     [31:0] n35420;
wire     [31:0] n35421;
wire     [31:0] n35422;
wire     [31:0] n35423;
wire     [31:0] n35424;
wire     [31:0] n35425;
wire     [31:0] n35426;
wire     [31:0] n35427;
wire     [31:0] n35428;
wire     [31:0] n35429;
wire     [31:0] n35430;
wire     [31:0] n35431;
wire     [31:0] n35432;
wire     [31:0] n35433;
wire     [31:0] n35434;
wire     [31:0] n35435;
wire     [31:0] n35436;
wire     [31:0] n35437;
wire     [31:0] n35438;
wire     [31:0] n35439;
wire     [31:0] n35440;
wire     [31:0] n35441;
wire     [31:0] n35442;
wire     [31:0] n35443;
wire     [31:0] n35444;
wire     [31:0] n35445;
wire     [31:0] n35446;
wire     [31:0] n35447;
wire     [31:0] n35448;
wire     [31:0] n35449;
wire     [31:0] n35450;
wire     [31:0] n35451;
wire     [31:0] n35452;
wire     [31:0] n35453;
wire     [31:0] n35454;
wire     [31:0] n35455;
wire     [31:0] n35456;
wire     [31:0] n35457;
wire     [31:0] n35458;
wire     [31:0] n35459;
wire     [31:0] n35460;
wire     [31:0] n35461;
wire     [31:0] n35462;
wire     [31:0] n35463;
wire     [31:0] n35464;
wire     [31:0] n35465;
wire     [31:0] n35466;
wire     [31:0] n35467;
wire     [31:0] n35468;
wire     [31:0] n35469;
wire     [31:0] n35470;
wire     [31:0] n35471;
wire     [31:0] n35472;
wire     [31:0] n35473;
wire     [31:0] n35474;
wire     [31:0] n35475;
wire     [31:0] n35476;
wire     [31:0] n35477;
wire     [31:0] n35478;
wire     [31:0] n35479;
wire     [31:0] n35480;
wire     [31:0] n35481;
wire     [31:0] n35482;
wire     [31:0] n35483;
wire     [31:0] n35484;
wire     [31:0] n35485;
wire     [31:0] n35486;
wire     [31:0] n35487;
wire     [31:0] n35488;
wire     [31:0] n35489;
wire     [31:0] n35490;
wire     [31:0] n35491;
wire     [31:0] n35492;
wire     [31:0] n35493;
wire     [31:0] n35494;
wire     [31:0] n35495;
wire     [31:0] n35496;
wire     [31:0] n35497;
wire     [31:0] n35498;
wire     [31:0] n35499;
wire     [31:0] n35500;
wire     [31:0] n35501;
wire     [31:0] n35502;
wire     [31:0] n35503;
wire     [31:0] n35504;
wire     [31:0] n35505;
wire     [31:0] n35506;
wire     [31:0] n35507;
wire     [31:0] n35508;
wire     [31:0] n35509;
wire     [31:0] n35510;
wire     [31:0] n35511;
wire     [31:0] n35512;
wire     [31:0] n35513;
wire     [31:0] n35514;
wire     [31:0] n35515;
wire     [31:0] n35516;
wire     [31:0] n35517;
wire     [31:0] n35518;
wire     [31:0] n35519;
wire     [31:0] n35520;
wire     [31:0] n35521;
wire     [31:0] n35522;
wire     [31:0] n35523;
wire     [31:0] n35524;
wire     [31:0] n35525;
wire     [31:0] n35526;
wire     [31:0] n35527;
wire     [31:0] n35528;
wire     [31:0] n35529;
wire     [31:0] n35530;
wire     [31:0] n35531;
wire     [31:0] n35532;
wire     [31:0] n35533;
wire     [31:0] n35534;
wire     [31:0] n35535;
wire     [31:0] n35536;
wire     [31:0] n35537;
wire     [31:0] n35538;
wire     [31:0] n35539;
wire     [31:0] n35540;
wire     [31:0] n35541;
wire     [31:0] n35542;
wire     [31:0] n35543;
wire     [31:0] n35544;
wire     [31:0] n35545;
wire     [31:0] n35546;
wire     [31:0] n35547;
wire     [31:0] n35548;
wire     [31:0] n35549;
wire     [31:0] n35550;
wire     [31:0] n35551;
wire     [31:0] n35552;
wire     [31:0] n35553;
wire     [31:0] n35554;
wire     [31:0] n35555;
wire     [31:0] n35556;
wire     [31:0] n35557;
wire     [31:0] n35558;
wire     [31:0] n35559;
wire     [31:0] n35560;
wire     [31:0] n35561;
wire     [31:0] n35562;
wire     [31:0] n35563;
wire     [31:0] n35564;
wire     [31:0] n35565;
wire     [31:0] n35566;
wire     [31:0] n35567;
wire     [31:0] n35568;
wire     [31:0] n35569;
wire     [31:0] n35570;
wire     [31:0] n35571;
wire     [31:0] n35572;
wire     [31:0] n35573;
wire     [31:0] n35574;
wire     [31:0] n35575;
wire     [31:0] n35576;
wire     [31:0] n35577;
wire     [31:0] n35578;
wire     [31:0] n35579;
wire     [31:0] n35580;
wire     [31:0] n35581;
wire     [31:0] n35582;
wire     [31:0] n35583;
wire     [31:0] n35584;
wire     [31:0] n35585;
wire     [31:0] n35586;
wire     [31:0] n35587;
wire     [31:0] n35588;
wire     [31:0] n35589;
wire     [31:0] n35590;
wire     [31:0] n35591;
wire     [31:0] n35592;
wire     [31:0] n35593;
wire     [31:0] n35594;
wire     [31:0] n35595;
wire     [31:0] n35596;
wire     [31:0] n35597;
wire     [31:0] n35598;
wire     [31:0] n35599;
wire     [31:0] n35600;
wire     [31:0] n35601;
wire     [31:0] n35602;
wire     [31:0] n35603;
wire     [31:0] n35604;
wire     [31:0] n35605;
wire     [31:0] n35606;
wire     [31:0] n35607;
wire     [31:0] n35608;
wire     [31:0] n35609;
wire     [31:0] n35610;
wire     [31:0] n35611;
wire     [31:0] n35612;
wire     [31:0] n35613;
wire     [31:0] n35614;
wire     [31:0] n35615;
wire     [31:0] n35616;
wire     [31:0] n35617;
wire     [31:0] n35618;
wire     [31:0] n35619;
wire     [31:0] n35620;
wire     [31:0] n35621;
wire     [31:0] n35622;
wire     [31:0] n35623;
wire     [31:0] n35624;
wire     [31:0] n35625;
wire     [31:0] n35626;
wire     [31:0] n35627;
wire     [31:0] n35628;
wire     [31:0] n35629;
wire     [31:0] n35630;
wire     [31:0] n35631;
wire     [31:0] n35632;
wire     [31:0] n35633;
wire     [31:0] n35634;
wire     [31:0] n35635;
wire     [31:0] n35636;
wire     [31:0] n35637;
wire     [31:0] n35638;
wire     [31:0] n35639;
wire     [31:0] n35640;
wire     [31:0] n35641;
wire     [31:0] n35642;
wire     [31:0] n35643;
wire     [31:0] n35644;
wire     [31:0] n35645;
wire     [31:0] n35646;
wire     [31:0] n35647;
wire     [31:0] n35648;
wire     [31:0] n35649;
wire     [31:0] n35650;
wire     [31:0] n35651;
wire     [31:0] n35652;
wire     [31:0] n35653;
wire     [31:0] n35654;
wire     [31:0] n35655;
wire     [31:0] n35656;
wire     [31:0] n35657;
wire     [31:0] n35658;
wire     [31:0] n35659;
wire     [31:0] n35660;
wire     [31:0] n35661;
wire     [31:0] n35662;
wire     [31:0] n35663;
wire     [31:0] n35664;
wire     [31:0] n35665;
wire     [31:0] n35666;
wire     [31:0] n35667;
wire     [31:0] n35668;
wire     [31:0] n35669;
wire     [31:0] n35670;
wire     [31:0] n35671;
wire     [31:0] n35672;
wire     [31:0] n35673;
wire     [31:0] n35674;
wire     [31:0] n35675;
wire     [31:0] n35676;
wire     [31:0] n35677;
wire     [31:0] n35678;
wire     [31:0] n35679;
wire     [31:0] n35680;
wire     [31:0] n35681;
wire     [31:0] n35682;
wire     [31:0] n35683;
wire     [31:0] n35684;
wire     [31:0] n35685;
wire     [31:0] n35686;
wire     [31:0] n35687;
wire     [31:0] n35688;
wire     [31:0] n35689;
wire     [31:0] n35690;
wire     [31:0] n35691;
wire     [31:0] n35692;
wire     [31:0] n35693;
wire     [31:0] n35694;
wire     [31:0] n35695;
wire     [31:0] n35696;
wire     [31:0] n35697;
wire     [31:0] n35698;
wire     [31:0] n35699;
wire     [31:0] n35700;
wire     [31:0] n35701;
wire     [31:0] n35702;
wire     [31:0] n35703;
wire     [31:0] n35704;
wire     [31:0] n35705;
wire     [31:0] n35706;
wire     [31:0] n35707;
wire     [31:0] n35708;
wire     [31:0] n35709;
wire     [31:0] n35710;
wire     [31:0] n35711;
wire     [31:0] n35712;
wire     [31:0] n35713;
wire     [31:0] n35714;
wire     [31:0] n35715;
wire     [31:0] n35716;
wire     [31:0] n35717;
wire     [31:0] n35718;
wire     [31:0] n35719;
wire     [31:0] n35720;
wire     [31:0] n35721;
wire     [31:0] n35722;
wire     [31:0] n35723;
wire     [31:0] n35724;
wire     [31:0] n35725;
wire     [31:0] n35726;
wire     [31:0] n35727;
wire     [31:0] n35728;
wire     [31:0] n35729;
wire     [31:0] n35730;
wire     [31:0] n35731;
wire     [31:0] n35732;
wire     [31:0] n35733;
wire     [31:0] n35734;
wire     [31:0] n35735;
wire     [31:0] n35736;
wire     [31:0] n35737;
wire     [31:0] n35738;
wire     [31:0] n35739;
wire     [31:0] n35740;
wire     [31:0] n35741;
wire     [31:0] n35742;
wire     [31:0] n35743;
wire     [31:0] n35744;
wire     [31:0] n35745;
wire     [31:0] n35746;
wire     [31:0] n35747;
wire     [31:0] n35748;
wire     [31:0] n35749;
wire     [31:0] n35750;
wire     [31:0] n35751;
wire     [31:0] n35752;
wire     [31:0] n35753;
wire     [31:0] n35754;
wire     [31:0] n35755;
wire     [31:0] n35756;
wire     [31:0] n35757;
wire     [31:0] n35758;
wire     [31:0] n35759;
wire     [31:0] n35760;
wire     [31:0] n35761;
wire     [31:0] n35762;
wire     [31:0] n35763;
wire     [31:0] n35764;
wire     [31:0] n35765;
wire     [31:0] n35766;
wire     [31:0] n35767;
wire     [31:0] n35768;
wire     [31:0] n35769;
wire     [31:0] n35770;
wire     [31:0] n35771;
wire     [31:0] n35772;
wire     [31:0] n35773;
wire     [31:0] n35774;
wire     [31:0] n35775;
wire     [31:0] n35776;
wire     [31:0] n35777;
wire     [31:0] n35778;
wire     [31:0] n35779;
wire     [31:0] n35780;
wire     [31:0] n35781;
wire     [31:0] n35782;
wire     [31:0] n35783;
wire     [31:0] n35784;
wire     [31:0] n35785;
wire     [31:0] n35786;
wire     [31:0] n35787;
wire     [31:0] n35788;
wire     [31:0] n35789;
wire     [31:0] n35790;
wire     [31:0] n35791;
wire     [31:0] n35792;
wire     [31:0] n35793;
wire     [31:0] n35794;
wire     [31:0] n35795;
wire     [31:0] n35796;
wire     [31:0] n35797;
wire     [31:0] n35798;
wire     [31:0] n35799;
wire     [31:0] n35800;
wire     [31:0] n35801;
wire     [31:0] n35802;
wire     [31:0] n35803;
wire     [31:0] n35804;
wire     [31:0] n35805;
wire     [31:0] n35806;
wire     [31:0] n35807;
wire     [31:0] n35808;
wire     [31:0] n35809;
wire     [31:0] n35810;
wire     [31:0] n35811;
wire     [31:0] n35812;
wire     [31:0] n35813;
wire     [31:0] n35814;
wire     [31:0] n35815;
wire     [31:0] n35816;
wire     [31:0] n35817;
wire     [31:0] n35818;
wire     [31:0] n35819;
wire     [31:0] n35820;
wire     [31:0] n35821;
wire     [31:0] n35822;
wire     [31:0] n35823;
wire     [31:0] n35824;
wire     [31:0] n35825;
wire     [31:0] n35826;
wire     [31:0] n35827;
wire     [31:0] n35828;
wire     [31:0] n35829;
wire     [31:0] n35830;
wire     [31:0] n35831;
wire     [31:0] n35832;
wire     [31:0] n35833;
wire     [31:0] n35834;
wire     [31:0] n35835;
wire     [31:0] n35836;
wire     [31:0] n35837;
wire     [31:0] n35838;
wire     [31:0] n35839;
wire     [31:0] n35840;
wire     [31:0] n35841;
wire     [31:0] n35842;
wire     [31:0] n35843;
wire     [31:0] n35844;
wire     [31:0] n35845;
wire     [31:0] n35846;
wire     [31:0] n35847;
wire     [31:0] n35848;
wire     [31:0] n35849;
wire     [31:0] n35850;
wire     [31:0] n35851;
wire     [31:0] n35852;
wire     [31:0] n35853;
wire     [31:0] n35854;
wire     [31:0] n35855;
wire     [31:0] n35856;
wire     [31:0] n35857;
wire     [31:0] n35858;
wire     [31:0] n35859;
wire     [31:0] n35860;
wire     [31:0] n35861;
wire     [31:0] n35862;
wire     [31:0] n35863;
wire     [31:0] n35864;
wire     [31:0] n35865;
wire     [31:0] n35866;
wire     [31:0] n35867;
wire     [31:0] n35868;
wire     [31:0] n35869;
wire     [31:0] n35870;
wire     [31:0] n35871;
wire     [31:0] n35872;
wire     [31:0] n35873;
wire     [31:0] n35874;
wire     [31:0] n35875;
wire     [31:0] n35876;
wire     [31:0] n35877;
wire     [31:0] n35878;
wire     [31:0] n35879;
wire     [31:0] n35880;
wire     [31:0] n35881;
wire     [31:0] n35882;
wire     [31:0] n35883;
wire     [31:0] n35884;
wire     [31:0] n35885;
wire     [31:0] n35886;
wire     [31:0] n35887;
wire     [31:0] n35888;
wire     [31:0] n35889;
wire     [31:0] n35890;
wire     [31:0] n35891;
wire     [31:0] n35892;
wire     [31:0] n35893;
wire     [31:0] n35894;
wire     [31:0] n35895;
wire     [31:0] n35896;
wire     [31:0] n35897;
wire     [31:0] n35898;
wire     [31:0] n35899;
wire     [31:0] n35900;
wire     [31:0] n35901;
wire     [31:0] n35902;
wire     [31:0] n35903;
wire     [31:0] n35904;
wire     [31:0] n35905;
wire     [31:0] n35906;
wire     [31:0] n35907;
wire     [31:0] n35908;
wire     [31:0] n35909;
wire     [31:0] n35910;
wire     [31:0] n35911;
wire     [31:0] n35912;
wire     [31:0] n35913;
wire     [31:0] n35914;
wire     [31:0] n35915;
wire     [31:0] n35916;
wire     [31:0] n35917;
wire     [31:0] n35918;
wire     [31:0] n35919;
wire     [31:0] n35920;
wire     [31:0] n35921;
wire     [31:0] n35922;
wire     [31:0] n35923;
wire     [31:0] n35924;
wire     [31:0] n35925;
wire     [31:0] n35926;
wire     [31:0] n35927;
wire     [31:0] n35928;
wire     [31:0] n35929;
wire     [31:0] n35930;
wire     [31:0] n35931;
wire     [31:0] n35932;
wire     [31:0] n35933;
wire     [31:0] n35934;
wire     [31:0] n35935;
wire     [31:0] n35936;
wire     [31:0] n35937;
wire     [31:0] n35938;
wire     [31:0] n35939;
wire     [31:0] n35940;
wire     [31:0] n35941;
wire     [31:0] n35942;
wire     [31:0] n35943;
wire     [31:0] n35944;
wire     [31:0] n35945;
wire     [31:0] n35946;
wire     [31:0] n35947;
wire     [31:0] n35948;
wire     [31:0] n35949;
wire     [31:0] n35950;
wire     [31:0] n35951;
wire     [31:0] n35952;
wire     [31:0] n35953;
wire     [31:0] n35954;
wire     [31:0] n35955;
wire     [31:0] n35956;
wire     [31:0] n35957;
wire     [31:0] n35958;
wire     [31:0] n35959;
wire     [31:0] n35960;
wire     [31:0] n35961;
wire     [31:0] n35962;
wire     [31:0] n35963;
wire     [31:0] n35964;
wire     [31:0] n35965;
wire     [31:0] n35966;
wire     [31:0] n35967;
wire     [31:0] n35968;
wire     [31:0] n35969;
wire     [31:0] n35970;
wire     [31:0] n35971;
wire     [31:0] n35972;
wire     [31:0] n35973;
wire     [31:0] n35974;
wire     [31:0] n35975;
wire     [31:0] n35976;
wire     [31:0] n35977;
wire     [31:0] n35978;
wire     [31:0] n35979;
wire     [31:0] n35980;
wire     [31:0] n35981;
wire     [31:0] n35982;
wire     [31:0] n35983;
wire     [31:0] n35984;
wire     [31:0] n35985;
wire     [31:0] n35986;
wire     [31:0] n35987;
wire     [31:0] n35988;
wire     [31:0] n35989;
wire     [31:0] n35990;
wire     [31:0] n35991;
wire     [31:0] n35992;
wire     [31:0] n35993;
wire     [31:0] n35994;
wire     [31:0] n35995;
wire     [31:0] n35996;
wire     [31:0] n35997;
wire     [31:0] n35998;
wire     [31:0] n35999;
wire     [31:0] n36000;
wire     [31:0] n36001;
wire     [31:0] n36002;
wire     [31:0] n36003;
wire     [31:0] n36004;
wire     [31:0] n36005;
wire     [31:0] n36006;
wire     [31:0] n36007;
wire     [31:0] n36008;
wire     [31:0] n36009;
wire     [31:0] n36010;
wire     [31:0] n36011;
wire     [31:0] n36012;
wire     [31:0] n36013;
wire     [31:0] n36014;
wire     [31:0] n36015;
wire     [31:0] n36016;
wire     [31:0] n36017;
wire     [31:0] n36018;
wire     [31:0] n36019;
wire     [31:0] n36020;
wire     [31:0] n36021;
wire     [31:0] n36022;
wire     [31:0] n36023;
wire     [31:0] n36024;
wire     [31:0] n36025;
wire     [31:0] n36026;
wire     [31:0] n36027;
wire     [31:0] n36028;
wire     [31:0] n36029;
wire     [31:0] n36030;
wire     [31:0] n36031;
wire     [31:0] n36032;
wire     [31:0] n36033;
wire     [31:0] n36034;
wire     [31:0] n36035;
wire     [31:0] n36036;
wire     [31:0] n36037;
wire     [31:0] n36038;
wire     [31:0] n36039;
wire     [31:0] n36040;
wire     [31:0] n36041;
wire     [31:0] n36042;
wire     [31:0] n36043;
wire     [31:0] n36044;
wire     [31:0] n36045;
wire     [31:0] n36046;
wire     [31:0] n36047;
wire     [31:0] n36048;
wire     [31:0] n36049;
wire     [31:0] n36050;
wire     [31:0] n36051;
wire     [31:0] n36052;
wire     [31:0] n36053;
wire     [31:0] n36054;
wire     [31:0] n36055;
wire     [31:0] n36056;
wire     [31:0] n36057;
wire     [31:0] n36058;
wire     [31:0] n36059;
wire     [31:0] n36060;
wire     [31:0] n36061;
wire     [31:0] n36062;
wire     [31:0] n36063;
wire     [31:0] n36064;
wire     [31:0] n36065;
wire     [31:0] n36066;
wire     [31:0] n36067;
wire     [31:0] n36068;
wire     [31:0] n36069;
wire     [31:0] n36070;
wire     [31:0] n36071;
wire     [31:0] n36072;
wire     [31:0] n36073;
wire     [31:0] n36074;
wire     [31:0] n36075;
wire     [31:0] n36076;
wire     [31:0] n36077;
wire     [31:0] n36078;
wire     [31:0] n36079;
wire     [31:0] n36080;
wire     [31:0] n36081;
wire     [31:0] n36082;
wire     [31:0] n36083;
wire     [31:0] n36084;
wire     [31:0] n36085;
wire     [31:0] n36086;
wire     [31:0] n36087;
wire     [31:0] n36088;
wire     [31:0] n36089;
wire     [31:0] n36090;
wire     [31:0] n36091;
wire     [31:0] n36092;
wire     [31:0] n36093;
wire     [31:0] n36094;
wire     [31:0] n36095;
wire     [31:0] n36096;
wire     [31:0] n36097;
wire     [31:0] n36098;
wire     [31:0] n36099;
wire     [31:0] n36100;
wire     [31:0] n36101;
wire     [31:0] n36102;
wire     [31:0] n36103;
wire     [31:0] n36104;
wire     [31:0] n36105;
wire     [31:0] n36106;
wire     [31:0] n36107;
wire     [31:0] n36108;
wire     [31:0] n36109;
wire     [31:0] n36110;
wire     [31:0] n36111;
wire     [31:0] n36112;
wire     [31:0] n36113;
wire     [31:0] n36114;
wire     [31:0] n36115;
wire     [31:0] n36116;
wire     [31:0] n36117;
wire     [31:0] n36118;
wire     [31:0] n36119;
wire     [31:0] n36120;
wire     [31:0] n36121;
wire     [31:0] n36122;
wire     [31:0] n36123;
wire     [31:0] n36124;
wire     [31:0] n36125;
wire     [31:0] n36126;
wire     [31:0] n36127;
wire     [31:0] n36128;
wire     [31:0] n36129;
wire     [31:0] n36130;
wire     [31:0] n36131;
wire     [31:0] n36132;
wire     [31:0] n36133;
wire     [31:0] n36134;
wire     [31:0] n36135;
wire     [31:0] n36136;
wire     [31:0] n36137;
wire     [31:0] n36138;
wire     [31:0] n36139;
wire     [31:0] n36140;
wire     [31:0] n36141;
wire     [31:0] n36142;
wire     [31:0] n36143;
wire     [31:0] n36144;
wire     [31:0] n36145;
wire     [31:0] n36146;
wire     [31:0] n36147;
wire     [31:0] n36148;
wire     [31:0] n36149;
wire     [31:0] n36150;
wire     [31:0] n36151;
wire     [31:0] n36152;
wire     [31:0] n36153;
wire     [31:0] n36154;
wire     [31:0] n36155;
wire     [31:0] n36156;
wire     [31:0] n36157;
wire     [31:0] n36158;
wire     [31:0] n36159;
wire     [31:0] n36160;
wire     [31:0] n36161;
wire     [31:0] n36162;
wire     [31:0] n36163;
wire     [31:0] n36164;
wire     [31:0] n36165;
wire     [31:0] n36166;
wire     [31:0] n36167;
wire     [31:0] n36168;
wire     [31:0] n36169;
wire     [31:0] n36170;
wire     [31:0] n36171;
wire     [31:0] n36172;
wire     [31:0] n36173;
wire     [31:0] n36174;
wire     [31:0] n36175;
wire     [31:0] n36176;
wire     [31:0] n36177;
wire     [31:0] n36178;
wire     [31:0] n36179;
wire     [31:0] n36180;
wire     [31:0] n36181;
wire     [31:0] n36182;
wire     [31:0] n36183;
wire     [31:0] n36184;
wire     [31:0] n36185;
wire     [31:0] n36186;
wire     [31:0] n36187;
wire     [31:0] n36188;
wire     [31:0] n36189;
wire     [31:0] n36190;
wire     [31:0] n36191;
wire     [31:0] n36192;
wire     [31:0] n36193;
wire     [31:0] n36194;
wire     [31:0] n36195;
wire     [31:0] n36196;
wire     [31:0] n36197;
wire     [31:0] n36198;
wire     [31:0] n36199;
wire     [31:0] n36200;
wire     [31:0] n36201;
wire     [31:0] n36202;
wire     [31:0] n36203;
wire     [31:0] n36204;
wire     [31:0] n36205;
wire     [31:0] n36206;
wire     [31:0] n36207;
wire     [31:0] n36208;
wire     [31:0] n36209;
wire     [31:0] n36210;
wire     [31:0] n36211;
wire     [31:0] n36212;
wire     [31:0] n36213;
wire     [31:0] n36214;
wire     [31:0] n36215;
wire     [31:0] n36216;
wire     [31:0] n36217;
wire     [31:0] n36218;
wire     [31:0] n36219;
wire     [31:0] n36220;
wire     [31:0] n36221;
wire     [31:0] n36222;
wire     [31:0] n36223;
wire     [31:0] n36224;
wire     [31:0] n36225;
wire     [31:0] n36226;
wire     [31:0] n36227;
wire     [31:0] n36228;
wire     [31:0] n36229;
wire     [31:0] n36230;
wire     [31:0] n36231;
wire     [31:0] n36232;
wire     [31:0] n36233;
wire     [31:0] n36234;
wire     [31:0] n36235;
wire     [31:0] n36236;
wire     [31:0] n36237;
wire     [31:0] n36238;
wire     [31:0] n36239;
wire     [31:0] n36240;
wire     [31:0] n36241;
wire     [31:0] n36242;
wire     [31:0] n36243;
wire     [31:0] n36244;
wire     [31:0] n36245;
wire     [31:0] n36246;
wire     [31:0] n36247;
wire     [31:0] n36248;
wire     [31:0] n36249;
wire     [31:0] n36250;
wire     [31:0] n36251;
wire     [31:0] n36252;
wire     [31:0] n36253;
wire     [31:0] n36254;
wire     [31:0] n36255;
wire     [31:0] n36256;
wire     [31:0] n36257;
wire     [31:0] n36258;
wire     [31:0] n36259;
wire     [31:0] n36260;
wire     [31:0] n36261;
wire     [31:0] n36262;
wire     [31:0] n36263;
wire     [31:0] n36264;
wire     [31:0] n36265;
wire     [31:0] n36266;
wire     [31:0] n36267;
wire     [31:0] n36268;
wire     [31:0] n36269;
wire     [31:0] n36270;
wire     [31:0] n36271;
wire     [31:0] n36272;
wire     [31:0] n36273;
wire     [31:0] n36274;
wire     [31:0] n36275;
wire     [31:0] n36276;
wire     [31:0] n36277;
wire     [31:0] n36278;
wire     [31:0] n36279;
wire     [31:0] n36280;
wire     [31:0] n36281;
wire     [31:0] n36282;
wire     [31:0] n36283;
wire     [31:0] n36284;
wire     [31:0] n36285;
wire     [31:0] n36286;
wire     [31:0] n36287;
wire     [31:0] n36288;
wire     [31:0] n36289;
wire     [31:0] n36290;
wire     [31:0] n36291;
wire     [31:0] n36292;
wire     [31:0] n36293;
wire     [31:0] n36294;
wire     [31:0] n36295;
wire     [31:0] n36296;
wire     [31:0] n36297;
wire     [31:0] n36298;
wire     [31:0] n36299;
wire     [31:0] n36300;
wire     [31:0] n36301;
wire     [31:0] n36302;
wire     [31:0] n36303;
wire     [31:0] n36304;
wire     [31:0] n36305;
wire     [31:0] n36306;
wire     [31:0] n36307;
wire     [31:0] n36308;
wire     [31:0] n36309;
wire     [31:0] n36310;
wire     [31:0] n36311;
wire     [31:0] n36312;
wire     [31:0] n36313;
wire     [31:0] n36314;
wire     [31:0] n36315;
wire     [31:0] n36316;
wire     [31:0] n36317;
wire     [31:0] n36318;
wire     [31:0] n36319;
wire     [31:0] n36320;
wire     [31:0] n36321;
wire     [31:0] n36322;
wire     [31:0] n36323;
wire     [31:0] n36324;
wire     [31:0] n36325;
wire     [31:0] n36326;
wire     [31:0] n36327;
wire     [31:0] n36328;
wire     [31:0] n36329;
wire     [31:0] n36330;
wire     [31:0] n36331;
wire     [31:0] n36332;
wire     [31:0] n36333;
wire     [31:0] n36334;
wire     [31:0] n36335;
wire     [31:0] n36336;
wire     [31:0] n36337;
wire     [31:0] n36338;
wire     [31:0] n36339;
wire     [31:0] n36340;
wire     [31:0] n36341;
wire     [31:0] n36342;
wire     [31:0] n36343;
wire     [31:0] n36344;
wire     [31:0] n36345;
wire     [31:0] n36346;
wire     [31:0] n36347;
wire     [31:0] n36348;
wire     [31:0] n36349;
wire     [31:0] n36350;
wire     [31:0] n36351;
wire     [31:0] n36352;
wire     [31:0] n36353;
wire     [31:0] n36354;
wire     [31:0] n36355;
wire     [31:0] n36356;
wire     [31:0] n36357;
wire     [31:0] n36358;
wire     [31:0] n36359;
wire     [31:0] n36360;
wire     [31:0] n36361;
wire     [31:0] n36362;
wire     [31:0] n36363;
wire     [31:0] n36364;
wire     [31:0] n36365;
wire     [31:0] n36366;
wire     [31:0] n36367;
wire     [31:0] n36368;
wire     [31:0] n36369;
wire     [31:0] n36370;
wire     [31:0] n36371;
wire     [31:0] n36372;
wire     [31:0] n36373;
wire     [31:0] n36374;
wire     [31:0] n36375;
wire     [31:0] n36376;
wire     [31:0] n36377;
wire     [31:0] n36378;
wire     [31:0] n36379;
wire     [31:0] n36380;
wire     [31:0] n36381;
wire     [31:0] n36382;
wire     [31:0] n36383;
wire     [31:0] n36384;
wire     [31:0] n36385;
wire     [31:0] n36386;
wire     [31:0] n36387;
wire     [31:0] n36388;
wire     [31:0] n36389;
wire     [31:0] n36390;
wire     [31:0] n36391;
wire     [31:0] n36392;
wire     [31:0] n36393;
wire     [31:0] n36394;
wire     [31:0] n36395;
wire     [31:0] n36396;
wire     [31:0] n36397;
wire     [31:0] n36398;
wire     [31:0] n36399;
wire     [31:0] n36400;
wire     [31:0] n36401;
wire     [31:0] n36402;
wire     [31:0] n36403;
wire     [31:0] n36404;
wire     [31:0] n36405;
wire     [31:0] n36406;
wire     [31:0] n36407;
wire     [31:0] n36408;
wire     [31:0] n36409;
wire     [31:0] n36410;
wire     [31:0] n36411;
wire     [31:0] n36412;
wire     [31:0] n36413;
wire     [31:0] n36414;
wire     [31:0] n36415;
wire     [31:0] n36416;
wire     [31:0] n36417;
wire     [31:0] n36418;
wire     [31:0] n36419;
wire     [31:0] n36420;
wire     [31:0] n36421;
wire     [31:0] n36422;
wire     [31:0] n36423;
wire     [31:0] n36424;
wire     [31:0] n36425;
wire     [31:0] n36426;
wire     [31:0] n36427;
wire     [31:0] n36428;
wire     [31:0] n36429;
wire     [31:0] n36430;
wire     [31:0] n36431;
wire     [31:0] n36432;
wire     [31:0] n36433;
wire     [31:0] n36434;
wire     [31:0] n36435;
wire     [31:0] n36436;
wire     [31:0] n36437;
wire     [31:0] n36438;
wire     [31:0] n36439;
wire     [31:0] n36440;
wire     [31:0] n36441;
wire     [31:0] n36442;
wire     [31:0] n36443;
wire     [31:0] n36444;
wire     [31:0] n36445;
wire     [31:0] n36446;
wire     [31:0] n36447;
wire     [31:0] n36448;
wire     [31:0] n36449;
wire     [31:0] n36450;
wire     [31:0] n36451;
wire     [31:0] n36452;
wire     [31:0] n36453;
wire     [31:0] n36454;
wire     [31:0] n36455;
wire     [31:0] n36456;
wire     [31:0] n36457;
wire     [31:0] n36458;
wire     [31:0] n36459;
wire     [31:0] n36460;
wire     [31:0] n36461;
wire     [31:0] n36462;
wire     [31:0] n36463;
wire     [31:0] n36464;
wire     [31:0] n36465;
wire     [31:0] n36466;
wire     [31:0] n36467;
wire     [31:0] n36468;
wire     [31:0] n36469;
wire     [31:0] n36470;
wire     [31:0] n36471;
wire     [31:0] n36472;
wire     [31:0] n36473;
wire     [31:0] n36474;
wire     [31:0] n36475;
wire     [31:0] n36476;
wire     [31:0] n36477;
wire     [31:0] n36478;
wire     [31:0] n36479;
wire     [31:0] n36480;
wire     [31:0] n36481;
wire     [31:0] n36482;
wire     [31:0] n36483;
wire     [31:0] n36484;
wire     [31:0] n36485;
wire     [31:0] n36486;
wire     [31:0] n36487;
wire     [31:0] n36488;
wire     [31:0] n36489;
wire     [31:0] n36490;
wire     [31:0] n36491;
wire     [31:0] n36492;
wire     [31:0] n36493;
wire     [31:0] n36494;
wire     [31:0] n36495;
wire     [31:0] n36496;
wire     [31:0] n36497;
wire     [31:0] n36498;
wire     [31:0] n36499;
wire     [31:0] n36500;
wire     [31:0] n36501;
wire     [31:0] n36502;
wire     [31:0] n36503;
wire     [31:0] n36504;
wire     [31:0] n36505;
wire     [31:0] n36506;
wire     [31:0] n36507;
wire     [31:0] n36508;
wire     [31:0] n36509;
wire     [31:0] n36510;
wire     [31:0] n36511;
wire     [31:0] n36512;
wire     [31:0] n36513;
wire     [31:0] n36514;
wire     [31:0] n36515;
wire     [31:0] n36516;
wire     [31:0] n36517;
wire     [31:0] n36518;
wire     [31:0] n36519;
wire     [31:0] n36520;
wire     [31:0] n36521;
wire     [31:0] n36522;
wire     [31:0] n36523;
wire     [31:0] n36524;
wire     [31:0] n36525;
wire     [31:0] n36526;
wire     [31:0] n36527;
wire     [31:0] n36528;
wire     [31:0] n36529;
wire     [31:0] n36530;
wire     [31:0] n36531;
wire     [31:0] n36532;
wire     [31:0] n36533;
wire     [31:0] n36534;
wire     [31:0] n36535;
wire     [31:0] n36536;
wire     [31:0] n36537;
wire     [31:0] n36538;
wire     [31:0] n36539;
wire     [31:0] n36540;
wire     [31:0] n36541;
wire     [31:0] n36542;
wire     [31:0] n36543;
wire     [31:0] n36544;
wire     [31:0] n36545;
wire     [31:0] n36546;
wire     [31:0] n36547;
wire     [31:0] n36548;
wire     [31:0] n36549;
wire     [31:0] n36550;
wire     [31:0] n36551;
wire     [31:0] n36552;
wire     [31:0] n36553;
wire     [31:0] n36554;
wire     [31:0] n36555;
wire     [31:0] n36556;
wire     [31:0] n36557;
wire     [31:0] n36558;
wire     [31:0] n36559;
wire     [31:0] n36560;
wire     [31:0] n36561;
wire     [31:0] n36562;
wire     [31:0] n36563;
wire     [31:0] n36564;
wire     [31:0] n36565;
wire     [31:0] n36566;
wire     [31:0] n36567;
wire     [31:0] n36568;
wire     [31:0] n36569;
wire     [31:0] n36570;
wire     [31:0] n36571;
wire     [31:0] n36572;
wire     [31:0] n36573;
wire     [31:0] n36574;
wire     [31:0] n36575;
wire     [31:0] n36576;
wire     [31:0] n36577;
wire     [31:0] n36578;
wire     [31:0] n36579;
wire     [31:0] n36580;
wire     [31:0] n36581;
wire     [31:0] n36582;
wire     [31:0] n36583;
wire     [31:0] n36584;
wire     [31:0] n36585;
wire     [31:0] n36586;
wire     [31:0] n36587;
wire     [31:0] n36588;
wire     [31:0] n36589;
wire     [31:0] n36590;
wire     [31:0] n36591;
wire     [31:0] n36592;
wire     [31:0] n36593;
wire     [31:0] n36594;
wire     [31:0] n36595;
wire     [31:0] n36596;
wire     [31:0] n36597;
wire     [31:0] n36598;
wire     [31:0] n36599;
wire     [31:0] n36600;
wire     [31:0] n36601;
wire     [31:0] n36602;
wire     [31:0] n36603;
wire     [31:0] n36604;
wire     [31:0] n36605;
wire     [31:0] n36606;
wire     [31:0] n36607;
wire     [31:0] n36608;
wire     [31:0] n36609;
wire     [31:0] n36610;
wire     [31:0] n36611;
wire     [31:0] n36612;
wire     [31:0] n36613;
wire     [31:0] n36614;
wire     [31:0] n36615;
wire     [31:0] n36616;
wire     [31:0] n36617;
wire     [31:0] n36618;
wire     [31:0] n36619;
wire     [31:0] n36620;
wire     [31:0] n36621;
wire     [31:0] n36622;
wire     [31:0] n36623;
wire     [31:0] n36624;
wire     [31:0] n36625;
wire     [31:0] n36626;
wire     [31:0] n36627;
wire     [31:0] n36628;
wire     [31:0] n36629;
wire     [31:0] n36630;
wire     [31:0] n36631;
wire     [31:0] n36632;
wire     [31:0] n36633;
wire     [31:0] n36634;
wire     [31:0] n36635;
wire     [31:0] n36636;
wire     [31:0] n36637;
wire     [31:0] n36638;
wire     [31:0] n36639;
wire     [31:0] n36640;
wire     [31:0] n36641;
wire     [31:0] n36642;
wire     [31:0] n36643;
wire     [31:0] n36644;
wire     [31:0] n36645;
wire     [31:0] n36646;
wire     [31:0] n36647;
wire     [31:0] n36648;
wire     [31:0] n36649;
wire     [31:0] n36650;
wire     [31:0] n36651;
wire     [31:0] n36652;
wire     [31:0] n36653;
wire     [31:0] n36654;
wire     [31:0] n36655;
wire     [31:0] n36656;
wire     [31:0] n36657;
wire     [31:0] n36658;
wire     [31:0] n36659;
wire     [31:0] n36660;
wire     [31:0] n36661;
wire     [31:0] n36662;
wire     [31:0] n36663;
wire     [31:0] n36664;
wire     [31:0] n36665;
wire     [31:0] n36666;
wire     [31:0] n36667;
wire     [31:0] n36668;
wire     [31:0] n36669;
wire     [31:0] n36670;
wire     [31:0] n36671;
wire     [31:0] n36672;
wire     [31:0] n36673;
wire     [31:0] n36674;
wire     [31:0] n36675;
wire     [31:0] n36676;
wire     [31:0] n36677;
wire     [31:0] n36678;
wire     [31:0] n36679;
wire     [31:0] n36680;
wire     [31:0] n36681;
wire     [31:0] n36682;
wire     [31:0] n36683;
wire     [31:0] n36684;
wire     [31:0] n36685;
wire     [31:0] n36686;
wire     [31:0] n36687;
wire     [31:0] n36688;
wire     [31:0] n36689;
wire     [31:0] n36690;
wire     [31:0] n36691;
wire     [31:0] n36692;
wire     [31:0] n36693;
wire     [31:0] n36694;
wire     [31:0] n36695;
wire     [31:0] n36696;
wire     [31:0] n36697;
wire     [31:0] n36698;
wire     [31:0] n36699;
wire     [31:0] n36700;
wire     [31:0] n36701;
wire     [31:0] n36702;
wire     [31:0] n36703;
wire     [31:0] n36704;
wire     [31:0] n36705;
wire     [31:0] n36706;
wire     [31:0] n36707;
wire     [31:0] n36708;
wire     [31:0] n36709;
wire     [31:0] n36710;
wire     [31:0] n36711;
wire     [31:0] n36712;
wire     [31:0] n36713;
wire     [31:0] n36714;
wire     [31:0] n36715;
wire     [31:0] n36716;
wire     [31:0] n36717;
wire     [31:0] n36718;
wire     [31:0] n36719;
wire     [31:0] n36720;
wire     [31:0] n36721;
wire     [31:0] n36722;
wire     [31:0] n36723;
wire     [31:0] n36724;
wire     [31:0] n36725;
wire     [31:0] n36726;
wire     [31:0] n36727;
wire     [31:0] n36728;
wire     [31:0] n36729;
wire     [31:0] n36730;
wire     [31:0] n36731;
wire     [31:0] n36732;
wire     [31:0] n36733;
wire     [31:0] n36734;
wire     [31:0] n36735;
wire     [31:0] n36736;
wire     [31:0] n36737;
wire     [31:0] n36738;
wire     [31:0] n36739;
wire     [31:0] n36740;
wire     [31:0] n36741;
wire     [31:0] n36742;
wire     [31:0] n36743;
wire     [31:0] n36744;
wire     [31:0] n36745;
wire     [31:0] n36746;
wire     [31:0] n36747;
wire     [31:0] n36748;
wire     [31:0] n36749;
wire     [31:0] n36750;
wire     [31:0] n36751;
wire     [31:0] n36752;
wire     [31:0] n36753;
wire     [31:0] n36754;
wire     [31:0] n36755;
wire     [31:0] n36756;
wire     [31:0] n36757;
wire     [31:0] n36758;
wire     [31:0] n36759;
wire     [31:0] n36760;
wire     [31:0] n36761;
wire     [31:0] n36762;
wire     [31:0] n36763;
wire     [31:0] n36764;
wire     [31:0] n36765;
wire     [31:0] n36766;
wire     [31:0] n36767;
wire     [31:0] n36768;
wire     [31:0] n36769;
wire     [31:0] n36770;
wire     [31:0] n36771;
wire     [31:0] n36772;
wire     [31:0] n36773;
wire     [31:0] n36774;
wire     [31:0] n36775;
wire     [31:0] n36776;
wire     [31:0] n36777;
wire     [31:0] n36778;
wire     [31:0] n36779;
wire     [31:0] n36780;
wire     [31:0] n36781;
wire     [31:0] n36782;
wire     [31:0] n36783;
wire     [31:0] n36784;
wire     [31:0] n36785;
wire     [31:0] n36786;
wire     [31:0] n36787;
wire     [31:0] n36788;
wire     [31:0] n36789;
wire     [31:0] n36790;
wire     [31:0] n36791;
wire     [31:0] n36792;
wire     [31:0] n36793;
wire     [31:0] n36794;
wire     [31:0] n36795;
wire     [31:0] n36796;
wire     [31:0] n36797;
wire     [31:0] n36798;
wire     [31:0] n36799;
wire     [31:0] n36800;
wire     [31:0] n36801;
wire     [31:0] n36802;
wire     [31:0] n36803;
wire     [31:0] n36804;
wire     [31:0] n36805;
wire     [31:0] n36806;
wire     [31:0] n36807;
wire     [31:0] n36808;
wire     [31:0] n36809;
wire     [31:0] n36810;
wire     [31:0] n36811;
wire     [31:0] n36812;
wire     [31:0] n36813;
wire     [31:0] n36814;
wire     [31:0] n36815;
wire     [31:0] n36816;
wire     [31:0] n36817;
wire     [31:0] n36818;
wire     [31:0] n36819;
wire     [31:0] n36820;
wire     [31:0] n36821;
wire     [31:0] n36822;
wire     [31:0] n36823;
wire     [31:0] n36824;
wire     [31:0] n36825;
wire     [31:0] n36826;
wire     [31:0] n36827;
wire     [31:0] n36828;
wire     [31:0] n36829;
wire     [31:0] n36830;
wire     [31:0] n36831;
wire     [31:0] n36832;
wire     [31:0] n36833;
wire     [31:0] n36834;
wire     [31:0] n36835;
wire     [31:0] n36836;
wire     [31:0] n36837;
wire     [31:0] n36838;
wire     [31:0] n36839;
wire     [31:0] n36840;
wire     [31:0] n36841;
wire     [31:0] n36842;
wire     [31:0] n36843;
wire     [31:0] n36844;
wire     [31:0] n36845;
wire     [31:0] n36846;
wire     [31:0] n36847;
wire     [31:0] n36848;
wire     [31:0] n36849;
wire     [31:0] n36850;
wire     [31:0] n36851;
wire     [31:0] n36852;
wire     [31:0] n36853;
wire     [31:0] n36854;
wire     [31:0] n36855;
wire     [31:0] n36856;
wire     [31:0] n36857;
wire     [31:0] n36858;
wire     [31:0] n36859;
wire     [31:0] n36860;
wire     [31:0] n36861;
wire     [31:0] n36862;
wire     [31:0] n36863;
wire     [31:0] n36864;
wire     [31:0] n36865;
wire     [31:0] n36866;
wire     [31:0] n36867;
wire     [31:0] n36868;
wire     [31:0] n36869;
wire     [31:0] n36870;
wire     [31:0] n36871;
wire     [31:0] n36872;
wire     [31:0] n36873;
wire     [31:0] n36874;
wire     [31:0] n36875;
wire     [31:0] n36876;
wire     [31:0] n36877;
wire     [31:0] n36878;
wire     [31:0] n36879;
wire     [31:0] n36880;
wire     [31:0] n36881;
wire     [31:0] n36882;
wire     [31:0] n36883;
wire     [31:0] n36884;
wire     [31:0] n36885;
wire     [31:0] n36886;
wire     [31:0] n36887;
wire     [31:0] n36888;
wire     [31:0] n36889;
wire     [31:0] n36890;
wire     [31:0] n36891;
wire     [31:0] n36892;
wire     [31:0] n36893;
wire     [31:0] n36894;
wire     [31:0] n36895;
wire     [31:0] n36896;
wire     [31:0] n36897;
wire     [31:0] n36898;
wire     [31:0] n36899;
wire     [31:0] n36900;
wire     [31:0] n36901;
wire     [31:0] n36902;
wire     [31:0] n36903;
wire     [31:0] n36904;
wire     [31:0] n36905;
wire     [31:0] n36906;
wire     [31:0] n36907;
wire     [31:0] n36908;
wire     [31:0] n36909;
wire     [31:0] n36910;
wire     [31:0] n36911;
wire     [31:0] n36912;
wire     [31:0] n36913;
wire     [31:0] n36914;
wire     [31:0] n36915;
wire     [31:0] n36916;
wire     [31:0] n36917;
wire     [31:0] n36918;
wire     [31:0] n36919;
wire     [31:0] n36920;
wire     [31:0] n36921;
wire     [31:0] n36922;
wire     [31:0] n36923;
wire     [31:0] n36924;
wire     [31:0] n36925;
wire     [31:0] n36926;
wire     [31:0] n36927;
wire     [31:0] n36928;
wire     [31:0] n36929;
wire     [31:0] n36930;
wire     [31:0] n36931;
wire     [31:0] n36932;
wire     [31:0] n36933;
wire     [31:0] n36934;
wire     [31:0] n36935;
wire     [31:0] n36936;
wire     [31:0] n36937;
wire     [31:0] n36938;
wire     [31:0] n36939;
wire     [31:0] n36940;
wire     [31:0] n36941;
wire     [31:0] n36942;
wire     [31:0] n36943;
wire     [31:0] n36944;
wire     [31:0] n36945;
wire     [31:0] n36946;
wire     [31:0] n36947;
wire     [31:0] n36948;
wire     [31:0] n36949;
wire     [31:0] n36950;
wire     [31:0] n36951;
wire     [31:0] n36952;
wire     [31:0] n36953;
wire     [31:0] n36954;
wire     [31:0] n36955;
wire     [31:0] n36956;
wire     [31:0] n36957;
wire     [31:0] n36958;
wire     [31:0] n36959;
wire     [31:0] n36960;
wire     [31:0] n36961;
wire     [31:0] n36962;
wire     [31:0] n36963;
wire     [31:0] n36964;
wire     [31:0] n36965;
wire     [31:0] n36966;
wire     [31:0] n36967;
wire     [31:0] n36968;
wire     [31:0] n36969;
wire     [31:0] n36970;
wire     [31:0] n36971;
wire     [31:0] n36972;
wire     [31:0] n36973;
wire     [31:0] n36974;
wire     [31:0] n36975;
wire     [31:0] n36976;
wire     [31:0] n36977;
wire     [31:0] n36978;
wire     [31:0] n36979;
wire     [31:0] n36980;
wire     [31:0] n36981;
wire     [31:0] n36982;
wire     [31:0] n36983;
wire     [31:0] n36984;
wire     [31:0] n36985;
wire     [31:0] n36986;
wire     [31:0] n36987;
wire     [31:0] n36988;
wire     [31:0] n36989;
wire     [31:0] n36990;
wire     [31:0] n36991;
wire     [31:0] n36992;
wire     [31:0] n36993;
wire     [31:0] n36994;
wire     [31:0] n36995;
wire     [31:0] n36996;
wire     [31:0] n36997;
wire     [31:0] n36998;
wire     [31:0] n36999;
wire     [31:0] n37000;
wire     [31:0] n37001;
wire     [31:0] n37002;
wire     [31:0] n37003;
wire     [31:0] n37004;
wire     [31:0] n37005;
wire     [31:0] n37006;
wire     [31:0] n37007;
wire     [31:0] n37008;
wire     [31:0] n37009;
wire     [31:0] n37010;
wire     [31:0] n37011;
wire     [31:0] n37012;
wire     [31:0] n37013;
wire     [31:0] n37014;
wire     [31:0] n37015;
wire     [31:0] n37016;
wire     [31:0] n37017;
wire     [31:0] n37018;
wire     [31:0] n37019;
wire     [31:0] n37020;
wire     [31:0] n37021;
wire     [31:0] n37022;
wire     [31:0] n37023;
wire     [31:0] n37024;
wire     [31:0] n37025;
wire     [31:0] n37026;
wire     [31:0] n37027;
wire     [31:0] n37028;
wire     [31:0] n37029;
wire     [31:0] n37030;
wire     [31:0] n37031;
wire     [31:0] n37032;
wire     [31:0] n37033;
wire     [31:0] n37034;
wire     [31:0] n37035;
wire     [31:0] n37036;
wire     [31:0] n37037;
wire     [31:0] n37038;
wire     [31:0] n37039;
wire     [31:0] n37040;
wire     [31:0] n37041;
wire     [31:0] n37042;
wire     [31:0] n37043;
wire     [31:0] n37044;
wire     [31:0] n37045;
wire     [31:0] n37046;
wire     [31:0] n37047;
wire     [31:0] n37048;
wire     [31:0] n37049;
wire     [31:0] n37050;
wire     [31:0] n37051;
wire     [31:0] n37052;
wire     [31:0] n37053;
wire     [31:0] n37054;
wire     [31:0] n37055;
wire     [31:0] n37056;
wire     [31:0] n37057;
wire     [31:0] n37058;
wire     [31:0] n37059;
wire     [31:0] n37060;
wire     [31:0] n37061;
wire     [31:0] n37062;
wire     [31:0] n37063;
wire     [31:0] n37064;
wire     [31:0] n37065;
wire     [31:0] n37066;
wire     [31:0] n37067;
wire     [31:0] n37068;
wire     [31:0] n37069;
wire     [31:0] n37070;
wire     [31:0] n37071;
wire     [31:0] n37072;
wire     [31:0] n37073;
wire     [31:0] n37074;
wire     [31:0] n37075;
wire     [31:0] n37076;
wire     [31:0] n37077;
wire     [31:0] n37078;
wire     [31:0] n37079;
wire     [31:0] n37080;
wire     [31:0] n37081;
wire     [31:0] n37082;
wire     [31:0] n37083;
wire     [31:0] n37084;
wire     [31:0] n37085;
wire     [31:0] n37086;
wire     [31:0] n37087;
wire     [31:0] n37088;
wire     [31:0] n37089;
wire     [31:0] n37090;
wire     [31:0] n37091;
wire     [31:0] n37092;
wire     [31:0] n37093;
wire     [31:0] n37094;
wire     [31:0] n37095;
wire     [31:0] n37096;
wire     [31:0] n37097;
wire     [31:0] n37098;
wire     [31:0] n37099;
wire     [31:0] n37100;
wire     [31:0] n37101;
wire     [31:0] n37102;
wire     [31:0] n37103;
wire     [31:0] n37104;
wire     [31:0] n37105;
wire     [31:0] n37106;
wire     [31:0] n37107;
wire     [31:0] n37108;
wire     [31:0] n37109;
wire     [31:0] n37110;
wire     [31:0] n37111;
wire     [31:0] n37112;
wire     [31:0] n37113;
wire     [31:0] n37114;
wire     [31:0] n37115;
wire     [31:0] n37116;
wire     [31:0] n37117;
wire     [31:0] n37118;
wire     [31:0] n37119;
wire     [31:0] n37120;
wire     [31:0] n37121;
wire     [31:0] n37122;
wire     [31:0] n37123;
wire     [31:0] n37124;
wire     [31:0] n37125;
wire     [31:0] n37126;
wire     [31:0] n37127;
wire     [31:0] n37128;
wire     [31:0] n37129;
wire     [31:0] n37130;
wire     [31:0] n37131;
wire     [31:0] n37132;
wire     [31:0] n37133;
wire     [31:0] n37134;
wire     [31:0] n37135;
wire     [31:0] n37136;
wire     [31:0] n37137;
wire     [31:0] n37138;
wire     [31:0] n37139;
wire     [31:0] n37140;
wire     [31:0] n37141;
wire     [31:0] n37142;
wire     [31:0] n37143;
wire     [31:0] n37144;
wire     [31:0] n37145;
wire     [31:0] n37146;
wire     [31:0] n37147;
wire     [31:0] n37148;
wire     [31:0] n37149;
wire     [31:0] n37150;
wire     [31:0] n37151;
wire     [31:0] n37152;
wire     [31:0] n37153;
wire     [31:0] n37154;
wire     [31:0] n37155;
wire     [31:0] n37156;
wire     [31:0] n37157;
wire     [31:0] n37158;
wire     [31:0] n37159;
wire     [31:0] n37160;
wire     [31:0] n37161;
wire     [31:0] n37162;
wire     [31:0] n37163;
wire     [31:0] n37164;
wire     [31:0] n37165;
wire     [31:0] n37166;
wire     [31:0] n37167;
wire     [31:0] n37168;
wire     [31:0] n37169;
wire     [31:0] n37170;
wire     [31:0] n37171;
wire     [31:0] n37172;
wire     [31:0] n37173;
wire     [31:0] n37174;
wire     [31:0] n37175;
wire     [31:0] n37176;
wire     [31:0] n37177;
wire     [31:0] n37178;
wire     [31:0] n37179;
wire     [31:0] n37180;
wire     [31:0] n37181;
wire     [31:0] n37182;
wire     [31:0] n37183;
wire     [31:0] n37184;
wire     [31:0] n37185;
wire     [31:0] n37186;
wire     [31:0] n37187;
wire     [31:0] n37188;
wire     [31:0] n37189;
wire     [31:0] n37190;
wire     [31:0] n37191;
wire     [31:0] n37192;
wire     [31:0] n37193;
wire     [31:0] n37194;
wire     [31:0] n37195;
wire     [31:0] n37196;
wire     [31:0] n37197;
wire     [31:0] n37198;
wire     [31:0] n37199;
wire     [31:0] n37200;
wire     [31:0] n37201;
wire     [31:0] n37202;
wire     [31:0] n37203;
wire     [31:0] n37204;
wire     [31:0] n37205;
wire     [31:0] n37206;
wire     [31:0] n37207;
wire     [31:0] n37208;
wire     [31:0] n37209;
wire     [31:0] n37210;
wire     [31:0] n37211;
wire     [31:0] n37212;
wire     [31:0] n37213;
wire     [31:0] n37214;
wire     [31:0] n37215;
wire     [31:0] n37216;
wire     [31:0] n37217;
wire     [31:0] n37218;
wire     [31:0] n37219;
wire     [31:0] n37220;
wire     [31:0] n37221;
wire     [31:0] n37222;
wire     [31:0] n37223;
wire     [31:0] n37224;
wire     [31:0] n37225;
wire     [31:0] n37226;
wire     [31:0] n37227;
wire     [31:0] n37228;
wire     [31:0] n37229;
wire     [31:0] n37230;
wire     [31:0] n37231;
wire     [31:0] n37232;
wire     [31:0] n37233;
wire     [31:0] n37234;
wire     [31:0] n37235;
wire     [31:0] n37236;
wire     [31:0] n37237;
wire     [31:0] n37238;
wire     [31:0] n37239;
wire     [31:0] n37240;
wire     [31:0] n37241;
wire     [31:0] n37242;
wire     [31:0] n37243;
wire     [31:0] n37244;
wire     [31:0] n37245;
wire     [31:0] n37246;
wire     [31:0] n37247;
wire     [31:0] n37248;
wire     [31:0] n37249;
wire     [31:0] n37250;
wire     [31:0] n37251;
wire     [31:0] n37252;
wire     [31:0] n37253;
wire     [31:0] n37254;
wire     [31:0] n37255;
wire     [31:0] n37256;
wire     [31:0] n37257;
wire     [31:0] n37258;
wire     [31:0] n37259;
wire     [31:0] n37260;
wire     [31:0] n37261;
wire     [31:0] n37262;
wire     [31:0] n37263;
wire     [31:0] n37264;
wire     [31:0] n37265;
wire     [31:0] n37266;
wire     [31:0] n37267;
wire     [31:0] n37268;
wire     [31:0] n37269;
wire     [31:0] n37270;
wire     [31:0] n37271;
wire     [31:0] n37272;
wire     [31:0] n37273;
wire     [31:0] n37274;
wire     [31:0] n37275;
wire     [31:0] n37276;
wire     [31:0] n37277;
wire     [31:0] n37278;
wire     [31:0] n37279;
wire     [31:0] n37280;
wire     [31:0] n37281;
wire     [31:0] n37282;
wire     [31:0] n37283;
wire     [31:0] n37284;
wire     [31:0] n37285;
wire     [31:0] n37286;
wire     [31:0] n37287;
wire     [31:0] n37288;
wire     [31:0] n37289;
wire     [31:0] n37290;
wire     [31:0] n37291;
wire     [31:0] n37292;
wire     [31:0] n37293;
wire     [31:0] n37294;
wire     [31:0] n37295;
wire     [31:0] n37296;
wire     [31:0] n37297;
wire     [31:0] n37298;
wire     [31:0] n37299;
wire     [31:0] n37300;
wire     [31:0] n37301;
wire     [31:0] n37302;
wire     [31:0] n37303;
wire     [31:0] n37304;
wire     [31:0] n37305;
wire     [31:0] n37306;
wire     [31:0] n37307;
wire     [31:0] n37308;
wire     [31:0] n37309;
wire     [31:0] n37310;
wire     [31:0] n37311;
wire     [31:0] n37312;
wire     [31:0] n37313;
wire     [31:0] n37314;
wire     [31:0] n37315;
wire     [31:0] n37316;
wire     [31:0] n37317;
wire     [31:0] n37318;
wire     [31:0] n37319;
wire     [31:0] n37320;
wire     [31:0] n37321;
wire     [31:0] n37322;
wire     [31:0] n37323;
wire     [31:0] n37324;
wire     [31:0] n37325;
wire     [31:0] n37326;
wire     [31:0] n37327;
wire     [31:0] n37328;
wire     [31:0] n37329;
wire     [31:0] n37330;
wire     [31:0] n37331;
wire     [31:0] n37332;
wire     [31:0] n37333;
wire     [31:0] n37334;
wire     [31:0] n37335;
wire     [31:0] n37336;
wire     [31:0] n37337;
wire     [31:0] n37338;
wire     [31:0] n37339;
wire     [31:0] n37340;
wire     [31:0] n37341;
wire     [31:0] n37342;
wire     [31:0] n37343;
wire     [31:0] n37344;
wire     [31:0] n37345;
wire     [31:0] n37346;
wire     [31:0] n37347;
wire     [31:0] n37348;
wire     [31:0] n37349;
wire     [31:0] n37350;
wire     [31:0] n37351;
wire     [31:0] n37352;
wire     [31:0] n37353;
wire     [31:0] n37354;
wire     [31:0] n37355;
wire     [31:0] n37356;
wire     [31:0] n37357;
wire     [31:0] n37358;
wire     [31:0] n37359;
wire     [31:0] n37360;
wire     [31:0] n37361;
wire     [31:0] n37362;
wire     [31:0] n37363;
wire     [31:0] n37364;
wire     [31:0] n37365;
wire     [31:0] n37366;
wire     [31:0] n37367;
wire     [31:0] n37368;
wire     [31:0] n37369;
wire     [31:0] n37370;
wire     [31:0] n37371;
wire     [31:0] n37372;
wire     [31:0] n37373;
wire     [31:0] n37374;
wire     [31:0] n37375;
wire     [31:0] n37376;
wire     [31:0] n37377;
wire     [31:0] n37378;
wire     [31:0] n37379;
wire     [31:0] n37380;
wire     [31:0] n37381;
wire     [31:0] n37382;
wire     [31:0] n37383;
wire     [31:0] n37384;
wire     [31:0] n37385;
wire     [31:0] n37386;
wire     [31:0] n37387;
wire     [31:0] n37388;
wire     [31:0] n37389;
wire     [31:0] n37390;
wire     [31:0] n37391;
wire     [31:0] n37392;
wire     [31:0] n37393;
wire     [31:0] n37394;
wire     [31:0] n37395;
wire     [31:0] n37396;
wire     [31:0] n37397;
wire     [31:0] n37398;
wire     [31:0] n37399;
wire     [31:0] n37400;
wire     [31:0] n37401;
wire     [31:0] n37402;
wire     [31:0] n37403;
wire     [31:0] n37404;
wire     [31:0] n37405;
wire     [31:0] n37406;
wire     [31:0] n37407;
wire     [31:0] n37408;
wire     [31:0] n37409;
wire     [31:0] n37410;
wire     [31:0] n37411;
wire     [31:0] n37412;
wire     [31:0] n37413;
wire     [31:0] n37414;
wire     [31:0] n37415;
wire     [31:0] n37416;
wire     [31:0] n37417;
wire     [31:0] n37418;
wire     [31:0] n37419;
wire     [31:0] n37420;
wire     [31:0] n37421;
wire     [31:0] n37422;
wire     [31:0] n37423;
wire     [31:0] n37424;
wire     [31:0] n37425;
wire     [31:0] n37426;
wire     [31:0] n37427;
wire     [31:0] n37428;
wire     [31:0] n37429;
wire     [31:0] n37430;
wire     [31:0] n37431;
wire     [31:0] n37432;
wire     [31:0] n37433;
wire     [31:0] n37434;
wire     [31:0] n37435;
wire     [31:0] n37436;
wire     [31:0] n37437;
wire     [31:0] n37438;
wire     [31:0] n37439;
wire     [31:0] n37440;
wire     [31:0] n37441;
wire     [31:0] n37442;
wire     [31:0] n37443;
wire     [31:0] n37444;
wire     [31:0] n37445;
wire     [31:0] n37446;
wire     [31:0] n37447;
wire     [31:0] n37448;
wire     [31:0] n37449;
wire     [31:0] n37450;
wire     [31:0] n37451;
wire     [31:0] n37452;
wire     [31:0] n37453;
wire     [31:0] n37454;
wire     [31:0] n37455;
wire     [31:0] n37456;
wire     [31:0] n37457;
wire     [31:0] n37458;
wire     [31:0] n37459;
wire     [31:0] n37460;
wire     [31:0] n37461;
wire     [31:0] n37462;
wire     [31:0] n37463;
wire     [31:0] n37464;
wire     [31:0] n37465;
wire     [31:0] n37466;
wire     [31:0] n37467;
wire     [31:0] n37468;
wire     [31:0] n37469;
wire     [31:0] n37470;
wire     [31:0] n37471;
wire     [31:0] n37472;
wire     [31:0] n37473;
wire     [31:0] n37474;
wire     [31:0] n37475;
wire     [31:0] n37476;
wire     [31:0] n37477;
wire     [31:0] n37478;
wire     [31:0] n37479;
wire     [31:0] n37480;
wire     [31:0] n37481;
wire     [31:0] n37482;
wire     [31:0] n37483;
wire     [31:0] n37484;
wire     [31:0] n37485;
wire     [31:0] n37486;
wire     [31:0] n37487;
wire     [31:0] n37488;
wire     [31:0] n37489;
wire     [31:0] n37490;
wire     [31:0] n37491;
wire     [31:0] n37492;
wire     [31:0] n37493;
wire     [31:0] n37494;
wire     [31:0] n37495;
wire     [31:0] n37496;
wire     [31:0] n37497;
wire     [31:0] n37498;
wire     [31:0] n37499;
wire     [31:0] n37500;
wire     [31:0] n37501;
wire     [31:0] n37502;
wire     [31:0] n37503;
wire     [31:0] n37504;
wire     [31:0] n37505;
wire     [31:0] n37506;
wire     [31:0] n37507;
wire     [31:0] n37508;
wire     [31:0] n37509;
wire     [31:0] n37510;
wire     [31:0] n37511;
wire     [31:0] n37512;
wire     [31:0] n37513;
wire     [31:0] n37514;
wire     [31:0] n37515;
wire     [31:0] n37516;
wire     [31:0] n37517;
wire     [31:0] n37518;
wire     [31:0] n37519;
wire     [31:0] n37520;
wire     [31:0] n37521;
wire     [31:0] n37522;
wire     [31:0] n37523;
wire     [31:0] n37524;
wire     [31:0] n37525;
wire     [31:0] n37526;
wire     [31:0] n37527;
wire     [31:0] n37528;
wire     [31:0] n37529;
wire     [31:0] n37530;
wire     [31:0] n37531;
wire     [31:0] n37532;
wire     [31:0] n37533;
wire     [31:0] n37534;
wire     [31:0] n37535;
wire     [31:0] n37536;
wire     [31:0] n37537;
wire     [31:0] n37538;
wire     [31:0] n37539;
wire     [31:0] n37540;
wire     [31:0] n37541;
wire     [31:0] n37542;
wire     [31:0] n37543;
wire     [31:0] n37544;
wire     [31:0] n37545;
wire     [31:0] n37546;
wire     [31:0] n37547;
wire     [31:0] n37548;
wire     [31:0] n37549;
wire     [31:0] n37550;
wire     [31:0] n37551;
wire     [31:0] n37552;
wire     [31:0] n37553;
wire     [31:0] n37554;
wire     [31:0] n37555;
wire     [31:0] n37556;
wire     [31:0] n37557;
wire     [31:0] n37558;
wire     [31:0] n37559;
wire     [31:0] n37560;
wire     [31:0] n37561;
wire     [31:0] n37562;
wire     [31:0] n37563;
wire     [31:0] n37564;
wire     [31:0] n37565;
wire     [31:0] n37566;
wire     [31:0] n37567;
wire     [31:0] n37568;
wire     [31:0] n37569;
wire     [31:0] n37570;
wire     [31:0] n37571;
wire     [31:0] n37572;
wire     [31:0] n37573;
wire     [31:0] n37574;
wire     [31:0] n37575;
wire     [31:0] n37576;
wire     [31:0] n37577;
wire     [31:0] n37578;
wire     [31:0] n37579;
wire     [31:0] n37580;
wire     [31:0] n37581;
wire     [31:0] n37582;
wire     [31:0] n37583;
wire     [31:0] n37584;
wire     [31:0] n37585;
wire     [31:0] n37586;
wire     [31:0] n37587;
wire     [31:0] n37588;
wire     [31:0] n37589;
wire     [31:0] n37590;
wire     [31:0] n37591;
wire     [31:0] n37592;
wire     [31:0] n37593;
wire     [31:0] n37594;
wire     [31:0] n37595;
wire     [31:0] n37596;
wire     [31:0] n37597;
wire     [31:0] n37598;
wire     [31:0] n37599;
wire     [31:0] n37600;
wire     [31:0] n37601;
wire     [31:0] n37602;
wire     [31:0] n37603;
wire     [31:0] n37604;
wire     [31:0] n37605;
wire     [31:0] n37606;
wire     [31:0] n37607;
wire     [31:0] n37608;
wire     [31:0] n37609;
wire     [31:0] n37610;
wire     [31:0] n37611;
wire     [31:0] n37612;
wire     [31:0] n37613;
wire     [31:0] n37614;
wire     [31:0] n37615;
wire     [31:0] n37616;
wire     [31:0] n37617;
wire     [31:0] n37618;
wire     [31:0] n37619;
wire     [31:0] n37620;
wire     [31:0] n37621;
wire     [31:0] n37622;
wire     [31:0] n37623;
wire     [31:0] n37624;
wire     [31:0] n37625;
wire     [31:0] n37626;
wire     [31:0] n37627;
wire     [31:0] n37628;
wire     [31:0] n37629;
wire     [31:0] n37630;
wire     [31:0] n37631;
wire     [31:0] n37632;
wire     [31:0] n37633;
wire     [31:0] n37634;
wire     [31:0] n37635;
wire     [31:0] n37636;
wire     [31:0] n37637;
wire     [31:0] n37638;
wire     [31:0] n37639;
wire     [31:0] n37640;
wire     [31:0] n37641;
wire     [31:0] n37642;
wire     [31:0] n37643;
wire     [31:0] n37644;
wire     [31:0] n37645;
wire     [31:0] n37646;
wire     [31:0] n37647;
wire     [31:0] n37648;
wire     [31:0] n37649;
wire     [31:0] n37650;
wire     [31:0] n37651;
wire     [31:0] n37652;
wire     [31:0] n37653;
wire     [31:0] n37654;
wire     [31:0] n37655;
wire     [31:0] n37656;
wire     [31:0] n37657;
wire     [31:0] n37658;
wire     [31:0] n37659;
wire     [31:0] n37660;
wire     [31:0] n37661;
wire     [31:0] n37662;
wire     [31:0] n37663;
wire     [31:0] n37664;
wire     [31:0] n37665;
wire     [31:0] n37666;
wire     [31:0] n37667;
wire     [31:0] n37668;
wire     [31:0] n37669;
wire     [31:0] n37670;
wire     [31:0] n37671;
wire     [31:0] n37672;
wire     [31:0] n37673;
wire     [31:0] n37674;
wire     [31:0] n37675;
wire     [31:0] n37676;
wire     [31:0] n37677;
wire     [31:0] n37678;
wire     [31:0] n37679;
wire     [31:0] n37680;
wire     [31:0] n37681;
wire     [31:0] n37682;
wire     [31:0] n37683;
wire     [31:0] n37684;
wire     [31:0] n37685;
wire     [31:0] n37686;
wire     [31:0] n37687;
wire     [31:0] n37688;
wire     [31:0] n37689;
wire     [31:0] n37690;
wire     [31:0] n37691;
wire     [31:0] n37692;
wire     [31:0] n37693;
wire     [31:0] n37694;
wire     [31:0] n37695;
wire     [31:0] n37696;
wire     [31:0] n37697;
wire     [31:0] n37698;
wire     [31:0] n37699;
wire     [31:0] n37700;
wire     [31:0] n37701;
wire     [31:0] n37702;
wire     [31:0] n37703;
wire     [31:0] n37704;
wire     [31:0] n37705;
wire     [31:0] n37706;
wire     [31:0] n37707;
wire     [31:0] n37708;
wire     [31:0] n37709;
wire     [31:0] n37710;
wire     [31:0] n37711;
wire     [31:0] n37712;
wire     [31:0] n37713;
wire     [31:0] n37714;
wire     [31:0] n37715;
wire     [31:0] n37716;
wire     [31:0] n37717;
wire     [31:0] n37718;
wire     [31:0] n37719;
wire     [31:0] n37720;
wire     [31:0] n37721;
wire     [31:0] n37722;
wire     [31:0] n37723;
wire     [31:0] n37724;
wire     [31:0] n37725;
wire     [31:0] n37726;
wire     [31:0] n37727;
wire     [31:0] n37728;
wire     [31:0] n37729;
wire     [31:0] n37730;
wire     [31:0] n37731;
wire     [31:0] n37732;
wire     [31:0] n37733;
wire     [31:0] n37734;
wire     [31:0] n37735;
wire     [31:0] n37736;
wire     [31:0] n37737;
wire     [31:0] n37738;
wire     [31:0] n37739;
wire     [31:0] n37740;
wire     [31:0] n37741;
wire     [31:0] n37742;
wire     [31:0] n37743;
wire     [31:0] n37744;
wire     [31:0] n37745;
wire     [31:0] n37746;
wire     [31:0] n37747;
wire     [31:0] n37748;
wire     [31:0] n37749;
wire     [31:0] n37750;
wire     [31:0] n37751;
wire     [31:0] n37752;
wire     [31:0] n37753;
wire     [31:0] n37754;
wire     [31:0] n37755;
wire     [31:0] n37756;
wire     [31:0] n37757;
wire     [31:0] n37758;
wire     [31:0] n37759;
wire     [31:0] n37760;
wire     [31:0] n37761;
wire     [31:0] n37762;
wire     [31:0] n37763;
wire     [31:0] n37764;
wire     [31:0] n37765;
wire     [31:0] n37766;
wire     [31:0] n37767;
wire     [31:0] n37768;
wire     [31:0] n37769;
wire     [31:0] n37770;
wire     [31:0] n37771;
wire     [31:0] n37772;
wire     [31:0] n37773;
wire     [31:0] n37774;
wire     [31:0] n37775;
wire     [31:0] n37776;
wire     [31:0] n37777;
wire     [31:0] n37778;
wire     [31:0] n37779;
wire     [31:0] n37780;
wire     [31:0] n37781;
wire     [31:0] n37782;
wire     [31:0] n37783;
wire     [31:0] n37784;
wire     [31:0] n37785;
wire     [31:0] n37786;
wire     [31:0] n37787;
wire     [31:0] n37788;
wire     [31:0] n37789;
wire     [31:0] n37790;
wire     [31:0] n37791;
wire     [31:0] n37792;
wire     [31:0] n37793;
wire     [31:0] n37794;
wire     [31:0] n37795;
wire     [31:0] n37796;
wire     [31:0] n37797;
wire     [31:0] n37798;
wire     [31:0] n37799;
wire     [31:0] n37800;
wire     [31:0] n37801;
wire     [31:0] n37802;
wire     [31:0] n37803;
wire     [31:0] n37804;
wire     [31:0] n37805;
wire     [31:0] n37806;
wire     [31:0] n37807;
wire     [31:0] n37808;
wire     [31:0] n37809;
wire     [31:0] n37810;
wire     [31:0] n37811;
wire     [31:0] n37812;
wire     [31:0] n37813;
wire     [31:0] n37814;
wire     [31:0] n37815;
wire     [31:0] n37816;
wire     [31:0] n37817;
wire     [31:0] n37818;
wire     [31:0] n37819;
wire     [31:0] n37820;
wire     [31:0] n37821;
wire     [31:0] n37822;
wire     [31:0] n37823;
wire     [31:0] n37824;
wire     [31:0] n37825;
wire     [31:0] n37826;
wire     [31:0] n37827;
wire     [31:0] n37828;
wire     [31:0] n37829;
wire     [31:0] n37830;
wire     [31:0] n37831;
wire     [31:0] n37832;
wire     [31:0] n37833;
wire     [31:0] n37834;
wire     [31:0] n37835;
wire     [31:0] n37836;
wire     [31:0] n37837;
wire     [31:0] n37838;
wire     [31:0] n37839;
wire     [31:0] n37840;
wire     [31:0] n37841;
wire     [31:0] n37842;
wire     [31:0] n37843;
wire     [31:0] n37844;
wire     [31:0] n37845;
wire     [31:0] n37846;
wire     [31:0] n37847;
wire     [31:0] n37848;
wire     [31:0] n37849;
wire     [31:0] n37850;
wire     [31:0] n37851;
wire     [31:0] n37852;
wire     [31:0] n37853;
wire     [31:0] n37854;
wire     [31:0] n37855;
wire     [31:0] n37856;
wire     [31:0] n37857;
wire     [31:0] n37858;
wire     [31:0] n37859;
wire     [31:0] n37860;
wire     [31:0] n37861;
wire     [31:0] n37862;
wire     [31:0] n37863;
wire     [31:0] n37864;
wire     [31:0] n37865;
wire     [31:0] n37866;
wire     [31:0] n37867;
wire     [31:0] n37868;
wire     [31:0] n37869;
wire     [31:0] n37870;
wire     [31:0] n37871;
wire     [31:0] n37872;
wire     [31:0] n37873;
wire     [31:0] n37874;
wire     [31:0] n37875;
wire     [31:0] n37876;
wire     [31:0] n37877;
wire     [31:0] n37878;
wire     [31:0] n37879;
wire     [31:0] n37880;
wire     [31:0] n37881;
wire     [31:0] n37882;
wire     [31:0] n37883;
wire     [31:0] n37884;
wire     [31:0] n37885;
wire     [31:0] n37886;
wire     [31:0] n37887;
wire     [31:0] n37888;
wire     [31:0] n37889;
wire     [31:0] n37890;
wire     [31:0] n37891;
wire     [31:0] n37892;
wire     [31:0] n37893;
wire     [31:0] n37894;
wire     [31:0] n37895;
wire     [31:0] n37896;
wire     [31:0] n37897;
wire     [31:0] n37898;
wire     [31:0] n37899;
wire     [31:0] n37900;
wire     [31:0] n37901;
wire     [31:0] n37902;
wire     [31:0] n37903;
wire     [31:0] n37904;
wire     [31:0] n37905;
wire     [31:0] n37906;
wire     [31:0] n37907;
wire     [31:0] n37908;
wire     [31:0] n37909;
wire     [31:0] n37910;
wire     [31:0] n37911;
wire     [31:0] n37912;
wire     [31:0] n37913;
wire     [31:0] n37914;
wire     [31:0] n37915;
wire     [31:0] n37916;
wire     [31:0] n37917;
wire     [31:0] n37918;
wire     [31:0] n37919;
wire     [31:0] n37920;
wire     [31:0] n37921;
wire     [31:0] n37922;
wire     [31:0] n37923;
wire     [31:0] n37924;
wire     [31:0] n37925;
wire     [31:0] n37926;
wire     [31:0] n37927;
wire     [31:0] n37928;
wire     [31:0] n37929;
wire     [31:0] n37930;
wire     [31:0] n37931;
wire     [31:0] n37932;
wire     [31:0] n37933;
wire     [31:0] n37934;
wire     [31:0] n37935;
wire     [31:0] n37936;
wire     [31:0] n37937;
wire     [31:0] n37938;
wire     [31:0] n37939;
wire     [31:0] n37940;
wire     [31:0] n37941;
wire     [31:0] n37942;
wire     [31:0] n37943;
wire     [31:0] n37944;
wire     [31:0] n37945;
wire     [31:0] n37946;
wire     [31:0] n37947;
wire     [31:0] n37948;
wire     [31:0] n37949;
wire     [31:0] n37950;
wire     [31:0] n37951;
wire     [31:0] n37952;
wire     [31:0] n37953;
wire     [31:0] n37954;
wire     [31:0] n37955;
wire     [31:0] n37956;
wire     [31:0] n37957;
wire     [31:0] n37958;
wire     [31:0] n37959;
wire     [31:0] n37960;
wire     [31:0] n37961;
wire     [31:0] n37962;
wire     [31:0] n37963;
wire     [31:0] n37964;
wire     [31:0] n37965;
wire     [31:0] n37966;
wire     [31:0] n37967;
wire     [31:0] n37968;
wire     [31:0] n37969;
wire     [31:0] n37970;
wire     [31:0] n37971;
wire     [31:0] n37972;
wire     [31:0] n37973;
wire     [31:0] n37974;
wire     [31:0] n37975;
wire     [31:0] n37976;
wire     [31:0] n37977;
wire     [31:0] n37978;
wire     [31:0] n37979;
wire     [31:0] n37980;
wire     [31:0] n37981;
wire     [31:0] n37982;
wire     [31:0] n37983;
wire     [31:0] n37984;
wire     [31:0] n37985;
wire     [31:0] n37986;
wire     [31:0] n37987;
wire     [31:0] n37988;
wire     [31:0] n37989;
wire     [31:0] n37990;
wire     [31:0] n37991;
wire     [31:0] n37992;
wire     [31:0] n37993;
wire     [31:0] n37994;
wire     [31:0] n37995;
wire     [31:0] n37996;
wire     [31:0] n37997;
wire     [31:0] n37998;
wire     [31:0] n37999;
wire     [31:0] n38000;
wire     [31:0] n38001;
wire     [31:0] n38002;
wire     [31:0] n38003;
wire     [31:0] n38004;
wire     [31:0] n38005;
wire     [31:0] n38006;
wire     [31:0] n38007;
wire     [31:0] n38008;
wire     [31:0] n38009;
wire     [31:0] n38010;
wire     [31:0] n38011;
wire     [31:0] n38012;
wire     [31:0] n38013;
wire     [31:0] n38014;
wire     [31:0] n38015;
wire     [31:0] n38016;
wire     [31:0] n38017;
wire     [31:0] n38018;
wire     [31:0] n38019;
wire     [31:0] n38020;
wire     [31:0] n38021;
wire     [31:0] n38022;
wire     [31:0] n38023;
wire     [31:0] n38024;
wire     [31:0] n38025;
wire     [31:0] n38026;
wire     [31:0] n38027;
wire     [31:0] n38028;
wire     [31:0] n38029;
wire     [31:0] n38030;
wire     [31:0] n38031;
wire     [31:0] n38032;
wire     [31:0] n38033;
wire     [31:0] n38034;
wire     [31:0] n38035;
wire     [31:0] n38036;
wire     [31:0] n38037;
wire     [31:0] n38038;
wire     [31:0] n38039;
wire     [31:0] n38040;
wire     [31:0] n38041;
wire     [31:0] n38042;
wire     [31:0] n38043;
wire     [31:0] n38044;
wire     [31:0] n38045;
wire     [31:0] n38046;
wire     [31:0] n38047;
wire     [31:0] n38048;
wire     [31:0] n38049;
wire     [31:0] n38050;
wire     [31:0] n38051;
wire     [31:0] n38052;
wire     [31:0] n38053;
wire     [31:0] n38054;
wire     [31:0] n38055;
wire     [31:0] n38056;
wire     [31:0] n38057;
wire     [31:0] n38058;
wire     [31:0] n38059;
wire     [31:0] n38060;
wire     [31:0] n38061;
wire     [31:0] n38062;
wire     [31:0] n38063;
wire     [31:0] n38064;
wire     [31:0] n38065;
wire     [31:0] n38066;
wire     [31:0] n38067;
wire     [31:0] n38068;
wire     [31:0] n38069;
wire     [31:0] n38070;
wire     [31:0] n38071;
wire     [31:0] n38072;
wire     [31:0] n38073;
wire     [31:0] n38074;
wire     [31:0] n38075;
wire     [31:0] n38076;
wire     [31:0] n38077;
wire     [31:0] n38078;
wire     [31:0] n38079;
wire     [31:0] n38080;
wire     [31:0] n38081;
wire     [31:0] n38082;
wire     [31:0] n38083;
wire     [31:0] n38084;
wire     [31:0] n38085;
wire     [31:0] n38086;
wire     [31:0] n38087;
wire     [31:0] n38088;
wire     [31:0] n38089;
wire     [31:0] n38090;
wire     [31:0] n38091;
wire     [31:0] n38092;
wire     [31:0] n38093;
wire     [31:0] n38094;
wire     [31:0] n38095;
wire     [31:0] n38096;
wire     [31:0] n38097;
wire     [31:0] n38098;
wire     [31:0] n38099;
wire     [31:0] n38100;
wire     [31:0] n38101;
wire     [31:0] n38102;
wire     [31:0] n38103;
wire     [31:0] n38104;
wire     [31:0] n38105;
wire     [31:0] n38106;
wire     [31:0] n38107;
wire     [31:0] n38108;
wire     [31:0] n38109;
wire     [31:0] n38110;
wire     [31:0] n38111;
wire     [31:0] n38112;
wire     [31:0] n38113;
wire     [31:0] n38114;
wire     [31:0] n38115;
wire     [31:0] n38116;
wire     [31:0] n38117;
wire     [31:0] n38118;
wire     [31:0] n38119;
wire     [31:0] n38120;
wire     [31:0] n38121;
wire     [31:0] n38122;
wire     [31:0] n38123;
wire     [31:0] n38124;
wire     [31:0] n38125;
wire     [31:0] n38126;
wire     [31:0] n38127;
wire     [31:0] n38128;
wire     [31:0] n38129;
wire     [31:0] n38130;
wire     [31:0] n38131;
wire     [31:0] n38132;
wire     [31:0] n38133;
wire     [31:0] n38134;
wire     [31:0] n38135;
wire     [31:0] n38136;
wire     [31:0] n38137;
wire     [31:0] n38138;
wire     [31:0] n38139;
wire     [31:0] n38140;
wire     [31:0] n38141;
wire     [31:0] n38142;
wire     [31:0] n38143;
wire     [31:0] n38144;
wire     [31:0] n38145;
wire     [31:0] n38146;
wire     [31:0] n38147;
wire     [31:0] n38148;
wire     [31:0] n38149;
wire     [31:0] n38150;
wire     [31:0] n38151;
wire     [31:0] n38152;
wire     [31:0] n38153;
wire     [31:0] n38154;
wire     [31:0] n38155;
wire     [31:0] n38156;
wire     [31:0] n38157;
wire     [31:0] n38158;
wire     [31:0] n38159;
wire     [31:0] n38160;
wire     [31:0] n38161;
wire     [31:0] n38162;
wire     [31:0] n38163;
wire     [31:0] n38164;
wire     [31:0] n38165;
wire     [31:0] n38166;
wire     [31:0] n38167;
wire     [31:0] n38168;
wire     [31:0] n38169;
wire     [31:0] n38170;
wire     [31:0] n38171;
wire     [31:0] n38172;
wire     [31:0] n38173;
wire     [31:0] n38174;
wire     [31:0] n38175;
wire     [31:0] n38176;
wire     [31:0] n38177;
wire     [31:0] n38178;
wire     [31:0] n38179;
wire     [31:0] n38180;
wire     [31:0] n38181;
wire     [31:0] n38182;
wire     [31:0] n38183;
wire     [31:0] n38184;
wire     [31:0] n38185;
wire     [31:0] n38186;
wire     [31:0] n38187;
wire     [31:0] n38188;
wire     [31:0] n38189;
wire     [31:0] n38190;
wire     [31:0] n38191;
wire     [31:0] n38192;
wire     [31:0] n38193;
wire     [31:0] n38194;
wire     [31:0] n38195;
wire     [31:0] n38196;
wire     [31:0] n38197;
wire     [31:0] n38198;
wire     [31:0] n38199;
wire     [31:0] n38200;
wire     [31:0] n38201;
wire     [31:0] n38202;
wire     [31:0] n38203;
wire     [31:0] n38204;
wire     [31:0] n38205;
wire     [31:0] n38206;
wire     [31:0] n38207;
wire     [31:0] n38208;
wire     [31:0] n38209;
wire     [31:0] n38210;
wire     [31:0] n38211;
wire     [31:0] n38212;
wire     [31:0] n38213;
wire     [31:0] n38214;
wire     [31:0] n38215;
wire     [31:0] n38216;
wire     [31:0] n38217;
wire     [31:0] n38218;
wire     [31:0] n38219;
wire     [31:0] n38220;
wire     [31:0] n38221;
wire     [31:0] n38222;
wire     [31:0] n38223;
wire     [31:0] n38224;
wire     [31:0] n38225;
wire     [31:0] n38226;
wire     [31:0] n38227;
wire     [31:0] n38228;
wire     [31:0] n38229;
wire     [31:0] n38230;
wire     [31:0] n38231;
wire     [31:0] n38232;
wire     [31:0] n38233;
wire     [31:0] n38234;
wire     [31:0] n38235;
wire     [31:0] n38236;
wire     [31:0] n38237;
wire     [31:0] n38238;
wire     [31:0] n38239;
wire     [31:0] n38240;
wire     [31:0] n38241;
wire     [31:0] n38242;
wire     [31:0] n38243;
wire     [31:0] n38244;
wire     [31:0] n38245;
wire     [31:0] n38246;
wire     [31:0] n38247;
wire     [31:0] n38248;
wire     [31:0] n38249;
wire     [31:0] n38250;
wire     [31:0] n38251;
wire     [31:0] n38252;
wire     [31:0] n38253;
wire     [31:0] n38254;
wire     [31:0] n38255;
wire     [31:0] n38256;
wire     [31:0] n38257;
wire     [31:0] n38258;
wire     [31:0] n38259;
wire     [31:0] n38260;
wire     [31:0] n38261;
wire     [31:0] n38262;
wire     [31:0] n38263;
wire     [31:0] n38264;
wire     [31:0] n38265;
wire     [31:0] n38266;
wire     [31:0] n38267;
wire     [31:0] n38268;
wire     [31:0] n38269;
wire     [31:0] n38270;
wire     [31:0] n38271;
wire     [31:0] n38272;
wire     [31:0] n38273;
wire     [31:0] n38274;
wire     [31:0] n38275;
wire     [31:0] n38276;
wire     [31:0] n38277;
wire     [31:0] n38278;
wire     [31:0] n38279;
wire     [31:0] n38280;
wire     [31:0] n38281;
wire     [31:0] n38282;
wire     [31:0] n38283;
wire     [31:0] n38284;
wire     [31:0] n38285;
wire     [31:0] n38286;
wire     [31:0] n38287;
wire     [31:0] n38288;
wire     [31:0] n38289;
wire     [31:0] n38290;
wire     [31:0] n38291;
wire     [31:0] n38292;
wire     [31:0] n38293;
wire     [31:0] n38294;
wire     [31:0] n38295;
wire     [31:0] n38296;
wire     [31:0] n38297;
wire     [31:0] n38298;
wire     [31:0] n38299;
wire     [31:0] n38300;
wire     [31:0] n38301;
wire     [31:0] n38302;
wire     [31:0] n38303;
wire     [31:0] n38304;
wire     [31:0] n38305;
wire     [31:0] n38306;
wire     [31:0] n38307;
wire     [31:0] n38308;
wire     [31:0] n38309;
wire     [31:0] n38310;
wire     [31:0] n38311;
wire     [31:0] n38312;
wire     [31:0] n38313;
wire     [31:0] n38314;
wire     [31:0] n38315;
wire     [31:0] n38316;
wire     [31:0] n38317;
wire     [31:0] n38318;
wire     [31:0] n38319;
wire     [31:0] n38320;
wire     [31:0] n38321;
wire     [31:0] n38322;
wire     [31:0] n38323;
wire     [31:0] n38324;
wire     [31:0] n38325;
wire     [31:0] n38326;
wire     [31:0] n38327;
wire     [31:0] n38328;
wire     [31:0] n38329;
wire     [31:0] n38330;
wire     [31:0] n38331;
wire     [31:0] n38332;
wire     [31:0] n38333;
wire     [31:0] n38334;
wire     [31:0] n38335;
wire     [31:0] n38336;
wire     [31:0] n38337;
wire     [31:0] n38338;
wire     [31:0] n38339;
wire     [31:0] n38340;
wire     [31:0] n38341;
wire     [31:0] n38342;
wire     [31:0] n38343;
wire     [31:0] n38344;
wire     [31:0] n38345;
wire     [31:0] n38346;
wire     [31:0] n38347;
wire     [31:0] n38348;
wire     [31:0] n38349;
wire     [31:0] n38350;
wire     [31:0] n38351;
wire     [31:0] n38352;
wire     [31:0] n38353;
wire     [31:0] n38354;
wire     [31:0] n38355;
wire     [31:0] n38356;
wire     [31:0] n38357;
wire     [31:0] n38358;
wire     [31:0] n38359;
wire     [31:0] n38360;
wire     [31:0] n38361;
wire     [31:0] n38362;
wire     [31:0] n38363;
wire     [31:0] n38364;
wire     [31:0] n38365;
wire     [31:0] n38366;
wire     [31:0] n38367;
wire     [31:0] n38368;
wire     [31:0] n38369;
wire     [31:0] n38370;
wire     [31:0] n38371;
wire     [31:0] n38372;
wire     [31:0] n38373;
wire     [31:0] n38374;
wire     [31:0] n38375;
wire     [31:0] n38376;
wire     [31:0] n38377;
wire     [31:0] n38378;
wire     [31:0] n38379;
wire     [31:0] n38380;
wire     [31:0] n38381;
wire     [31:0] n38382;
wire     [31:0] n38383;
wire     [31:0] n38384;
wire     [31:0] n38385;
wire     [31:0] n38386;
wire     [31:0] n38387;
wire     [31:0] n38388;
wire     [31:0] n38389;
wire     [31:0] n38390;
wire     [31:0] n38391;
wire     [31:0] n38392;
wire     [31:0] n38393;
wire     [31:0] n38394;
wire     [31:0] n38395;
wire     [31:0] n38396;
wire     [31:0] n38397;
wire     [31:0] n38398;
wire     [31:0] n38399;
wire     [31:0] n38400;
wire     [31:0] n38401;
wire     [31:0] n38402;
wire     [31:0] n38403;
wire     [31:0] n38404;
wire     [31:0] n38405;
wire     [31:0] n38406;
wire     [31:0] n38407;
wire     [31:0] n38408;
wire     [31:0] n38409;
wire     [31:0] n38410;
wire     [31:0] n38411;
wire     [31:0] n38412;
wire     [31:0] n38413;
wire     [31:0] n38414;
wire     [31:0] n38415;
wire     [31:0] n38416;
wire     [31:0] n38417;
wire     [31:0] n38418;
wire     [31:0] n38419;
wire     [31:0] n38420;
wire     [31:0] n38421;
wire     [31:0] n38422;
wire     [31:0] n38423;
wire     [31:0] n38424;
wire     [31:0] n38425;
wire     [31:0] n38426;
wire     [31:0] n38427;
wire     [31:0] n38428;
wire     [31:0] n38429;
wire     [31:0] n38430;
wire     [31:0] n38431;
wire     [31:0] n38432;
wire     [31:0] n38433;
wire     [31:0] n38434;
wire     [31:0] n38435;
wire     [31:0] n38436;
wire     [31:0] n38437;
wire     [31:0] n38438;
wire     [31:0] n38439;
wire     [31:0] n38440;
wire     [31:0] n38441;
wire     [31:0] n38442;
wire     [31:0] n38443;
wire     [31:0] n38444;
wire     [31:0] n38445;
wire     [31:0] n38446;
wire     [31:0] n38447;
wire     [31:0] n38448;
wire     [31:0] n38449;
wire     [31:0] n38450;
wire     [31:0] n38451;
wire     [31:0] n38452;
wire     [31:0] n38453;
wire     [31:0] n38454;
wire     [31:0] n38455;
wire     [31:0] n38456;
wire     [31:0] n38457;
wire     [31:0] n38458;
wire     [31:0] n38459;
wire     [31:0] n38460;
wire     [31:0] n38461;
wire     [31:0] n38462;
wire     [31:0] n38463;
wire     [31:0] n38464;
wire     [31:0] n38465;
wire     [31:0] n38466;
wire     [31:0] n38467;
wire     [31:0] n38468;
wire     [31:0] n38469;
wire     [31:0] n38470;
wire     [31:0] n38471;
wire     [31:0] n38472;
wire     [31:0] n38473;
wire     [31:0] n38474;
wire     [31:0] n38475;
wire     [31:0] n38476;
wire     [31:0] n38477;
wire     [31:0] n38478;
wire     [31:0] n38479;
wire     [31:0] n38480;
wire     [31:0] n38481;
wire     [31:0] n38482;
wire     [31:0] n38483;
wire     [31:0] n38484;
wire     [31:0] n38485;
wire     [31:0] n38486;
wire     [31:0] n38487;
wire     [31:0] n38488;
wire     [31:0] n38489;
wire     [31:0] n38490;
wire     [31:0] n38491;
wire     [31:0] n38492;
wire     [31:0] n38493;
wire     [31:0] n38494;
wire     [31:0] n38495;
wire     [31:0] n38496;
wire     [31:0] n38497;
wire     [31:0] n38498;
wire     [31:0] n38499;
wire     [31:0] n38500;
wire     [31:0] n38501;
wire     [31:0] n38502;
wire     [31:0] n38503;
wire     [31:0] n38504;
wire     [31:0] n38505;
wire     [31:0] n38506;
wire     [31:0] n38507;
wire     [31:0] n38508;
wire     [31:0] n38509;
wire     [31:0] n38510;
wire     [31:0] n38511;
wire     [31:0] n38512;
wire     [31:0] n38513;
wire     [31:0] n38514;
wire     [31:0] n38515;
wire     [31:0] n38516;
wire     [31:0] n38517;
wire     [31:0] n38518;
wire     [31:0] n38519;
wire     [31:0] n38520;
wire     [31:0] n38521;
wire     [31:0] n38522;
wire     [31:0] n38523;
wire     [31:0] n38524;
wire     [31:0] n38525;
wire     [31:0] n38526;
wire     [31:0] n38527;
wire     [31:0] n38528;
wire     [31:0] n38529;
wire     [31:0] n38530;
wire     [31:0] n38531;
wire     [31:0] n38532;
wire     [31:0] n38533;
wire     [31:0] n38534;
wire     [31:0] n38535;
wire     [31:0] n38536;
wire     [31:0] n38537;
wire     [31:0] n38538;
wire     [31:0] n38539;
wire     [31:0] n38540;
wire     [31:0] n38541;
wire     [31:0] n38542;
wire     [31:0] n38543;
wire     [31:0] n38544;
wire     [31:0] n38545;
wire     [31:0] n38546;
wire     [31:0] n38547;
wire     [31:0] n38548;
wire     [31:0] n38549;
wire     [31:0] n38550;
wire     [31:0] n38551;
wire     [31:0] n38552;
wire     [31:0] n38553;
wire     [31:0] n38554;
wire     [31:0] n38555;
wire     [31:0] n38556;
wire     [31:0] n38557;
wire     [31:0] n38558;
wire     [31:0] n38559;
wire     [31:0] n38560;
wire     [31:0] n38561;
wire     [31:0] n38562;
wire     [31:0] n38563;
wire     [31:0] n38564;
wire     [31:0] n38565;
wire     [31:0] n38566;
wire     [31:0] n38567;
wire     [31:0] n38568;
wire     [31:0] n38569;
wire     [31:0] n38570;
wire     [31:0] n38571;
wire     [31:0] n38572;
wire     [31:0] n38573;
wire     [31:0] n38574;
wire     [31:0] n38575;
wire     [31:0] n38576;
wire     [31:0] n38577;
wire     [31:0] n38578;
wire     [31:0] n38579;
wire     [31:0] n38580;
wire     [31:0] n38581;
wire     [31:0] n38582;
wire     [31:0] n38583;
wire     [31:0] n38584;
wire     [31:0] n38585;
wire     [31:0] n38586;
wire     [31:0] n38587;
wire     [31:0] n38588;
wire     [31:0] n38589;
wire     [31:0] n38590;
wire     [31:0] n38591;
wire     [31:0] n38592;
wire     [31:0] n38593;
wire     [31:0] n38594;
wire     [31:0] n38595;
wire     [31:0] n38596;
wire     [31:0] n38597;
wire     [31:0] n38598;
wire     [31:0] n38599;
wire     [31:0] n38600;
wire     [31:0] n38601;
wire     [31:0] n38602;
wire     [31:0] n38603;
wire     [31:0] n38604;
wire     [31:0] n38605;
wire     [31:0] n38606;
wire     [31:0] n38607;
wire     [31:0] n38608;
wire     [31:0] n38609;
wire     [31:0] n38610;
wire     [31:0] n38611;
wire     [31:0] n38612;
wire     [31:0] n38613;
wire     [31:0] n38614;
wire     [31:0] n38615;
wire     [31:0] n38616;
wire     [31:0] n38617;
wire     [31:0] n38618;
wire     [31:0] n38619;
wire     [31:0] n38620;
wire     [31:0] n38621;
wire     [31:0] n38622;
wire     [31:0] n38623;
wire     [31:0] n38624;
wire     [31:0] n38625;
wire     [31:0] n38626;
wire     [31:0] n38627;
wire     [31:0] n38628;
wire     [31:0] n38629;
wire     [31:0] n38630;
wire     [31:0] n38631;
wire     [31:0] n38632;
wire     [31:0] n38633;
wire     [31:0] n38634;
wire     [31:0] n38635;
wire     [31:0] n38636;
wire     [31:0] n38637;
wire     [31:0] n38638;
wire     [31:0] n38639;
wire     [31:0] n38640;
wire     [31:0] n38641;
wire     [31:0] n38642;
wire     [31:0] n38643;
wire     [31:0] n38644;
wire     [31:0] n38645;
wire     [31:0] n38646;
wire     [31:0] n38647;
wire     [31:0] n38648;
wire     [31:0] n38649;
wire     [31:0] n38650;
wire     [31:0] n38651;
wire     [31:0] n38652;
wire     [31:0] n38653;
wire     [31:0] n38654;
wire     [31:0] n38655;
wire     [31:0] n38656;
wire     [31:0] n38657;
wire     [31:0] n38658;
wire     [31:0] n38659;
wire     [31:0] n38660;
wire     [31:0] n38661;
wire     [31:0] n38662;
wire     [31:0] n38663;
wire     [31:0] n38664;
wire     [31:0] n38665;
wire     [31:0] n38666;
wire     [31:0] n38667;
wire     [31:0] n38668;
wire     [31:0] n38669;
wire     [31:0] n38670;
wire     [31:0] n38671;
wire     [31:0] n38672;
wire     [31:0] n38673;
wire     [31:0] n38674;
wire     [31:0] n38675;
wire     [31:0] n38676;
wire     [31:0] n38677;
wire     [31:0] n38678;
wire     [31:0] n38679;
wire     [31:0] n38680;
wire     [31:0] n38681;
wire     [31:0] n38682;
wire     [31:0] n38683;
wire     [31:0] n38684;
wire     [31:0] n38685;
wire     [31:0] n38686;
wire     [31:0] n38687;
wire     [31:0] n38688;
wire     [31:0] n38689;
wire     [31:0] n38690;
wire     [31:0] n38691;
wire     [31:0] n38692;
wire     [31:0] n38693;
wire     [31:0] n38694;
wire     [31:0] n38695;
wire     [31:0] n38696;
wire     [31:0] n38697;
wire     [31:0] n38698;
wire     [31:0] n38699;
wire     [31:0] n38700;
wire     [31:0] n38701;
wire     [31:0] n38702;
wire     [31:0] n38703;
wire     [31:0] n38704;
wire     [31:0] n38705;
wire     [31:0] n38706;
wire     [31:0] n38707;
wire     [31:0] n38708;
wire     [31:0] n38709;
wire     [31:0] n38710;
wire     [31:0] n38711;
wire     [31:0] n38712;
wire     [31:0] n38713;
wire     [31:0] n38714;
wire     [31:0] n38715;
wire     [31:0] n38716;
wire     [31:0] n38717;
wire     [31:0] n38718;
wire     [31:0] n38719;
wire     [31:0] n38720;
wire     [31:0] n38721;
wire     [31:0] n38722;
wire     [31:0] n38723;
wire     [31:0] n38724;
wire     [31:0] n38725;
wire     [31:0] n38726;
wire     [31:0] n38727;
wire     [31:0] n38728;
wire     [31:0] n38729;
wire     [31:0] n38730;
wire     [31:0] n38731;
wire     [31:0] n38732;
wire     [31:0] n38733;
wire     [31:0] n38734;
wire     [31:0] n38735;
wire     [31:0] n38736;
wire     [31:0] n38737;
wire     [31:0] n38738;
wire     [31:0] n38739;
wire     [31:0] n38740;
wire     [31:0] n38741;
wire     [31:0] n38742;
wire     [31:0] n38743;
wire     [31:0] n38744;
wire     [31:0] n38745;
wire     [31:0] n38746;
wire     [31:0] n38747;
wire     [31:0] n38748;
wire     [31:0] n38749;
wire     [31:0] n38750;
wire     [31:0] n38751;
wire     [31:0] n38752;
wire     [31:0] n38753;
wire     [31:0] n38754;
wire     [31:0] n38755;
wire     [31:0] n38756;
wire     [31:0] n38757;
wire     [31:0] n38758;
wire     [31:0] n38759;
wire     [31:0] n38760;
wire     [31:0] n38761;
wire     [31:0] n38762;
wire     [31:0] n38763;
wire     [31:0] n38764;
wire     [31:0] n38765;
wire     [31:0] n38766;
wire     [31:0] n38767;
wire     [31:0] n38768;
wire     [31:0] n38769;
wire     [31:0] n38770;
wire     [31:0] n38771;
wire     [31:0] n38772;
wire     [31:0] n38773;
wire     [31:0] n38774;
wire     [31:0] n38775;
wire     [31:0] n38776;
wire     [31:0] n38777;
wire     [31:0] n38778;
wire     [31:0] n38779;
wire     [31:0] n38780;
wire     [31:0] n38781;
wire     [31:0] n38782;
wire     [31:0] n38783;
wire     [31:0] n38784;
wire     [31:0] n38785;
wire     [31:0] n38786;
wire     [31:0] n38787;
wire     [31:0] n38788;
wire     [31:0] n38789;
wire     [31:0] n38790;
wire     [31:0] n38791;
wire     [31:0] n38792;
wire     [31:0] n38793;
wire     [31:0] n38794;
wire     [31:0] n38795;
wire     [31:0] n38796;
wire     [31:0] n38797;
wire     [31:0] n38798;
wire     [31:0] n38799;
wire     [31:0] n38800;
wire     [31:0] n38801;
wire     [31:0] n38802;
wire     [31:0] n38803;
wire     [31:0] n38804;
wire     [31:0] n38805;
wire     [31:0] n38806;
wire     [31:0] n38807;
wire     [31:0] n38808;
wire     [31:0] n38809;
wire     [31:0] n38810;
wire     [31:0] n38811;
wire     [31:0] n38812;
wire     [31:0] n38813;
wire     [31:0] n38814;
wire     [31:0] n38815;
wire     [31:0] n38816;
wire     [31:0] n38817;
wire     [31:0] n38818;
wire     [31:0] n38819;
wire     [31:0] n38820;
wire     [31:0] n38821;
wire     [31:0] n38822;
wire     [31:0] n38823;
wire     [31:0] n38824;
wire     [31:0] n38825;
wire     [31:0] n38826;
wire     [31:0] n38827;
wire     [31:0] n38828;
wire     [31:0] n38829;
wire     [31:0] n38830;
wire     [31:0] n38831;
wire     [31:0] n38832;
wire     [31:0] n38833;
wire     [31:0] n38834;
wire     [31:0] n38835;
wire     [31:0] n38836;
wire     [31:0] n38837;
wire     [31:0] n38838;
wire     [31:0] n38839;
wire     [31:0] n38840;
wire     [31:0] n38841;
wire     [31:0] n38842;
wire     [31:0] n38843;
wire     [31:0] n38844;
wire     [31:0] n38845;
wire     [31:0] n38846;
wire     [31:0] n38847;
wire     [31:0] n38848;
wire     [31:0] n38849;
wire     [31:0] n38850;
wire     [31:0] n38851;
wire     [31:0] n38852;
wire     [31:0] n38853;
wire     [31:0] n38854;
wire     [31:0] n38855;
wire     [31:0] n38856;
wire     [31:0] n38857;
wire     [31:0] n38858;
wire     [31:0] n38859;
wire     [31:0] n38860;
wire     [31:0] n38861;
wire     [31:0] n38862;
wire     [31:0] n38863;
wire     [31:0] n38864;
wire     [31:0] n38865;
wire     [31:0] n38866;
wire     [31:0] n38867;
wire     [31:0] n38868;
wire     [31:0] n38869;
wire     [31:0] n38870;
wire     [31:0] n38871;
wire     [31:0] n38872;
wire     [31:0] n38873;
wire     [31:0] n38874;
wire     [31:0] n38875;
wire     [31:0] n38876;
wire     [31:0] n38877;
wire     [31:0] n38878;
wire     [31:0] n38879;
wire     [31:0] n38880;
wire     [31:0] n38881;
wire     [31:0] n38882;
wire     [31:0] n38883;
wire     [31:0] n38884;
wire     [31:0] n38885;
wire     [31:0] n38886;
wire     [31:0] n38887;
wire     [31:0] n38888;
wire     [31:0] n38889;
wire     [31:0] n38890;
wire     [31:0] n38891;
wire     [31:0] n38892;
wire     [31:0] n38893;
wire     [31:0] n38894;
wire     [31:0] n38895;
wire     [31:0] n38896;
wire     [31:0] n38897;
wire     [31:0] n38898;
wire     [31:0] n38899;
wire     [31:0] n38900;
wire     [31:0] n38901;
wire     [31:0] n38902;
wire     [31:0] n38903;
wire     [31:0] n38904;
wire     [31:0] n38905;
wire     [31:0] n38906;
wire     [31:0] n38907;
wire     [31:0] n38908;
wire     [31:0] n38909;
wire     [31:0] n38910;
wire     [31:0] n38911;
wire     [31:0] n38912;
wire     [31:0] n38913;
wire     [31:0] n38914;
wire     [31:0] n38915;
wire     [31:0] n38916;
wire     [31:0] n38917;
wire     [31:0] n38918;
wire     [31:0] n38919;
wire     [31:0] n38920;
wire     [31:0] n38921;
wire     [31:0] n38922;
wire     [31:0] n38923;
wire     [31:0] n38924;
wire     [31:0] n38925;
wire     [31:0] n38926;
wire     [31:0] n38927;
wire     [31:0] n38928;
wire     [31:0] n38929;
wire     [31:0] n38930;
wire     [31:0] n38931;
wire     [31:0] n38932;
wire     [31:0] n38933;
wire     [31:0] n38934;
wire     [31:0] n38935;
wire     [31:0] n38936;
wire     [31:0] n38937;
wire     [31:0] n38938;
wire     [31:0] n38939;
wire     [31:0] n38940;
wire     [31:0] n38941;
wire     [31:0] n38942;
wire     [31:0] n38943;
wire     [31:0] n38944;
wire     [31:0] n38945;
wire     [31:0] n38946;
wire     [31:0] n38947;
wire     [31:0] n38948;
wire     [31:0] n38949;
wire     [31:0] n38950;
wire     [31:0] n38951;
wire     [31:0] n38952;
wire     [31:0] n38953;
wire     [31:0] n38954;
wire     [31:0] n38955;
wire     [31:0] n38956;
wire     [31:0] n38957;
wire     [31:0] n38958;
wire     [31:0] n38959;
wire     [31:0] n38960;
wire     [31:0] n38961;
wire     [31:0] n38962;
wire     [31:0] n38963;
wire     [31:0] n38964;
wire     [31:0] n38965;
wire     [31:0] n38966;
wire     [31:0] n38967;
wire     [31:0] n38968;
wire     [31:0] n38969;
wire     [31:0] n38970;
wire     [31:0] n38971;
wire     [31:0] n38972;
wire     [31:0] n38973;
wire     [31:0] n38974;
wire     [31:0] n38975;
wire     [31:0] n38976;
wire     [31:0] n38977;
wire     [31:0] n38978;
wire     [31:0] n38979;
wire     [31:0] n38980;
wire     [31:0] n38981;
wire     [31:0] n38982;
wire     [31:0] n38983;
wire     [31:0] n38984;
wire     [31:0] n38985;
wire     [31:0] n38986;
wire     [31:0] n38987;
wire     [31:0] n38988;
wire     [31:0] n38989;
wire     [31:0] n38990;
wire     [31:0] n38991;
wire     [31:0] n38992;
wire     [31:0] n38993;
wire     [31:0] n38994;
wire     [31:0] n38995;
wire     [31:0] n38996;
wire     [31:0] n38997;
wire     [31:0] n38998;
wire     [31:0] n38999;
wire     [31:0] n39000;
wire     [31:0] n39001;
wire     [31:0] n39002;
wire     [31:0] n39003;
wire     [31:0] n39004;
wire     [31:0] n39005;
wire     [31:0] n39006;
wire     [31:0] n39007;
wire     [31:0] n39008;
wire     [31:0] n39009;
wire     [31:0] n39010;
wire     [31:0] n39011;
wire     [31:0] n39012;
wire     [31:0] n39013;
wire     [31:0] n39014;
wire     [31:0] n39015;
wire     [31:0] n39016;
wire     [31:0] n39017;
wire     [31:0] n39018;
wire     [31:0] n39019;
wire     [31:0] n39020;
wire     [31:0] n39021;
wire     [31:0] n39022;
wire     [31:0] n39023;
wire     [31:0] n39024;
wire     [31:0] n39025;
wire     [31:0] n39026;
wire     [31:0] n39027;
wire     [31:0] n39028;
wire     [31:0] n39029;
wire     [31:0] n39030;
wire     [31:0] n39031;
wire     [31:0] n39032;
wire     [31:0] n39033;
wire     [31:0] n39034;
wire     [31:0] n39035;
wire     [31:0] n39036;
wire     [31:0] n39037;
wire     [31:0] n39038;
wire     [31:0] n39039;
wire     [31:0] n39040;
wire     [31:0] n39041;
wire     [31:0] n39042;
wire     [31:0] n39043;
wire     [31:0] n39044;
wire     [31:0] n39045;
wire     [31:0] n39046;
wire     [31:0] n39047;
wire     [31:0] n39048;
wire     [31:0] n39049;
wire     [31:0] n39050;
wire     [31:0] n39051;
wire     [31:0] n39052;
wire     [31:0] n39053;
wire     [31:0] n39054;
wire     [31:0] n39055;
wire     [31:0] n39056;
wire     [31:0] n39057;
wire     [31:0] n39058;
wire     [31:0] n39059;
wire     [31:0] n39060;
wire     [31:0] n39061;
wire     [31:0] n39062;
wire     [31:0] n39063;
wire     [31:0] n39064;
wire     [31:0] n39065;
wire     [31:0] n39066;
wire     [31:0] n39067;
wire     [31:0] n39068;
wire     [31:0] n39069;
wire     [31:0] n39070;
wire     [31:0] n39071;
wire     [31:0] n39072;
wire     [31:0] n39073;
wire     [31:0] n39074;
wire     [31:0] n39075;
wire     [31:0] n39076;
wire     [31:0] n39077;
wire     [31:0] n39078;
wire     [31:0] n39079;
wire     [31:0] n39080;
wire     [31:0] n39081;
wire     [31:0] n39082;
wire     [31:0] n39083;
wire     [31:0] n39084;
wire     [31:0] n39085;
wire     [31:0] n39086;
wire     [31:0] n39087;
wire     [31:0] n39088;
wire     [31:0] n39089;
wire     [31:0] n39090;
wire     [31:0] n39091;
wire     [31:0] n39092;
wire     [31:0] n39093;
wire     [31:0] n39094;
wire     [31:0] n39095;
wire     [31:0] n39096;
wire     [31:0] n39097;
wire     [31:0] n39098;
wire     [31:0] n39099;
wire     [31:0] n39100;
wire     [31:0] n39101;
wire     [31:0] n39102;
wire     [31:0] n39103;
wire     [31:0] n39104;
wire     [31:0] n39105;
wire     [31:0] n39106;
wire     [31:0] n39107;
wire     [31:0] n39108;
wire     [31:0] n39109;
wire     [31:0] n39110;
wire     [31:0] n39111;
wire     [31:0] n39112;
wire     [31:0] n39113;
wire     [31:0] n39114;
wire     [31:0] n39115;
wire     [31:0] n39116;
wire     [31:0] n39117;
wire     [31:0] n39118;
wire     [31:0] n39119;
wire     [31:0] n39120;
wire     [31:0] n39121;
wire     [31:0] n39122;
wire     [31:0] n39123;
wire     [31:0] n39124;
wire     [31:0] n39125;
wire     [31:0] n39126;
wire     [31:0] n39127;
wire     [31:0] n39128;
wire     [31:0] n39129;
wire     [31:0] n39130;
wire     [31:0] n39131;
wire     [31:0] n39132;
wire     [31:0] n39133;
wire     [31:0] n39134;
wire     [31:0] n39135;
wire     [31:0] n39136;
wire     [31:0] n39137;
wire     [31:0] n39138;
wire     [31:0] n39139;
wire     [31:0] n39140;
wire     [31:0] n39141;
wire     [31:0] n39142;
wire     [31:0] n39143;
wire     [31:0] n39144;
wire     [31:0] n39145;
wire     [31:0] n39146;
wire     [31:0] n39147;
wire     [31:0] n39148;
wire     [31:0] n39149;
wire     [31:0] n39150;
wire     [31:0] n39151;
wire     [31:0] n39152;
wire     [31:0] n39153;
wire     [31:0] n39154;
wire     [31:0] n39155;
wire     [31:0] n39156;
wire     [31:0] n39157;
wire     [31:0] n39158;
wire     [31:0] n39159;
wire     [31:0] n39160;
wire     [31:0] n39161;
wire     [31:0] n39162;
wire     [31:0] n39163;
wire     [31:0] n39164;
wire     [31:0] n39165;
wire     [31:0] n39166;
wire     [31:0] n39167;
wire     [31:0] n39168;
wire     [31:0] n39169;
wire     [31:0] n39170;
wire     [31:0] n39171;
wire     [31:0] n39172;
wire     [31:0] n39173;
wire     [31:0] n39174;
wire     [31:0] n39175;
wire     [31:0] n39176;
wire     [31:0] n39177;
wire     [31:0] n39178;
wire     [31:0] n39179;
wire     [31:0] n39180;
wire     [31:0] n39181;
wire     [31:0] n39182;
wire     [31:0] n39183;
wire     [31:0] n39184;
wire     [31:0] n39185;
wire     [31:0] n39186;
wire     [31:0] n39187;
wire     [31:0] n39188;
wire     [31:0] n39189;
wire     [31:0] n39190;
wire     [31:0] n39191;
wire     [31:0] n39192;
wire     [31:0] n39193;
wire     [31:0] n39194;
wire     [31:0] n39195;
wire     [31:0] n39196;
wire     [31:0] n39197;
wire     [31:0] n39198;
wire     [31:0] n39199;
wire     [31:0] n39200;
wire     [31:0] n39201;
wire     [31:0] n39202;
wire     [31:0] n39203;
wire     [31:0] n39204;
wire     [31:0] n39205;
wire     [31:0] n39206;
wire     [31:0] n39207;
wire     [31:0] n39208;
wire     [31:0] n39209;
wire     [31:0] n39210;
wire     [31:0] n39211;
wire     [31:0] n39212;
wire     [31:0] n39213;
wire     [31:0] n39214;
wire     [31:0] n39215;
wire     [31:0] n39216;
wire     [31:0] n39217;
wire     [31:0] n39218;
wire     [31:0] n39219;
wire     [31:0] n39220;
wire     [31:0] n39221;
wire     [31:0] n39222;
wire     [31:0] n39223;
wire     [31:0] n39224;
wire     [31:0] n39225;
wire     [31:0] n39226;
wire     [31:0] n39227;
wire     [31:0] n39228;
wire     [31:0] n39229;
wire     [31:0] n39230;
wire     [31:0] n39231;
wire     [31:0] n39232;
wire     [31:0] n39233;
wire     [31:0] n39234;
wire     [31:0] n39235;
wire     [31:0] n39236;
wire     [31:0] n39237;
wire     [31:0] n39238;
wire     [31:0] n39239;
wire     [31:0] n39240;
wire     [31:0] n39241;
wire     [31:0] n39242;
wire     [31:0] n39243;
wire     [31:0] n39244;
wire     [31:0] n39245;
wire     [31:0] n39246;
wire     [31:0] n39247;
wire     [31:0] n39248;
wire     [31:0] n39249;
wire     [31:0] n39250;
wire     [31:0] n39251;
wire     [31:0] n39252;
wire     [31:0] n39253;
wire     [31:0] n39254;
wire     [31:0] n39255;
wire     [31:0] n39256;
wire     [31:0] n39257;
wire     [31:0] n39258;
wire     [31:0] n39259;
wire     [31:0] n39260;
wire     [31:0] n39261;
wire     [31:0] n39262;
wire     [31:0] n39263;
wire     [31:0] n39264;
wire     [31:0] n39265;
wire     [31:0] n39266;
wire     [31:0] n39267;
wire     [31:0] n39268;
wire     [31:0] n39269;
wire     [31:0] n39270;
wire     [31:0] n39271;
wire     [31:0] n39272;
wire     [31:0] n39273;
wire     [31:0] n39274;
wire     [31:0] n39275;
wire     [31:0] n39276;
wire     [31:0] n39277;
wire     [31:0] n39278;
wire     [31:0] n39279;
wire     [31:0] n39280;
wire     [31:0] n39281;
wire     [31:0] n39282;
wire     [31:0] n39283;
wire     [31:0] n39284;
wire     [31:0] n39285;
wire     [31:0] n39286;
wire     [31:0] n39287;
wire     [31:0] n39288;
wire     [31:0] n39289;
wire     [31:0] n39290;
wire     [31:0] n39291;
wire     [31:0] n39292;
wire     [31:0] n39293;
wire     [31:0] n39294;
wire     [31:0] n39295;
wire     [31:0] n39296;
wire     [31:0] n39297;
wire     [31:0] n39298;
wire     [31:0] n39299;
wire     [31:0] n39300;
wire     [31:0] n39301;
wire     [31:0] n39302;
wire     [31:0] n39303;
wire     [31:0] n39304;
wire     [31:0] n39305;
wire     [31:0] n39306;
wire     [31:0] n39307;
wire     [31:0] n39308;
wire     [31:0] n39309;
wire     [31:0] n39310;
wire     [31:0] n39311;
wire     [31:0] n39312;
wire     [31:0] n39313;
wire     [31:0] n39314;
wire     [31:0] n39315;
wire     [31:0] n39316;
wire     [31:0] n39317;
wire     [31:0] n39318;
wire     [31:0] n39319;
wire     [31:0] n39320;
wire     [31:0] n39321;
wire     [31:0] n39322;
wire     [31:0] n39323;
wire     [31:0] n39324;
wire     [31:0] n39325;
wire     [31:0] n39326;
wire     [31:0] n39327;
wire     [31:0] n39328;
wire     [31:0] n39329;
wire     [31:0] n39330;
wire     [31:0] n39331;
wire     [31:0] n39332;
wire     [31:0] n39333;
wire     [31:0] n39334;
wire     [31:0] n39335;
wire     [31:0] n39336;
wire     [31:0] n39337;
wire     [31:0] n39338;
wire     [31:0] n39339;
wire     [31:0] n39340;
wire     [31:0] n39341;
wire     [31:0] n39342;
wire     [31:0] n39343;
wire     [31:0] n39344;
wire     [31:0] n39345;
wire     [31:0] n39346;
wire     [31:0] n39347;
wire     [31:0] n39348;
wire     [31:0] n39349;
wire     [31:0] n39350;
wire     [31:0] n39351;
wire     [31:0] n39352;
wire     [31:0] n39353;
wire     [31:0] n39354;
wire     [31:0] n39355;
wire     [31:0] n39356;
wire     [31:0] n39357;
wire     [31:0] n39358;
wire     [31:0] n39359;
wire     [31:0] n39360;
wire     [31:0] n39361;
wire     [31:0] n39362;
wire     [31:0] n39363;
wire     [31:0] n39364;
wire     [31:0] n39365;
wire     [31:0] n39366;
wire     [31:0] n39367;
wire     [31:0] n39368;
wire     [31:0] n39369;
wire     [31:0] n39370;
wire     [31:0] n39371;
wire     [31:0] n39372;
wire     [31:0] n39373;
wire     [31:0] n39374;
wire     [31:0] n39375;
wire     [31:0] n39376;
wire     [31:0] n39377;
wire     [31:0] n39378;
wire     [31:0] n39379;
wire     [31:0] n39380;
wire     [31:0] n39381;
wire     [31:0] n39382;
wire     [31:0] n39383;
wire     [31:0] n39384;
wire     [31:0] n39385;
wire     [31:0] n39386;
wire     [31:0] n39387;
wire     [31:0] n39388;
wire     [31:0] n39389;
wire     [31:0] n39390;
wire     [31:0] n39391;
wire     [31:0] n39392;
wire     [31:0] n39393;
wire     [31:0] n39394;
wire     [31:0] n39395;
wire     [31:0] n39396;
wire     [31:0] n39397;
wire     [31:0] n39398;
wire     [31:0] n39399;
wire     [31:0] n39400;
wire     [31:0] n39401;
wire     [31:0] n39402;
wire     [31:0] n39403;
wire     [31:0] n39404;
wire     [31:0] n39405;
wire     [31:0] n39406;
wire     [31:0] n39407;
wire     [31:0] n39408;
wire     [31:0] n39409;
wire     [31:0] n39410;
wire     [31:0] n39411;
wire     [31:0] n39412;
wire     [31:0] n39413;
wire     [31:0] n39414;
wire     [31:0] n39415;
wire     [31:0] n39416;
wire     [31:0] n39417;
wire     [31:0] n39418;
wire     [31:0] n39419;
wire     [31:0] n39420;
wire     [31:0] n39421;
wire     [31:0] n39422;
wire     [31:0] n39423;
wire     [31:0] n39424;
wire     [31:0] n39425;
wire     [31:0] n39426;
wire     [31:0] n39427;
wire     [31:0] n39428;
wire     [31:0] n39429;
wire     [31:0] n39430;
wire     [31:0] n39431;
wire     [31:0] n39432;
wire     [31:0] n39433;
wire     [31:0] n39434;
wire     [31:0] n39435;
wire     [31:0] n39436;
wire     [31:0] n39437;
wire     [31:0] n39438;
wire     [31:0] n39439;
wire     [31:0] n39440;
wire     [31:0] n39441;
wire     [31:0] n39442;
wire     [31:0] n39443;
wire     [31:0] n39444;
wire     [31:0] n39445;
wire     [31:0] n39446;
wire     [31:0] n39447;
wire     [31:0] n39448;
wire     [31:0] n39449;
wire     [31:0] n39450;
wire     [31:0] n39451;
wire     [31:0] n39452;
wire     [31:0] n39453;
wire     [31:0] n39454;
wire     [31:0] n39455;
wire     [31:0] n39456;
wire     [31:0] n39457;
wire     [31:0] n39458;
wire     [31:0] n39459;
wire     [31:0] n39460;
wire     [31:0] n39461;
wire     [31:0] n39462;
wire     [31:0] n39463;
wire     [31:0] n39464;
wire     [31:0] n39465;
wire     [31:0] n39466;
wire     [31:0] n39467;
wire     [31:0] n39468;
wire     [31:0] n39469;
wire     [31:0] n39470;
wire     [31:0] n39471;
wire     [31:0] n39472;
wire     [31:0] n39473;
wire     [31:0] n39474;
wire     [31:0] n39475;
wire     [31:0] n39476;
wire     [31:0] n39477;
wire     [31:0] n39478;
wire     [31:0] n39479;
wire     [31:0] n39480;
wire     [31:0] n39481;
wire     [31:0] n39482;
wire     [31:0] n39483;
wire     [31:0] n39484;
wire     [31:0] n39485;
wire     [31:0] n39486;
wire     [31:0] n39487;
wire     [31:0] n39488;
wire     [31:0] n39489;
wire     [31:0] n39490;
wire     [31:0] n39491;
wire     [31:0] n39492;
wire     [31:0] n39493;
wire     [31:0] n39494;
wire     [31:0] n39495;
wire     [31:0] n39496;
wire     [31:0] n39497;
wire     [31:0] n39498;
wire     [31:0] n39499;
wire     [31:0] n39500;
wire     [31:0] n39501;
wire     [31:0] n39502;
wire     [31:0] n39503;
wire     [31:0] n39504;
wire     [31:0] n39505;
wire     [31:0] n39506;
wire     [31:0] n39507;
wire     [31:0] n39508;
wire     [31:0] n39509;
wire     [31:0] n39510;
wire     [31:0] n39511;
wire     [31:0] n39512;
wire     [31:0] n39513;
wire     [31:0] n39514;
wire     [31:0] n39515;
wire     [31:0] n39516;
wire     [31:0] n39517;
wire     [31:0] n39518;
wire     [31:0] n39519;
wire     [31:0] n39520;
wire     [31:0] n39521;
wire     [31:0] n39522;
wire     [31:0] n39523;
wire     [31:0] n39524;
wire     [31:0] n39525;
wire     [31:0] n39526;
wire     [31:0] n39527;
wire     [31:0] n39528;
wire     [31:0] n39529;
wire     [31:0] n39530;
wire     [31:0] n39531;
wire     [31:0] n39532;
wire     [31:0] n39533;
wire     [31:0] n39534;
wire     [31:0] n39535;
wire     [31:0] n39536;
wire     [31:0] n39537;
wire     [31:0] n39538;
wire     [31:0] n39539;
wire     [31:0] n39540;
wire     [31:0] n39541;
wire     [31:0] n39542;
wire     [31:0] n39543;
wire     [31:0] n39544;
wire     [31:0] n39545;
wire     [31:0] n39546;
wire     [31:0] n39547;
wire     [31:0] n39548;
wire     [31:0] n39549;
wire     [31:0] n39550;
wire     [31:0] n39551;
wire     [31:0] n39552;
wire     [31:0] n39553;
wire     [31:0] n39554;
wire     [31:0] n39555;
wire     [31:0] n39556;
wire     [31:0] n39557;
wire     [31:0] n39558;
wire     [31:0] n39559;
wire     [31:0] n39560;
wire     [31:0] n39561;
wire     [31:0] n39562;
wire     [31:0] n39563;
wire     [31:0] n39564;
wire     [31:0] n39565;
wire     [31:0] n39566;
wire     [31:0] n39567;
wire     [31:0] n39568;
wire     [31:0] n39569;
wire     [31:0] n39570;
wire     [31:0] n39571;
wire     [31:0] n39572;
wire     [31:0] n39573;
wire     [31:0] n39574;
wire     [31:0] n39575;
wire     [31:0] n39576;
wire     [31:0] n39577;
wire     [31:0] n39578;
wire     [31:0] n39579;
wire     [31:0] n39580;
wire     [31:0] n39581;
wire     [31:0] n39582;
wire     [31:0] n39583;
wire     [31:0] n39584;
wire     [31:0] n39585;
wire     [31:0] n39586;
wire     [31:0] n39587;
wire     [31:0] n39588;
wire     [31:0] n39589;
wire     [31:0] n39590;
wire     [31:0] n39591;
wire     [31:0] n39592;
wire     [31:0] n39593;
wire     [31:0] n39594;
wire     [31:0] n39595;
wire     [31:0] n39596;
wire     [31:0] n39597;
wire     [31:0] n39598;
wire     [31:0] n39599;
wire     [31:0] n39600;
wire     [31:0] n39601;
wire     [31:0] n39602;
wire     [31:0] n39603;
wire     [31:0] n39604;
wire     [31:0] n39605;
wire     [31:0] n39606;
wire     [31:0] n39607;
wire     [31:0] n39608;
wire     [31:0] n39609;
wire     [31:0] n39610;
wire     [31:0] n39611;
wire     [31:0] n39612;
wire     [31:0] n39613;
wire     [31:0] n39614;
wire     [31:0] n39615;
wire     [31:0] n39616;
wire     [31:0] n39617;
wire     [31:0] n39618;
wire     [31:0] n39619;
wire     [31:0] n39620;
wire     [31:0] n39621;
wire     [31:0] n39622;
wire     [31:0] n39623;
wire     [31:0] n39624;
wire     [31:0] n39625;
wire     [31:0] n39626;
wire     [31:0] n39627;
wire     [31:0] n39628;
wire     [31:0] n39629;
wire     [31:0] n39630;
wire     [31:0] n39631;
wire     [31:0] n39632;
wire     [31:0] n39633;
wire     [31:0] n39634;
wire     [31:0] n39635;
wire     [31:0] n39636;
wire     [31:0] n39637;
wire     [31:0] n39638;
wire     [31:0] n39639;
wire     [31:0] n39640;
wire     [31:0] n39641;
wire     [31:0] n39642;
wire     [31:0] n39643;
wire     [31:0] n39644;
wire     [31:0] n39645;
wire     [31:0] n39646;
wire     [31:0] n39647;
wire     [31:0] n39648;
wire     [31:0] n39649;
wire     [31:0] n39650;
wire     [31:0] n39651;
wire     [31:0] n39652;
wire     [31:0] n39653;
wire     [31:0] n39654;
wire     [31:0] n39655;
wire     [31:0] n39656;
wire     [31:0] n39657;
wire     [31:0] n39658;
wire     [31:0] n39659;
wire     [31:0] n39660;
wire     [31:0] n39661;
wire     [31:0] n39662;
wire     [31:0] n39663;
wire     [31:0] n39664;
wire     [31:0] n39665;
wire     [31:0] n39666;
wire     [31:0] n39667;
wire     [31:0] n39668;
wire     [31:0] n39669;
wire     [31:0] n39670;
wire     [31:0] n39671;
wire     [31:0] n39672;
wire     [31:0] n39673;
wire     [31:0] n39674;
wire     [31:0] n39675;
wire     [31:0] n39676;
wire     [31:0] n39677;
wire     [31:0] n39678;
wire     [31:0] n39679;
wire     [31:0] n39680;
wire     [31:0] n39681;
wire     [31:0] n39682;
wire     [31:0] n39683;
wire     [31:0] n39684;
wire     [31:0] n39685;
wire     [31:0] n39686;
wire     [31:0] n39687;
wire     [31:0] n39688;
wire     [31:0] n39689;
wire     [31:0] n39690;
wire     [31:0] n39691;
wire     [31:0] n39692;
wire     [31:0] n39693;
wire     [31:0] n39694;
wire     [31:0] n39695;
wire     [31:0] n39696;
wire     [31:0] n39697;
wire     [31:0] n39698;
wire     [31:0] n39699;
wire     [31:0] n39700;
wire     [31:0] n39701;
wire     [31:0] n39702;
wire     [31:0] n39703;
wire     [31:0] n39704;
wire     [31:0] n39705;
wire     [31:0] n39706;
wire     [31:0] n39707;
wire     [31:0] n39708;
wire     [31:0] n39709;
wire     [31:0] n39710;
wire     [31:0] n39711;
wire     [31:0] n39712;
wire     [31:0] n39713;
wire     [31:0] n39714;
wire     [31:0] n39715;
wire     [31:0] n39716;
wire     [31:0] n39717;
wire     [31:0] n39718;
wire     [31:0] n39719;
wire     [31:0] n39720;
wire     [31:0] n39721;
wire     [31:0] n39722;
wire     [31:0] n39723;
wire     [31:0] n39724;
wire     [31:0] n39725;
wire     [31:0] n39726;
wire     [31:0] n39727;
wire     [31:0] n39728;
wire     [31:0] n39729;
wire     [31:0] n39730;
wire     [31:0] n39731;
wire     [31:0] n39732;
wire     [31:0] n39733;
wire     [31:0] n39734;
wire     [31:0] n39735;
wire     [31:0] n39736;
wire     [31:0] n39737;
wire     [31:0] n39738;
wire     [31:0] n39739;
wire     [31:0] n39740;
wire     [31:0] n39741;
wire     [31:0] n39742;
wire     [31:0] n39743;
wire     [31:0] n39744;
wire     [31:0] n39745;
wire     [31:0] n39746;
wire     [31:0] n39747;
wire     [31:0] n39748;
wire     [31:0] n39749;
wire     [31:0] n39750;
wire     [31:0] n39751;
wire     [31:0] n39752;
wire     [31:0] n39753;
wire     [31:0] n39754;
wire     [31:0] n39755;
wire     [31:0] n39756;
wire     [31:0] n39757;
wire     [31:0] n39758;
wire     [31:0] n39759;
wire     [31:0] n39760;
wire     [31:0] n39761;
wire     [31:0] n39762;
wire     [31:0] n39763;
wire     [31:0] n39764;
wire     [31:0] n39765;
wire     [31:0] n39766;
wire     [31:0] n39767;
wire     [31:0] n39768;
wire     [31:0] n39769;
wire     [31:0] n39770;
wire     [31:0] n39771;
wire     [31:0] n39772;
wire     [31:0] n39773;
wire     [31:0] n39774;
wire     [31:0] n39775;
wire     [31:0] n39776;
wire     [31:0] n39777;
wire     [31:0] n39778;
wire     [31:0] n39779;
wire     [31:0] n39780;
wire     [31:0] n39781;
wire     [31:0] n39782;
wire     [31:0] n39783;
wire     [31:0] n39784;
wire     [31:0] n39785;
wire     [31:0] n39786;
wire     [31:0] n39787;
wire     [31:0] n39788;
wire     [31:0] n39789;
wire     [31:0] n39790;
wire     [31:0] n39791;
wire     [31:0] n39792;
wire     [31:0] n39793;
wire     [31:0] n39794;
wire     [31:0] n39795;
wire     [31:0] n39796;
wire     [31:0] n39797;
wire     [31:0] n39798;
wire     [31:0] n39799;
wire     [31:0] n39800;
wire     [31:0] n39801;
wire     [31:0] n39802;
wire     [31:0] n39803;
wire     [31:0] n39804;
wire     [31:0] n39805;
wire     [31:0] n39806;
wire     [31:0] n39807;
wire     [31:0] n39808;
wire     [31:0] n39809;
wire     [31:0] n39810;
wire     [31:0] n39811;
wire     [31:0] n39812;
wire     [31:0] n39813;
wire     [31:0] n39814;
wire     [31:0] n39815;
wire     [31:0] n39816;
wire     [31:0] n39817;
wire     [31:0] n39818;
wire     [31:0] n39819;
wire     [31:0] n39820;
wire     [31:0] n39821;
wire     [31:0] n39822;
wire     [31:0] n39823;
wire     [31:0] n39824;
wire     [31:0] n39825;
wire     [31:0] n39826;
wire     [31:0] n39827;
wire     [31:0] n39828;
wire     [31:0] n39829;
wire     [31:0] n39830;
wire     [31:0] n39831;
wire     [31:0] n39832;
wire     [31:0] n39833;
wire     [31:0] n39834;
wire     [31:0] n39835;
wire     [31:0] n39836;
wire     [31:0] n39837;
wire     [31:0] n39838;
wire     [31:0] n39839;
wire     [31:0] n39840;
wire     [31:0] n39841;
wire     [31:0] n39842;
wire     [31:0] n39843;
wire     [31:0] n39844;
wire     [31:0] n39845;
wire     [31:0] n39846;
wire     [31:0] n39847;
wire     [31:0] n39848;
wire     [31:0] n39849;
wire     [31:0] n39850;
wire     [31:0] n39851;
wire     [31:0] n39852;
wire     [31:0] n39853;
wire     [31:0] n39854;
wire     [31:0] n39855;
wire     [31:0] n39856;
wire     [31:0] n39857;
wire     [31:0] n39858;
wire     [31:0] n39859;
wire     [31:0] n39860;
wire     [31:0] n39861;
wire     [31:0] n39862;
wire     [31:0] n39863;
wire     [31:0] n39864;
wire     [31:0] n39865;
wire     [31:0] n39866;
wire     [31:0] n39867;
wire     [31:0] n39868;
wire     [31:0] n39869;
wire     [31:0] n39870;
wire     [31:0] n39871;
wire     [31:0] n39872;
wire     [31:0] n39873;
wire     [31:0] n39874;
wire     [31:0] n39875;
wire     [31:0] n39876;
wire     [31:0] n39877;
wire     [31:0] n39878;
wire     [31:0] n39879;
wire     [31:0] n39880;
wire     [31:0] n39881;
wire     [31:0] n39882;
wire     [31:0] n39883;
wire     [31:0] n39884;
wire     [31:0] n39885;
wire     [31:0] n39886;
wire     [31:0] n39887;
wire     [31:0] n39888;
wire     [31:0] n39889;
wire     [31:0] n39890;
wire     [31:0] n39891;
wire     [31:0] n39892;
wire     [31:0] n39893;
wire     [31:0] n39894;
wire     [31:0] n39895;
wire     [31:0] n39896;
wire     [31:0] n39897;
wire     [31:0] n39898;
wire     [31:0] n39899;
wire     [31:0] n39900;
wire     [31:0] n39901;
wire     [31:0] n39902;
wire     [31:0] n39903;
wire     [31:0] n39904;
wire     [31:0] n39905;
wire     [31:0] n39906;
wire     [31:0] n39907;
wire     [31:0] n39908;
wire     [31:0] n39909;
wire     [31:0] n39910;
wire     [31:0] n39911;
wire     [31:0] n39912;
wire     [31:0] n39913;
wire     [31:0] n39914;
wire     [31:0] n39915;
wire     [31:0] n39916;
wire     [31:0] n39917;
wire     [31:0] n39918;
wire     [31:0] n39919;
wire     [31:0] n39920;
wire     [31:0] n39921;
wire     [31:0] n39922;
wire     [31:0] n39923;
wire     [31:0] n39924;
wire     [31:0] n39925;
wire     [31:0] n39926;
wire     [31:0] n39927;
wire     [31:0] n39928;
wire     [31:0] n39929;
wire     [31:0] n39930;
wire     [31:0] n39931;
wire     [31:0] n39932;
wire     [31:0] n39933;
wire     [31:0] n39934;
wire     [31:0] n39935;
wire     [31:0] n39936;
wire     [31:0] n39937;
wire     [31:0] n39938;
wire     [31:0] n39939;
wire     [31:0] n39940;
wire     [31:0] n39941;
wire     [31:0] n39942;
wire     [31:0] n39943;
wire     [31:0] n39944;
wire     [31:0] n39945;
wire     [31:0] n39946;
wire     [31:0] n39947;
wire     [31:0] n39948;
wire     [31:0] n39949;
wire     [31:0] n39950;
wire     [31:0] n39951;
wire     [31:0] n39952;
wire     [31:0] n39953;
wire     [31:0] n39954;
wire     [31:0] n39955;
wire     [31:0] n39956;
wire     [31:0] n39957;
wire     [31:0] n39958;
wire     [31:0] n39959;
wire     [31:0] n39960;
wire     [31:0] n39961;
wire     [31:0] n39962;
wire     [31:0] n39963;
wire     [31:0] n39964;
wire     [31:0] n39965;
wire     [31:0] n39966;
wire     [31:0] n39967;
wire     [31:0] n39968;
wire     [31:0] n39969;
wire     [31:0] n39970;
wire     [31:0] n39971;
wire     [31:0] n39972;
wire     [31:0] n39973;
wire     [31:0] n39974;
wire     [31:0] n39975;
wire     [31:0] n39976;
wire     [31:0] n39977;
wire     [31:0] n39978;
wire     [31:0] n39979;
wire     [31:0] n39980;
wire     [31:0] n39981;
wire     [31:0] n39982;
wire     [31:0] n39983;
wire     [31:0] n39984;
wire     [31:0] n39985;
wire     [31:0] n39986;
wire     [31:0] n39987;
wire     [31:0] n39988;
wire     [31:0] n39989;
wire     [31:0] n39990;
wire     [31:0] n39991;
wire     [31:0] n39992;
wire     [31:0] n39993;
wire     [31:0] n39994;
wire     [31:0] n39995;
wire     [31:0] n39996;
wire     [31:0] n39997;
wire     [31:0] n39998;
wire     [31:0] n39999;
wire     [31:0] n40000;
wire     [31:0] n40001;
wire     [31:0] n40002;
wire     [31:0] n40003;
wire     [31:0] n40004;
wire     [31:0] n40005;
wire     [31:0] n40006;
wire     [31:0] n40007;
wire     [31:0] n40008;
wire     [31:0] n40009;
wire     [31:0] n40010;
wire     [31:0] n40011;
wire     [31:0] n40012;
wire     [31:0] n40013;
wire     [31:0] n40014;
wire     [31:0] n40015;
wire     [31:0] n40016;
wire     [31:0] n40017;
wire     [31:0] n40018;
wire     [31:0] n40019;
wire     [31:0] n40020;
wire     [31:0] n40021;
wire     [31:0] n40022;
wire     [31:0] n40023;
wire     [31:0] n40024;
wire     [31:0] n40025;
wire     [31:0] n40026;
wire     [31:0] n40027;
wire     [31:0] n40028;
wire     [31:0] n40029;
wire     [31:0] n40030;
wire     [31:0] n40031;
wire     [31:0] n40032;
wire     [31:0] n40033;
wire     [31:0] n40034;
wire     [31:0] n40035;
wire     [31:0] n40036;
wire     [31:0] n40037;
wire     [31:0] n40038;
wire     [31:0] n40039;
wire     [31:0] n40040;
wire     [31:0] n40041;
wire     [31:0] n40042;
wire     [31:0] n40043;
wire     [31:0] n40044;
wire     [31:0] n40045;
wire     [31:0] n40046;
wire     [31:0] n40047;
wire     [31:0] n40048;
wire     [31:0] n40049;
wire     [31:0] n40050;
wire     [31:0] n40051;
wire     [31:0] n40052;
wire     [31:0] n40053;
wire     [31:0] n40054;
wire     [31:0] n40055;
wire     [31:0] n40056;
wire     [31:0] n40057;
wire     [31:0] n40058;
wire     [31:0] n40059;
wire     [31:0] n40060;
wire     [31:0] n40061;
wire     [31:0] n40062;
wire     [31:0] n40063;
wire     [31:0] n40064;
wire     [31:0] n40065;
wire     [31:0] n40066;
wire     [31:0] n40067;
wire     [31:0] n40068;
wire     [31:0] n40069;
wire     [31:0] n40070;
wire     [31:0] n40071;
wire     [31:0] n40072;
wire     [31:0] n40073;
wire     [31:0] n40074;
wire     [31:0] n40075;
wire     [31:0] n40076;
wire     [31:0] n40077;
wire     [31:0] n40078;
wire     [31:0] n40079;
wire     [31:0] n40080;
wire     [31:0] n40081;
wire     [31:0] n40082;
wire     [31:0] n40083;
wire     [31:0] n40084;
wire     [31:0] n40085;
wire     [31:0] n40086;
wire     [31:0] n40087;
wire     [31:0] n40088;
wire     [31:0] n40089;
wire     [31:0] n40090;
wire     [31:0] n40091;
wire     [31:0] n40092;
wire     [31:0] n40093;
wire     [31:0] n40094;
wire     [31:0] n40095;
wire     [31:0] n40096;
wire     [31:0] n40097;
wire     [31:0] n40098;
wire     [31:0] n40099;
wire     [31:0] n40100;
wire     [31:0] n40101;
wire     [31:0] n40102;
wire     [31:0] n40103;
wire     [31:0] n40104;
wire     [31:0] n40105;
wire     [31:0] n40106;
wire     [31:0] n40107;
wire     [31:0] n40108;
wire     [31:0] n40109;
wire     [31:0] n40110;
wire     [31:0] n40111;
wire     [31:0] n40112;
wire     [31:0] n40113;
wire     [31:0] n40114;
wire     [31:0] n40115;
wire     [31:0] n40116;
wire     [31:0] n40117;
wire     [31:0] n40118;
wire     [31:0] n40119;
wire     [31:0] n40120;
wire     [31:0] n40121;
wire     [31:0] n40122;
wire     [31:0] n40123;
wire     [31:0] n40124;
wire     [31:0] n40125;
wire     [31:0] n40126;
wire     [31:0] n40127;
wire     [31:0] n40128;
wire     [31:0] n40129;
wire     [31:0] n40130;
wire     [31:0] n40131;
wire     [31:0] n40132;
wire     [31:0] n40133;
wire     [31:0] n40134;
wire     [31:0] n40135;
wire     [31:0] n40136;
wire     [31:0] n40137;
wire     [31:0] n40138;
wire     [31:0] n40139;
wire     [31:0] n40140;
wire     [31:0] n40141;
wire     [31:0] n40142;
wire     [31:0] n40143;
wire     [31:0] n40144;
wire     [31:0] n40145;
wire     [31:0] n40146;
wire     [31:0] n40147;
wire     [31:0] n40148;
wire     [31:0] n40149;
wire     [31:0] n40150;
wire     [31:0] n40151;
wire     [31:0] n40152;
wire     [31:0] n40153;
wire     [31:0] n40154;
wire     [31:0] n40155;
wire     [31:0] n40156;
wire     [31:0] n40157;
wire     [31:0] n40158;
wire     [31:0] n40159;
wire     [31:0] n40160;
wire     [31:0] n40161;
wire     [31:0] n40162;
wire     [31:0] n40163;
wire     [31:0] n40164;
wire     [31:0] n40165;
wire     [31:0] n40166;
wire     [31:0] n40167;
wire     [31:0] n40168;
wire     [31:0] n40169;
wire     [31:0] n40170;
wire     [31:0] n40171;
wire     [31:0] n40172;
wire     [31:0] n40173;
wire     [31:0] n40174;
wire     [31:0] n40175;
wire     [31:0] n40176;
wire     [31:0] n40177;
wire     [31:0] n40178;
wire     [31:0] n40179;
wire     [31:0] n40180;
wire     [31:0] n40181;
wire     [31:0] n40182;
wire     [31:0] n40183;
wire     [31:0] n40184;
wire     [31:0] n40185;
wire     [31:0] n40186;
wire     [31:0] n40187;
wire     [31:0] n40188;
wire     [31:0] n40189;
wire     [31:0] n40190;
wire     [31:0] n40191;
wire     [31:0] n40192;
wire     [31:0] n40193;
wire     [31:0] n40194;
wire     [31:0] n40195;
wire     [31:0] n40196;
wire     [31:0] n40197;
wire     [31:0] n40198;
wire     [31:0] n40199;
wire     [31:0] n40200;
wire     [31:0] n40201;
wire     [31:0] n40202;
wire     [31:0] n40203;
wire     [31:0] n40204;
wire     [31:0] n40205;
wire     [31:0] n40206;
wire     [31:0] n40207;
wire     [31:0] n40208;
wire     [31:0] n40209;
wire     [31:0] n40210;
wire     [31:0] n40211;
wire     [31:0] n40212;
wire     [31:0] n40213;
wire     [31:0] n40214;
wire     [31:0] n40215;
wire     [31:0] n40216;
wire     [31:0] n40217;
wire     [31:0] n40218;
wire     [31:0] n40219;
wire     [31:0] n40220;
wire     [31:0] n40221;
wire     [31:0] n40222;
wire     [31:0] n40223;
wire     [31:0] n40224;
wire     [31:0] n40225;
wire     [31:0] n40226;
wire     [31:0] n40227;
wire     [31:0] n40228;
wire     [31:0] n40229;
wire     [31:0] n40230;
wire     [31:0] n40231;
wire     [31:0] n40232;
wire     [31:0] n40233;
wire     [31:0] n40234;
wire     [31:0] n40235;
wire     [31:0] n40236;
wire     [31:0] n40237;
wire     [31:0] n40238;
wire     [31:0] n40239;
wire     [31:0] n40240;
wire     [31:0] n40241;
wire     [31:0] n40242;
wire     [31:0] n40243;
wire     [31:0] n40244;
wire     [31:0] n40245;
wire     [31:0] n40246;
wire     [31:0] n40247;
wire     [31:0] n40248;
wire     [31:0] n40249;
wire     [31:0] n40250;
wire     [31:0] n40251;
wire     [31:0] n40252;
wire     [31:0] n40253;
wire     [31:0] n40254;
wire     [31:0] n40255;
wire     [31:0] n40256;
wire     [31:0] n40257;
wire     [31:0] n40258;
wire     [31:0] n40259;
wire     [31:0] n40260;
wire     [31:0] n40261;
wire     [31:0] n40262;
wire     [31:0] n40263;
wire     [31:0] n40264;
wire     [31:0] n40265;
wire     [31:0] n40266;
wire     [31:0] n40267;
wire     [31:0] n40268;
wire     [31:0] n40269;
wire     [31:0] n40270;
wire     [31:0] n40271;
wire     [31:0] n40272;
wire     [31:0] n40273;
wire     [31:0] n40274;
wire     [31:0] n40275;
wire     [31:0] n40276;
wire     [31:0] n40277;
wire     [31:0] n40278;
wire     [31:0] n40279;
wire     [31:0] n40280;
wire     [31:0] n40281;
wire     [31:0] n40282;
wire     [31:0] n40283;
wire     [31:0] n40284;
wire     [31:0] n40285;
wire     [31:0] n40286;
wire     [31:0] n40287;
wire     [31:0] n40288;
wire     [31:0] n40289;
wire     [31:0] n40290;
wire     [31:0] n40291;
wire     [31:0] n40292;
wire     [31:0] n40293;
wire     [31:0] n40294;
wire     [31:0] n40295;
wire     [31:0] n40296;
wire     [31:0] n40297;
wire     [31:0] n40298;
wire     [31:0] n40299;
wire     [31:0] n40300;
wire     [31:0] n40301;
wire     [31:0] n40302;
wire     [31:0] n40303;
wire     [31:0] n40304;
wire     [31:0] n40305;
wire     [31:0] n40306;
wire     [31:0] n40307;
wire     [31:0] n40308;
wire     [31:0] n40309;
wire     [31:0] n40310;
wire     [31:0] n40311;
wire     [31:0] n40312;
wire     [31:0] n40313;
wire     [31:0] n40314;
wire     [31:0] n40315;
wire     [31:0] n40316;
wire     [31:0] n40317;
wire     [31:0] n40318;
wire     [31:0] n40319;
wire     [31:0] n40320;
wire     [31:0] n40321;
wire     [31:0] n40322;
wire     [31:0] n40323;
wire     [31:0] n40324;
wire     [31:0] n40325;
wire     [31:0] n40326;
wire     [31:0] n40327;
wire     [31:0] n40328;
wire     [31:0] n40329;
wire     [31:0] n40330;
wire     [31:0] n40331;
wire     [31:0] n40332;
wire     [31:0] n40333;
wire     [31:0] n40334;
wire     [31:0] n40335;
wire     [31:0] n40336;
wire     [31:0] n40337;
wire     [31:0] n40338;
wire     [31:0] n40339;
wire     [31:0] n40340;
wire     [31:0] n40341;
wire     [31:0] n40342;
wire     [31:0] n40343;
wire     [31:0] n40344;
wire     [31:0] n40345;
wire     [31:0] n40346;
wire     [31:0] n40347;
wire     [31:0] n40348;
wire     [31:0] n40349;
wire     [31:0] n40350;
wire     [31:0] n40351;
wire     [31:0] n40352;
wire     [31:0] n40353;
wire     [31:0] n40354;
wire     [31:0] n40355;
wire     [31:0] n40356;
wire     [31:0] n40357;
wire     [31:0] n40358;
wire     [31:0] n40359;
wire     [31:0] n40360;
wire     [31:0] n40361;
wire     [31:0] n40362;
wire     [31:0] n40363;
wire     [31:0] n40364;
wire     [31:0] n40365;
wire     [31:0] n40366;
wire     [31:0] n40367;
wire     [31:0] n40368;
wire     [31:0] n40369;
wire     [31:0] n40370;
wire     [31:0] n40371;
wire     [31:0] n40372;
wire     [31:0] n40373;
wire     [31:0] n40374;
wire     [31:0] n40375;
wire     [31:0] n40376;
wire     [31:0] n40377;
wire     [31:0] n40378;
wire     [31:0] n40379;
wire     [31:0] n40380;
wire     [31:0] n40381;
wire     [31:0] n40382;
wire     [31:0] n40383;
wire     [31:0] n40384;
wire     [31:0] n40385;
wire     [31:0] n40386;
wire     [31:0] n40387;
wire     [31:0] n40388;
wire     [31:0] n40389;
wire     [31:0] n40390;
wire     [31:0] n40391;
wire     [31:0] n40392;
wire     [31:0] n40393;
wire     [31:0] n40394;
wire     [31:0] n40395;
wire     [31:0] n40396;
wire     [31:0] n40397;
wire     [31:0] n40398;
wire     [31:0] n40399;
wire     [31:0] n40400;
wire     [31:0] n40401;
wire     [31:0] n40402;
wire     [31:0] n40403;
wire     [31:0] n40404;
wire     [31:0] n40405;
wire     [31:0] n40406;
wire     [31:0] n40407;
wire     [31:0] n40408;
wire     [31:0] n40409;
wire     [31:0] n40410;
wire     [31:0] n40411;
wire     [31:0] n40412;
wire     [31:0] n40413;
wire     [31:0] n40414;
wire     [31:0] n40415;
wire     [31:0] n40416;
wire     [31:0] n40417;
wire     [31:0] n40418;
wire     [31:0] n40419;
wire     [31:0] n40420;
wire     [31:0] n40421;
wire     [31:0] n40422;
wire     [31:0] n40423;
wire     [31:0] n40424;
wire     [31:0] n40425;
wire     [31:0] n40426;
wire     [31:0] n40427;
wire     [31:0] n40428;
wire     [31:0] n40429;
wire     [31:0] n40430;
wire     [31:0] n40431;
wire     [31:0] n40432;
wire     [31:0] n40433;
wire     [31:0] n40434;
wire     [31:0] n40435;
wire     [31:0] n40436;
wire     [31:0] n40437;
wire     [31:0] n40438;
wire     [31:0] n40439;
wire     [31:0] n40440;
wire     [31:0] n40441;
wire     [31:0] n40442;
wire     [31:0] n40443;
wire     [31:0] n40444;
wire     [31:0] n40445;
wire     [31:0] n40446;
wire     [31:0] n40447;
wire     [31:0] n40448;
wire     [31:0] n40449;
wire     [31:0] n40450;
wire     [31:0] n40451;
wire     [31:0] n40452;
wire     [31:0] n40453;
wire     [31:0] n40454;
wire     [31:0] n40455;
wire     [31:0] n40456;
wire     [31:0] n40457;
wire     [31:0] n40458;
wire     [31:0] n40459;
wire     [31:0] n40460;
wire     [31:0] n40461;
wire     [31:0] n40462;
wire     [31:0] n40463;
wire     [31:0] n40464;
wire     [31:0] n40465;
wire     [31:0] n40466;
wire     [31:0] n40467;
wire     [31:0] n40468;
wire     [31:0] n40469;
wire     [31:0] n40470;
wire     [31:0] n40471;
wire     [31:0] n40472;
wire     [31:0] n40473;
wire     [31:0] n40474;
wire     [31:0] n40475;
wire     [31:0] n40476;
wire     [31:0] n40477;
wire     [31:0] n40478;
wire     [31:0] n40479;
wire     [31:0] n40480;
wire     [31:0] n40481;
wire     [31:0] n40482;
wire     [31:0] n40483;
wire     [31:0] n40484;
wire     [31:0] n40485;
wire     [31:0] n40486;
wire     [31:0] n40487;
wire     [31:0] n40488;
wire     [31:0] n40489;
wire     [31:0] n40490;
wire     [31:0] n40491;
wire     [31:0] n40492;
wire     [31:0] n40493;
wire     [31:0] n40494;
wire     [31:0] n40495;
wire     [31:0] n40496;
wire     [31:0] n40497;
wire     [31:0] n40498;
wire     [31:0] n40499;
wire     [31:0] n40500;
wire     [31:0] n40501;
wire     [31:0] n40502;
wire     [31:0] n40503;
wire     [31:0] n40504;
wire     [31:0] n40505;
wire     [31:0] n40506;
wire     [31:0] n40507;
wire     [31:0] n40508;
wire     [31:0] n40509;
wire     [31:0] n40510;
wire     [31:0] n40511;
wire     [31:0] n40512;
wire     [31:0] n40513;
wire     [31:0] n40514;
wire     [31:0] n40515;
wire     [31:0] n40516;
wire     [31:0] n40517;
wire     [31:0] n40518;
wire     [31:0] n40519;
wire     [31:0] n40520;
wire     [31:0] n40521;
wire     [31:0] n40522;
wire     [31:0] n40523;
wire     [31:0] n40524;
wire     [31:0] n40525;
wire     [31:0] n40526;
wire     [31:0] n40527;
wire     [31:0] n40528;
wire     [31:0] n40529;
wire     [31:0] n40530;
wire     [31:0] n40531;
wire     [31:0] n40532;
wire     [31:0] n40533;
wire     [31:0] n40534;
wire     [31:0] n40535;
wire     [31:0] n40536;
wire     [31:0] n40537;
wire     [31:0] n40538;
wire     [31:0] n40539;
wire     [31:0] n40540;
wire     [31:0] n40541;
wire     [31:0] n40542;
wire     [31:0] n40543;
wire     [31:0] n40544;
wire     [31:0] n40545;
wire     [31:0] n40546;
wire     [31:0] n40547;
wire     [31:0] n40548;
wire     [31:0] n40549;
wire     [31:0] n40550;
wire     [31:0] n40551;
wire     [31:0] n40552;
wire     [31:0] n40553;
wire     [31:0] n40554;
wire     [31:0] n40555;
wire     [31:0] n40556;
wire     [31:0] n40557;
wire     [31:0] n40558;
wire     [31:0] n40559;
wire     [31:0] n40560;
wire     [31:0] n40561;
wire     [31:0] n40562;
wire     [31:0] n40563;
wire     [31:0] n40564;
wire     [31:0] n40565;
wire     [31:0] n40566;
wire     [31:0] n40567;
wire     [31:0] n40568;
wire     [31:0] n40569;
wire     [31:0] n40570;
wire     [31:0] n40571;
wire     [31:0] n40572;
wire     [31:0] n40573;
wire     [31:0] n40574;
wire     [31:0] n40575;
wire     [31:0] n40576;
wire     [31:0] n40577;
wire     [31:0] n40578;
wire     [31:0] n40579;
wire     [31:0] n40580;
wire     [31:0] n40581;
wire     [31:0] n40582;
wire     [31:0] n40583;
wire     [31:0] n40584;
wire     [31:0] n40585;
wire     [31:0] n40586;
wire     [31:0] n40587;
wire     [31:0] n40588;
wire     [31:0] n40589;
wire     [31:0] n40590;
wire     [31:0] n40591;
wire     [31:0] n40592;
wire     [31:0] n40593;
wire     [31:0] n40594;
wire     [31:0] n40595;
wire     [31:0] n40596;
wire     [31:0] n40597;
wire     [31:0] n40598;
wire     [31:0] n40599;
wire     [31:0] n40600;
wire     [31:0] n40601;
wire     [31:0] n40602;
wire     [31:0] n40603;
wire     [31:0] n40604;
wire     [31:0] n40605;
wire     [31:0] n40606;
wire     [31:0] n40607;
wire     [31:0] n40608;
wire     [31:0] n40609;
wire     [31:0] n40610;
wire     [31:0] n40611;
wire     [31:0] n40612;
wire     [31:0] n40613;
wire     [31:0] n40614;
wire     [31:0] n40615;
wire     [31:0] n40616;
wire     [31:0] n40617;
wire     [31:0] n40618;
wire     [31:0] n40619;
wire     [31:0] n40620;
wire     [31:0] n40621;
wire     [31:0] n40622;
wire     [31:0] n40623;
wire     [31:0] n40624;
wire     [31:0] n40625;
wire     [31:0] n40626;
wire     [31:0] n40627;
wire     [31:0] n40628;
wire     [31:0] n40629;
wire     [31:0] n40630;
wire     [31:0] n40631;
wire     [31:0] n40632;
wire     [31:0] n40633;
wire     [31:0] n40634;
wire     [31:0] n40635;
wire     [31:0] n40636;
wire     [31:0] n40637;
wire     [31:0] n40638;
wire     [31:0] n40639;
wire     [31:0] n40640;
wire     [31:0] n40641;
wire     [31:0] n40642;
wire     [31:0] n40643;
wire     [31:0] n40644;
wire     [31:0] n40645;
wire     [31:0] n40646;
wire     [31:0] n40647;
wire     [31:0] n40648;
wire     [31:0] n40649;
wire     [31:0] n40650;
wire     [31:0] n40651;
wire     [31:0] n40652;
wire     [31:0] n40653;
wire     [31:0] n40654;
wire     [31:0] n40655;
wire     [31:0] n40656;
wire     [31:0] n40657;
wire     [31:0] n40658;
wire     [31:0] n40659;
wire     [31:0] n40660;
wire     [31:0] n40661;
wire     [31:0] n40662;
wire     [31:0] n40663;
wire     [31:0] n40664;
wire     [31:0] n40665;
wire     [31:0] n40666;
wire     [31:0] n40667;
wire     [31:0] n40668;
wire     [31:0] n40669;
wire     [31:0] n40670;
wire     [31:0] n40671;
wire     [31:0] n40672;
wire     [31:0] n40673;
wire     [31:0] n40674;
wire     [31:0] n40675;
wire     [31:0] n40676;
wire     [31:0] n40677;
wire     [31:0] n40678;
wire     [31:0] n40679;
wire     [31:0] n40680;
wire     [31:0] n40681;
wire     [31:0] n40682;
wire     [31:0] n40683;
wire     [31:0] n40684;
wire     [31:0] n40685;
wire     [31:0] n40686;
wire     [31:0] n40687;
wire     [31:0] n40688;
wire     [31:0] n40689;
wire     [31:0] n40690;
wire     [31:0] n40691;
wire     [31:0] n40692;
wire     [31:0] n40693;
wire     [31:0] n40694;
wire     [31:0] n40695;
wire     [31:0] n40696;
wire     [31:0] n40697;
wire     [31:0] n40698;
wire     [31:0] n40699;
wire     [31:0] n40700;
wire     [31:0] n40701;
wire     [31:0] n40702;
wire     [31:0] n40703;
wire     [31:0] n40704;
wire     [31:0] n40705;
wire     [31:0] n40706;
wire     [31:0] n40707;
wire     [31:0] n40708;
wire     [31:0] n40709;
wire     [31:0] n40710;
wire     [31:0] n40711;
wire     [31:0] n40712;
wire     [31:0] n40713;
wire     [31:0] n40714;
wire     [31:0] n40715;
wire     [31:0] n40716;
wire     [31:0] n40717;
wire     [31:0] n40718;
wire     [31:0] n40719;
wire     [31:0] n40720;
wire     [31:0] n40721;
wire     [31:0] n40722;
wire     [31:0] n40723;
wire     [31:0] n40724;
wire     [31:0] n40725;
wire     [31:0] n40726;
wire     [31:0] n40727;
wire     [31:0] n40728;
wire     [31:0] n40729;
wire     [31:0] n40730;
wire     [31:0] n40731;
wire     [31:0] n40732;
wire     [31:0] n40733;
wire     [31:0] n40734;
wire     [31:0] n40735;
wire     [31:0] n40736;
wire     [31:0] n40737;
wire     [31:0] n40738;
wire     [31:0] n40739;
wire     [31:0] n40740;
wire     [31:0] n40741;
wire     [31:0] n40742;
wire     [31:0] n40743;
wire     [31:0] n40744;
wire     [31:0] n40745;
wire     [31:0] n40746;
wire     [31:0] n40747;
wire     [31:0] n40748;
wire     [31:0] n40749;
wire     [31:0] n40750;
wire     [31:0] n40751;
wire     [31:0] n40752;
wire     [31:0] n40753;
wire     [31:0] n40754;
wire     [31:0] n40755;
wire     [31:0] n40756;
wire     [31:0] n40757;
wire     [31:0] n40758;
wire     [31:0] n40759;
wire     [31:0] n40760;
wire     [31:0] n40761;
wire     [31:0] n40762;
wire     [31:0] n40763;
wire     [31:0] n40764;
wire     [31:0] n40765;
wire     [31:0] n40766;
wire     [31:0] n40767;
wire     [31:0] n40768;
wire     [31:0] n40769;
wire     [31:0] n40770;
wire     [31:0] n40771;
wire     [31:0] n40772;
wire     [31:0] n40773;
wire     [31:0] n40774;
wire     [31:0] n40775;
wire     [31:0] n40776;
wire     [31:0] n40777;
wire     [31:0] n40778;
wire     [31:0] n40779;
wire     [31:0] n40780;
wire     [31:0] n40781;
wire     [31:0] n40782;
wire     [31:0] n40783;
wire     [31:0] n40784;
wire     [31:0] n40785;
wire     [31:0] n40786;
wire     [31:0] n40787;
wire     [31:0] n40788;
wire     [31:0] n40789;
wire     [31:0] n40790;
wire     [31:0] n40791;
wire     [31:0] n40792;
wire     [31:0] n40793;
wire     [31:0] n40794;
wire     [31:0] n40795;
wire     [31:0] n40796;
wire     [31:0] n40797;
wire     [31:0] n40798;
wire     [31:0] n40799;
wire     [31:0] n40800;
wire     [31:0] n40801;
wire     [31:0] n40802;
wire     [31:0] n40803;
wire     [31:0] n40804;
wire     [31:0] n40805;
wire     [31:0] n40806;
wire     [31:0] n40807;
wire     [31:0] n40808;
wire     [31:0] n40809;
wire     [31:0] n40810;
wire     [31:0] n40811;
wire     [31:0] n40812;
wire     [31:0] n40813;
wire     [31:0] n40814;
wire     [31:0] n40815;
wire     [31:0] n40816;
wire     [31:0] n40817;
wire     [31:0] n40818;
wire     [31:0] n40819;
wire     [31:0] n40820;
wire     [31:0] n40821;
wire     [31:0] n40822;
wire     [31:0] n40823;
wire     [31:0] n40824;
wire     [31:0] n40825;
wire     [31:0] n40826;
wire     [31:0] n40827;
wire     [31:0] n40828;
wire     [31:0] n40829;
wire     [31:0] n40830;
wire     [31:0] n40831;
wire     [31:0] n40832;
wire     [31:0] n40833;
wire     [31:0] n40834;
wire     [31:0] n40835;
wire     [31:0] n40836;
wire     [31:0] n40837;
wire     [31:0] n40838;
wire     [31:0] n40839;
wire     [31:0] n40840;
wire     [31:0] n40841;
wire     [31:0] n40842;
wire     [31:0] n40843;
wire     [31:0] n40844;
wire     [31:0] n40845;
wire     [31:0] n40846;
wire     [31:0] n40847;
wire     [31:0] n40848;
wire     [31:0] n40849;
wire     [31:0] n40850;
wire     [31:0] n40851;
wire     [31:0] n40852;
wire     [31:0] n40853;
wire     [31:0] n40854;
wire     [31:0] n40855;
wire     [31:0] n40856;
wire     [31:0] n40857;
wire     [31:0] n40858;
wire     [31:0] n40859;
wire     [31:0] n40860;
wire     [31:0] n40861;
wire     [31:0] n40862;
wire     [31:0] n40863;
wire     [31:0] n40864;
wire     [31:0] n40865;
wire     [31:0] n40866;
wire     [31:0] n40867;
wire     [31:0] n40868;
wire     [31:0] n40869;
wire     [31:0] n40870;
wire     [31:0] n40871;
wire     [31:0] n40872;
wire     [31:0] n40873;
wire     [31:0] n40874;
wire     [31:0] n40875;
wire     [31:0] n40876;
wire     [31:0] n40877;
wire     [31:0] n40878;
wire     [31:0] n40879;
wire     [31:0] n40880;
wire     [31:0] n40881;
wire     [31:0] n40882;
wire     [31:0] n40883;
wire     [31:0] n40884;
wire     [31:0] n40885;
wire     [31:0] n40886;
wire     [31:0] n40887;
wire     [31:0] n40888;
wire     [31:0] n40889;
wire     [31:0] n40890;
wire     [31:0] n40891;
wire     [31:0] n40892;
wire     [31:0] n40893;
wire     [31:0] n40894;
wire     [31:0] n40895;
wire     [31:0] n40896;
wire     [31:0] n40897;
wire     [31:0] n40898;
wire     [31:0] n40899;
wire     [31:0] n40900;
wire     [31:0] n40901;
wire     [31:0] n40902;
wire     [31:0] n40903;
wire     [31:0] n40904;
wire     [31:0] n40905;
wire     [31:0] n40906;
wire     [31:0] n40907;
wire     [31:0] n40908;
wire     [31:0] n40909;
wire     [31:0] n40910;
wire     [31:0] n40911;
wire     [31:0] n40912;
wire     [31:0] n40913;
wire     [31:0] n40914;
wire     [31:0] n40915;
wire     [31:0] n40916;
wire     [31:0] n40917;
wire     [31:0] n40918;
wire     [31:0] n40919;
wire     [31:0] n40920;
wire     [31:0] n40921;
wire     [31:0] n40922;
wire     [31:0] n40923;
wire     [31:0] n40924;
wire     [31:0] n40925;
wire     [31:0] n40926;
wire     [31:0] n40927;
wire     [31:0] n40928;
wire     [31:0] n40929;
wire     [31:0] n40930;
wire     [31:0] n40931;
wire     [31:0] n40932;
wire     [31:0] n40933;
wire     [31:0] n40934;
wire     [31:0] n40935;
wire     [31:0] n40936;
wire     [31:0] n40937;
wire     [31:0] n40938;
wire     [31:0] n40939;
wire     [31:0] n40940;
wire     [31:0] n40941;
wire     [31:0] n40942;
wire     [31:0] n40943;
wire     [31:0] n40944;
wire     [31:0] n40945;
wire     [31:0] n40946;
wire     [31:0] n40947;
wire     [31:0] n40948;
wire     [31:0] n40949;
wire     [31:0] n40950;
wire     [31:0] n40951;
wire     [31:0] n40952;
wire     [31:0] n40953;
wire     [31:0] n40954;
wire     [31:0] n40955;
wire     [31:0] n40956;
wire     [31:0] n40957;
wire     [31:0] n40958;
wire     [31:0] n40959;
wire     [31:0] n40960;
wire     [31:0] n40961;
wire     [31:0] n40962;
wire     [31:0] n40963;
wire     [31:0] n40964;
wire     [31:0] n40965;
wire     [31:0] n40966;
wire     [31:0] n40967;
wire     [31:0] n40968;
wire     [31:0] n40969;
wire     [31:0] n40970;
wire     [31:0] n40971;
wire     [31:0] n40972;
wire     [31:0] n40973;
wire     [31:0] n40974;
wire     [31:0] n40975;
wire     [31:0] n40976;
wire     [31:0] n40977;
wire     [31:0] n40978;
wire     [31:0] n40979;
wire     [31:0] n40980;
wire     [31:0] n40981;
wire     [31:0] n40982;
wire     [31:0] n40983;
wire     [31:0] n40984;
wire     [31:0] n40985;
wire     [31:0] n40986;
wire     [31:0] n40987;
wire     [31:0] n40988;
wire     [31:0] n40989;
wire     [31:0] n40990;
wire     [31:0] n40991;
wire     [31:0] n40992;
wire     [31:0] n40993;
wire     [31:0] n40994;
wire     [31:0] n40995;
wire     [31:0] n40996;
wire     [31:0] n40997;
wire     [31:0] n40998;
wire     [31:0] n40999;
wire     [31:0] n41000;
wire     [31:0] n41001;
wire     [31:0] n41002;
wire     [31:0] n41003;
wire     [31:0] n41004;
wire     [31:0] n41005;
wire     [31:0] n41006;
wire     [31:0] n41007;
wire     [31:0] n41008;
wire     [31:0] n41009;
wire     [31:0] n41010;
wire     [31:0] n41011;
wire     [31:0] n41012;
wire     [31:0] n41013;
wire     [31:0] n41014;
wire     [31:0] n41015;
wire     [31:0] n41016;
wire     [31:0] n41017;
wire     [31:0] n41018;
wire     [31:0] n41019;
wire     [31:0] n41020;
wire     [31:0] n41021;
wire     [31:0] n41022;
wire     [31:0] n41023;
wire     [31:0] n41024;
wire     [31:0] n41025;
wire     [31:0] n41026;
wire     [31:0] n41027;
wire     [31:0] n41028;
wire     [31:0] n41029;
wire     [31:0] n41030;
wire     [31:0] n41031;
wire     [31:0] n41032;
wire     [31:0] n41033;
wire     [31:0] n41034;
wire     [31:0] n41035;
wire     [31:0] n41036;
wire     [31:0] n41037;
wire     [31:0] n41038;
wire     [31:0] n41039;
wire     [31:0] n41040;
wire     [31:0] n41041;
wire     [31:0] n41042;
wire     [31:0] n41043;
wire     [31:0] n41044;
wire     [31:0] n41045;
wire     [31:0] n41046;
wire     [31:0] n41047;
wire     [31:0] n41048;
wire     [31:0] n41049;
wire     [31:0] n41050;
wire     [31:0] n41051;
wire     [31:0] n41052;
wire     [31:0] n41053;
wire     [31:0] n41054;
wire     [31:0] n41055;
wire     [31:0] n41056;
wire     [31:0] n41057;
wire     [31:0] n41058;
wire     [31:0] n41059;
wire     [31:0] n41060;
wire     [31:0] n41061;
wire     [31:0] n41062;
wire     [31:0] n41063;
wire     [31:0] n41064;
wire     [31:0] n41065;
wire     [31:0] n41066;
wire     [31:0] n41067;
wire     [31:0] n41068;
wire     [31:0] n41069;
wire     [31:0] n41070;
wire     [31:0] n41071;
wire     [31:0] n41072;
wire     [31:0] n41073;
wire     [31:0] n41074;
wire     [31:0] n41075;
wire     [31:0] n41076;
wire     [31:0] n41077;
wire     [31:0] n41078;
wire     [31:0] n41079;
wire     [31:0] n41080;
wire     [31:0] n41081;
wire     [31:0] n41082;
wire     [31:0] n41083;
wire     [31:0] n41084;
wire     [31:0] n41085;
wire     [31:0] n41086;
wire     [31:0] n41087;
wire     [31:0] n41088;
wire     [31:0] n41089;
wire     [31:0] n41090;
wire     [31:0] n41091;
wire     [31:0] n41092;
wire     [31:0] n41093;
wire     [31:0] n41094;
wire     [31:0] n41095;
wire     [31:0] n41096;
wire     [31:0] n41097;
wire     [31:0] n41098;
wire     [31:0] n41099;
wire     [31:0] n41100;
wire     [31:0] n41101;
wire     [31:0] n41102;
wire     [31:0] n41103;
wire     [31:0] n41104;
wire     [31:0] n41105;
wire     [31:0] n41106;
wire     [31:0] n41107;
wire     [31:0] n41108;
wire     [31:0] n41109;
wire     [31:0] n41110;
wire     [31:0] n41111;
wire     [31:0] n41112;
wire     [31:0] n41113;
wire     [31:0] n41114;
wire     [31:0] n41115;
wire     [31:0] n41116;
wire     [31:0] n41117;
wire     [31:0] n41118;
wire     [31:0] n41119;
wire     [31:0] n41120;
wire     [31:0] n41121;
wire     [31:0] n41122;
wire     [31:0] n41123;
wire     [31:0] n41124;
wire     [31:0] n41125;
wire     [31:0] n41126;
wire     [31:0] n41127;
wire     [31:0] n41128;
wire     [31:0] n41129;
wire     [31:0] n41130;
wire     [31:0] n41131;
wire     [31:0] n41132;
wire     [31:0] n41133;
wire     [31:0] n41134;
wire     [31:0] n41135;
wire     [31:0] n41136;
wire     [31:0] n41137;
wire     [31:0] n41138;
wire     [31:0] n41139;
wire     [31:0] n41140;
wire     [31:0] n41141;
wire     [31:0] n41142;
wire     [31:0] n41143;
wire     [31:0] n41144;
wire     [31:0] n41145;
wire     [31:0] n41146;
wire     [31:0] n41147;
wire     [31:0] n41148;
wire     [31:0] n41149;
wire     [31:0] n41150;
wire     [31:0] n41151;
wire     [31:0] n41152;
wire     [31:0] n41153;
wire     [31:0] n41154;
wire     [31:0] n41155;
wire     [31:0] n41156;
wire     [31:0] n41157;
wire     [31:0] n41158;
wire     [31:0] n41159;
wire     [31:0] n41160;
wire     [31:0] n41161;
wire     [31:0] n41162;
wire     [31:0] n41163;
wire     [31:0] n41164;
wire     [31:0] n41165;
wire     [31:0] n41166;
wire     [31:0] n41167;
wire     [31:0] n41168;
wire     [31:0] n41169;
wire     [31:0] n41170;
wire     [31:0] n41171;
wire     [31:0] n41172;
wire     [31:0] n41173;
wire     [31:0] n41174;
wire     [31:0] n41175;
wire     [31:0] n41176;
wire     [31:0] n41177;
wire     [31:0] n41178;
wire     [31:0] n41179;
wire     [31:0] n41180;
wire     [31:0] n41181;
wire     [31:0] n41182;
wire     [31:0] n41183;
wire     [31:0] n41184;
wire     [31:0] n41185;
wire     [31:0] n41186;
wire     [31:0] n41187;
wire     [31:0] n41188;
wire     [31:0] n41189;
wire     [31:0] n41190;
wire     [31:0] n41191;
wire     [31:0] n41192;
wire     [31:0] n41193;
wire     [31:0] n41194;
wire     [31:0] n41195;
wire     [31:0] n41196;
wire     [31:0] n41197;
wire     [31:0] n41198;
wire     [31:0] n41199;
wire     [31:0] n41200;
wire     [31:0] n41201;
wire     [31:0] n41202;
wire     [31:0] n41203;
wire     [31:0] n41204;
wire     [31:0] n41205;
wire     [31:0] n41206;
wire     [31:0] n41207;
wire     [31:0] n41208;
wire     [31:0] n41209;
wire     [31:0] n41210;
wire     [31:0] n41211;
wire     [31:0] n41212;
wire     [31:0] n41213;
wire     [31:0] n41214;
wire     [31:0] n41215;
wire     [31:0] n41216;
wire     [31:0] n41217;
wire     [31:0] n41218;
wire     [31:0] n41219;
wire     [31:0] n41220;
wire     [31:0] n41221;
wire     [31:0] n41222;
wire     [31:0] n41223;
wire     [31:0] n41224;
wire     [31:0] n41225;
wire     [31:0] n41226;
wire     [31:0] n41227;
wire     [31:0] n41228;
wire     [31:0] n41229;
wire     [31:0] n41230;
wire     [31:0] n41231;
wire     [31:0] n41232;
wire     [31:0] n41233;
wire     [31:0] n41234;
wire     [31:0] n41235;
wire     [31:0] n41236;
wire     [31:0] n41237;
wire     [31:0] n41238;
wire     [31:0] n41239;
wire     [31:0] n41240;
wire     [31:0] n41241;
wire     [31:0] n41242;
wire     [31:0] n41243;
wire     [31:0] n41244;
wire     [31:0] n41245;
wire     [31:0] n41246;
wire     [31:0] n41247;
wire     [31:0] n41248;
wire     [31:0] n41249;
wire     [31:0] n41250;
wire     [31:0] n41251;
wire     [31:0] n41252;
wire     [31:0] n41253;
wire     [31:0] n41254;
wire     [31:0] n41255;
wire     [31:0] n41256;
wire     [31:0] n41257;
wire     [31:0] n41258;
wire     [31:0] n41259;
wire     [31:0] n41260;
wire     [31:0] n41261;
wire     [31:0] n41262;
wire     [31:0] n41263;
wire     [31:0] n41264;
wire     [31:0] n41265;
wire     [31:0] n41266;
wire     [31:0] n41267;
wire     [31:0] n41268;
wire     [31:0] n41269;
wire     [31:0] n41270;
wire     [31:0] n41271;
wire     [31:0] n41272;
wire     [31:0] n41273;
wire     [31:0] n41274;
wire     [31:0] n41275;
wire     [31:0] n41276;
wire     [31:0] n41277;
wire     [31:0] n41278;
wire     [31:0] n41279;
wire     [31:0] n41280;
wire     [31:0] n41281;
wire     [31:0] n41282;
wire     [31:0] n41283;
wire     [31:0] n41284;
wire     [31:0] n41285;
wire     [31:0] n41286;
wire     [31:0] n41287;
wire     [31:0] n41288;
wire     [31:0] n41289;
wire     [31:0] n41290;
wire     [31:0] n41291;
wire     [31:0] n41292;
wire     [31:0] n41293;
wire     [31:0] n41294;
wire     [31:0] n41295;
wire     [31:0] n41296;
wire     [31:0] n41297;
wire     [31:0] n41298;
wire     [31:0] n41299;
wire     [31:0] n41300;
wire     [31:0] n41301;
wire     [31:0] n41302;
wire     [31:0] n41303;
wire     [31:0] n41304;
wire     [31:0] n41305;
wire     [31:0] n41306;
wire     [31:0] n41307;
wire     [31:0] n41308;
wire     [31:0] n41309;
wire     [31:0] n41310;
wire     [31:0] n41311;
wire     [31:0] n41312;
wire     [31:0] n41313;
wire     [31:0] n41314;
wire     [31:0] n41315;
wire     [31:0] n41316;
wire     [31:0] n41317;
wire     [31:0] n41318;
wire     [31:0] n41319;
wire     [31:0] n41320;
wire     [31:0] n41321;
wire     [31:0] n41322;
wire     [31:0] n41323;
wire     [31:0] n41324;
wire     [31:0] n41325;
wire     [31:0] n41326;
wire     [31:0] n41327;
wire     [31:0] n41328;
wire     [31:0] n41329;
wire     [31:0] n41330;
wire     [31:0] n41331;
wire     [31:0] n41332;
wire     [31:0] n41333;
wire     [31:0] n41334;
wire     [31:0] n41335;
wire     [31:0] n41336;
wire     [31:0] n41337;
wire     [31:0] n41338;
wire     [31:0] n41339;
wire     [31:0] n41340;
wire     [31:0] n41341;
wire     [31:0] n41342;
wire     [31:0] n41343;
wire     [31:0] n41344;
wire     [31:0] n41345;
wire     [31:0] n41346;
wire     [31:0] n41347;
wire     [31:0] n41348;
wire     [31:0] n41349;
wire     [31:0] n41350;
wire     [31:0] n41351;
wire     [31:0] n41352;
wire     [31:0] n41353;
wire     [31:0] n41354;
wire     [31:0] n41355;
wire     [31:0] n41356;
wire     [31:0] n41357;
wire     [31:0] n41358;
wire     [31:0] n41359;
wire     [31:0] n41360;
wire     [31:0] n41361;
wire     [31:0] n41362;
wire     [31:0] n41363;
wire     [31:0] n41364;
wire     [31:0] n41365;
wire     [31:0] n41366;
wire     [31:0] n41367;
wire     [31:0] n41368;
wire     [31:0] n41369;
wire     [31:0] n41370;
wire     [31:0] n41371;
wire     [31:0] n41372;
wire     [31:0] n41373;
wire     [31:0] n41374;
wire     [31:0] n41375;
wire     [31:0] n41376;
wire     [31:0] n41377;
wire     [31:0] n41378;
wire     [31:0] n41379;
wire     [31:0] n41380;
wire     [31:0] n41381;
wire     [31:0] n41382;
wire     [31:0] n41383;
wire     [31:0] n41384;
wire     [31:0] n41385;
wire     [31:0] n41386;
wire     [31:0] n41387;
wire     [31:0] n41388;
wire     [31:0] n41389;
wire     [31:0] n41390;
wire     [31:0] n41391;
wire     [31:0] n41392;
wire     [31:0] n41393;
wire     [31:0] n41394;
wire     [31:0] n41395;
wire     [31:0] n41396;
wire     [31:0] n41397;
wire     [31:0] n41398;
wire     [31:0] n41399;
wire     [31:0] n41400;
wire     [31:0] n41401;
wire     [31:0] n41402;
wire     [31:0] n41403;
wire     [31:0] n41404;
wire     [31:0] n41405;
wire     [31:0] n41406;
wire     [31:0] n41407;
wire     [31:0] n41408;
wire     [31:0] n41409;
wire     [31:0] n41410;
wire     [31:0] n41411;
wire     [31:0] n41412;
wire     [31:0] n41413;
wire     [31:0] n41414;
wire     [31:0] n41415;
wire     [31:0] n41416;
wire     [31:0] n41417;
wire     [31:0] n41418;
wire     [31:0] n41419;
wire     [31:0] n41420;
wire     [31:0] n41421;
wire     [31:0] n41422;
wire     [31:0] n41423;
wire     [31:0] n41424;
wire     [31:0] n41425;
wire     [31:0] n41426;
wire     [31:0] n41427;
wire     [31:0] n41428;
wire     [31:0] n41429;
wire     [31:0] n41430;
wire     [31:0] n41431;
wire     [31:0] n41432;
wire     [31:0] n41433;
wire     [31:0] n41434;
wire     [31:0] n41435;
wire     [31:0] n41436;
wire     [31:0] n41437;
wire     [31:0] n41438;
wire     [31:0] n41439;
wire     [31:0] n41440;
wire     [31:0] n41441;
wire     [31:0] n41442;
wire     [31:0] n41443;
wire     [31:0] n41444;
wire     [31:0] n41445;
wire     [31:0] n41446;
wire     [31:0] n41447;
wire     [31:0] n41448;
wire     [31:0] n41449;
wire     [31:0] n41450;
wire     [31:0] n41451;
wire     [31:0] n41452;
wire     [31:0] n41453;
wire     [31:0] n41454;
wire     [31:0] n41455;
wire     [31:0] n41456;
wire     [31:0] n41457;
wire     [31:0] n41458;
wire     [31:0] n41459;
wire     [31:0] n41460;
wire     [31:0] n41461;
wire     [31:0] n41462;
wire     [31:0] n41463;
wire     [31:0] n41464;
wire     [31:0] n41465;
wire     [31:0] n41466;
wire     [31:0] n41467;
wire     [31:0] n41468;
wire     [31:0] n41469;
wire     [31:0] n41470;
wire     [31:0] n41471;
wire     [31:0] n41472;
wire     [31:0] n41473;
wire     [31:0] n41474;
wire     [31:0] n41475;
wire     [31:0] n41476;
wire     [31:0] n41477;
wire     [31:0] n41478;
wire     [31:0] n41479;
wire     [31:0] n41480;
wire     [31:0] n41481;
wire     [31:0] n41482;
wire     [31:0] n41483;
wire     [31:0] n41484;
wire     [31:0] n41485;
wire     [31:0] n41486;
wire     [31:0] n41487;
wire     [31:0] n41488;
wire     [31:0] n41489;
wire     [31:0] n41490;
wire     [31:0] n41491;
wire     [31:0] n41492;
wire     [31:0] n41493;
wire     [31:0] n41494;
wire     [31:0] n41495;
wire     [31:0] n41496;
wire     [31:0] n41497;
wire     [31:0] n41498;
wire     [31:0] n41499;
wire     [31:0] n41500;
wire     [31:0] n41501;
wire     [31:0] n41502;
wire     [31:0] n41503;
wire     [31:0] n41504;
wire     [31:0] n41505;
wire     [31:0] n41506;
wire     [31:0] n41507;
wire     [31:0] n41508;
wire     [31:0] n41509;
wire     [31:0] n41510;
wire     [31:0] n41511;
wire     [31:0] n41512;
wire     [31:0] n41513;
wire     [31:0] n41514;
wire     [31:0] n41515;
wire     [31:0] n41516;
wire     [31:0] n41517;
wire     [31:0] n41518;
wire     [31:0] n41519;
wire     [31:0] n41520;
wire     [31:0] n41521;
wire     [31:0] n41522;
wire     [31:0] n41523;
wire     [31:0] n41524;
wire     [31:0] n41525;
wire     [31:0] n41526;
wire     [31:0] n41527;
wire     [31:0] n41528;
wire     [31:0] n41529;
wire     [31:0] n41530;
wire     [31:0] n41531;
wire     [31:0] n41532;
wire     [31:0] n41533;
wire     [31:0] n41534;
wire     [31:0] n41535;
wire     [31:0] n41536;
wire     [31:0] n41537;
wire     [31:0] n41538;
wire     [31:0] n41539;
wire     [31:0] n41540;
wire     [31:0] n41541;
wire     [31:0] n41542;
wire     [31:0] n41543;
wire     [31:0] n41544;
wire     [31:0] n41545;
wire     [31:0] n41546;
wire     [31:0] n41547;
wire     [31:0] n41548;
wire     [31:0] n41549;
wire     [31:0] n41550;
wire     [31:0] n41551;
wire     [31:0] n41552;
wire     [31:0] n41553;
wire     [31:0] n41554;
wire     [31:0] n41555;
wire     [31:0] n41556;
wire     [31:0] n41557;
wire     [31:0] n41558;
wire     [31:0] n41559;
wire     [31:0] n41560;
wire     [31:0] n41561;
wire     [31:0] n41562;
wire     [31:0] n41563;
wire     [31:0] n41564;
wire     [31:0] n41565;
wire     [31:0] n41566;
wire     [31:0] n41567;
wire     [31:0] n41568;
wire     [31:0] n41569;
wire     [31:0] n41570;
wire     [31:0] n41571;
wire     [31:0] n41572;
wire     [31:0] n41573;
wire     [31:0] n41574;
wire     [31:0] n41575;
wire     [31:0] n41576;
wire     [31:0] n41577;
wire     [31:0] n41578;
wire     [31:0] n41579;
wire     [31:0] n41580;
wire     [31:0] n41581;
wire     [31:0] n41582;
wire     [31:0] n41583;
wire     [31:0] n41584;
wire     [31:0] n41585;
wire     [31:0] n41586;
wire     [31:0] n41587;
wire     [31:0] n41588;
wire     [31:0] n41589;
wire     [31:0] n41590;
wire     [31:0] n41591;
wire     [31:0] n41592;
wire     [31:0] n41593;
wire     [31:0] n41594;
wire     [31:0] n41595;
wire     [31:0] n41596;
wire     [31:0] n41597;
wire     [31:0] n41598;
wire     [31:0] n41599;
wire     [31:0] n41600;
wire     [31:0] n41601;
wire     [31:0] n41602;
wire     [31:0] n41603;
wire     [31:0] n41604;
wire     [31:0] n41605;
wire     [31:0] n41606;
wire     [31:0] n41607;
wire     [31:0] n41608;
wire     [31:0] n41609;
wire     [31:0] n41610;
wire     [31:0] n41611;
wire     [31:0] n41612;
wire     [31:0] n41613;
wire     [31:0] n41614;
wire     [31:0] n41615;
wire     [31:0] n41616;
wire     [31:0] n41617;
wire     [31:0] n41618;
wire     [31:0] n41619;
wire     [31:0] n41620;
wire     [31:0] n41621;
wire     [31:0] n41622;
wire     [31:0] n41623;
wire     [31:0] n41624;
wire     [31:0] n41625;
wire     [31:0] n41626;
wire     [31:0] n41627;
wire     [31:0] n41628;
wire     [31:0] n41629;
wire     [31:0] n41630;
wire     [31:0] n41631;
wire     [31:0] n41632;
wire     [31:0] n41633;
wire     [31:0] n41634;
wire     [31:0] n41635;
wire     [31:0] n41636;
wire     [31:0] n41637;
wire     [31:0] n41638;
wire     [31:0] n41639;
wire     [31:0] n41640;
wire     [31:0] n41641;
wire     [31:0] n41642;
wire     [31:0] n41643;
wire     [31:0] n41644;
wire     [31:0] n41645;
wire     [31:0] n41646;
wire     [31:0] n41647;
wire     [31:0] n41648;
wire     [31:0] n41649;
wire     [31:0] n41650;
wire     [31:0] n41651;
wire     [31:0] n41652;
wire     [31:0] n41653;
wire     [31:0] n41654;
wire     [31:0] n41655;
wire     [31:0] n41656;
wire     [31:0] n41657;
wire     [31:0] n41658;
wire     [31:0] n41659;
wire     [31:0] n41660;
wire     [31:0] n41661;
wire     [31:0] n41662;
wire     [31:0] n41663;
wire     [31:0] n41664;
wire     [31:0] n41665;
wire     [31:0] n41666;
wire     [31:0] n41667;
wire     [31:0] n41668;
wire     [31:0] n41669;
wire     [31:0] n41670;
wire     [31:0] n41671;
wire     [31:0] n41672;
wire     [31:0] n41673;
wire     [31:0] n41674;
wire     [31:0] n41675;
wire     [31:0] n41676;
wire     [31:0] n41677;
wire     [31:0] n41678;
wire     [31:0] n41679;
wire     [31:0] n41680;
wire     [31:0] n41681;
wire     [31:0] n41682;
wire     [31:0] n41683;
wire     [31:0] n41684;
wire     [31:0] n41685;
wire     [31:0] n41686;
wire     [31:0] n41687;
wire     [31:0] n41688;
wire     [31:0] n41689;
wire     [31:0] n41690;
wire     [31:0] n41691;
wire     [31:0] n41692;
wire     [31:0] n41693;
wire     [31:0] n41694;
wire     [31:0] n41695;
wire     [31:0] n41696;
wire     [31:0] n41697;
wire     [31:0] n41698;
wire     [31:0] n41699;
wire     [31:0] n41700;
wire     [31:0] n41701;
wire     [31:0] n41702;
wire     [31:0] n41703;
wire     [31:0] n41704;
wire     [31:0] n41705;
wire     [31:0] n41706;
wire     [31:0] n41707;
wire     [31:0] n41708;
wire     [31:0] n41709;
wire     [31:0] n41710;
wire     [31:0] n41711;
wire     [31:0] n41712;
wire     [31:0] n41713;
wire     [31:0] n41714;
wire     [31:0] n41715;
wire     [31:0] n41716;
wire     [31:0] n41717;
wire     [31:0] n41718;
wire     [31:0] n41719;
wire     [31:0] n41720;
wire     [31:0] n41721;
wire     [31:0] n41722;
wire     [31:0] n41723;
wire     [31:0] n41724;
wire     [31:0] n41725;
wire     [31:0] n41726;
wire     [31:0] n41727;
wire     [31:0] n41728;
wire     [31:0] n41729;
wire     [31:0] n41730;
wire     [31:0] n41731;
wire     [31:0] n41732;
wire     [31:0] n41733;
wire     [31:0] n41734;
wire     [31:0] n41735;
wire     [31:0] n41736;
wire     [31:0] n41737;
wire     [31:0] n41738;
wire     [31:0] n41739;
wire     [31:0] n41740;
wire     [31:0] n41741;
wire     [31:0] n41742;
wire     [31:0] n41743;
wire     [31:0] n41744;
wire     [31:0] n41745;
wire     [31:0] n41746;
wire     [31:0] n41747;
wire     [31:0] n41748;
wire     [31:0] n41749;
wire     [31:0] n41750;
wire     [31:0] n41751;
wire     [31:0] n41752;
wire     [31:0] n41753;
wire     [31:0] n41754;
wire     [31:0] n41755;
wire     [31:0] n41756;
wire     [31:0] n41757;
wire     [31:0] n41758;
wire     [31:0] n41759;
wire     [31:0] n41760;
wire     [31:0] n41761;
wire     [31:0] n41762;
wire     [31:0] n41763;
wire     [31:0] n41764;
wire     [31:0] n41765;
wire     [31:0] n41766;
wire     [31:0] n41767;
wire     [31:0] n41768;
wire     [31:0] n41769;
wire     [31:0] n41770;
wire     [31:0] n41771;
wire     [31:0] n41772;
wire     [31:0] n41773;
wire     [31:0] n41774;
wire     [31:0] n41775;
wire     [31:0] n41776;
wire     [31:0] n41777;
wire     [31:0] n41778;
wire     [31:0] n41779;
wire     [31:0] n41780;
wire     [31:0] n41781;
wire     [31:0] n41782;
wire     [31:0] n41783;
wire     [31:0] n41784;
wire     [31:0] n41785;
wire     [31:0] n41786;
wire     [31:0] n41787;
wire     [31:0] n41788;
wire     [31:0] n41789;
wire     [31:0] n41790;
wire     [31:0] n41791;
wire     [31:0] n41792;
wire     [31:0] n41793;
wire     [31:0] n41794;
wire     [31:0] n41795;
wire     [31:0] n41796;
wire     [31:0] n41797;
wire     [31:0] n41798;
wire     [31:0] n41799;
wire     [31:0] n41800;
wire     [31:0] n41801;
wire     [31:0] n41802;
wire     [31:0] n41803;
wire     [31:0] n41804;
wire     [31:0] n41805;
wire     [31:0] n41806;
wire     [31:0] n41807;
wire     [31:0] n41808;
wire     [31:0] n41809;
wire     [31:0] n41810;
wire     [31:0] n41811;
wire     [31:0] n41812;
wire     [31:0] n41813;
wire     [31:0] n41814;
wire     [31:0] n41815;
wire     [31:0] n41816;
wire     [31:0] n41817;
wire     [31:0] n41818;
wire     [31:0] n41819;
wire     [31:0] n41820;
wire     [31:0] n41821;
wire     [31:0] n41822;
wire     [31:0] n41823;
wire     [31:0] n41824;
wire     [31:0] n41825;
wire     [31:0] n41826;
wire     [31:0] n41827;
wire     [31:0] n41828;
wire     [31:0] n41829;
wire     [31:0] n41830;
wire     [31:0] n41831;
wire     [31:0] n41832;
wire     [31:0] n41833;
wire     [31:0] n41834;
wire     [31:0] n41835;
wire     [31:0] n41836;
wire     [31:0] n41837;
wire     [31:0] n41838;
wire     [31:0] n41839;
wire     [31:0] n41840;
wire     [31:0] n41841;
wire     [31:0] n41842;
wire     [31:0] n41843;
wire     [31:0] n41844;
wire     [31:0] n41845;
wire     [31:0] n41846;
wire     [31:0] n41847;
wire     [31:0] n41848;
wire     [31:0] n41849;
wire     [31:0] n41850;
wire     [31:0] n41851;
wire     [31:0] n41852;
wire     [31:0] n41853;
wire     [31:0] n41854;
wire     [31:0] n41855;
wire     [31:0] n41856;
wire     [31:0] n41857;
wire     [31:0] n41858;
wire     [31:0] n41859;
wire     [31:0] n41860;
wire     [31:0] n41861;
wire     [31:0] n41862;
wire     [31:0] n41863;
wire     [31:0] n41864;
wire     [31:0] n41865;
wire     [31:0] n41866;
wire     [31:0] n41867;
wire     [31:0] n41868;
wire     [31:0] n41869;
wire     [31:0] n41870;
wire     [31:0] n41871;
wire     [31:0] n41872;
wire     [31:0] n41873;
wire     [31:0] n41874;
wire     [31:0] n41875;
wire     [31:0] n41876;
wire     [31:0] n41877;
wire     [31:0] n41878;
wire     [31:0] n41879;
wire     [31:0] n41880;
wire     [31:0] n41881;
wire     [31:0] n41882;
wire     [31:0] n41883;
wire     [31:0] n41884;
wire     [31:0] n41885;
wire     [31:0] n41886;
wire     [31:0] n41887;
wire     [31:0] n41888;
wire     [31:0] n41889;
wire     [31:0] n41890;
wire     [31:0] n41891;
wire     [31:0] n41892;
wire     [31:0] n41893;
wire     [31:0] n41894;
wire     [31:0] n41895;
wire     [31:0] n41896;
wire     [31:0] n41897;
wire     [31:0] n41898;
wire     [31:0] n41899;
wire     [31:0] n41900;
wire     [31:0] n41901;
wire     [31:0] n41902;
wire     [31:0] n41903;
wire     [31:0] n41904;
wire     [31:0] n41905;
wire     [31:0] n41906;
wire     [31:0] n41907;
wire     [31:0] n41908;
wire     [31:0] n41909;
wire     [31:0] n41910;
wire     [31:0] n41911;
wire     [31:0] n41912;
wire     [31:0] n41913;
wire     [31:0] n41914;
wire     [31:0] n41915;
wire     [31:0] n41916;
wire     [31:0] n41917;
wire     [31:0] n41918;
wire     [31:0] n41919;
wire     [31:0] n41920;
wire     [31:0] n41921;
wire     [31:0] n41922;
wire     [31:0] n41923;
wire     [31:0] n41924;
wire     [31:0] n41925;
wire     [31:0] n41926;
wire     [31:0] n41927;
wire     [31:0] n41928;
wire     [31:0] n41929;
wire     [31:0] n41930;
wire     [31:0] n41931;
wire     [31:0] n41932;
wire     [31:0] n41933;
wire     [31:0] n41934;
wire     [31:0] n41935;
wire     [31:0] n41936;
wire     [31:0] n41937;
wire     [31:0] n41938;
wire     [31:0] n41939;
wire     [31:0] n41940;
wire     [31:0] n41941;
wire     [31:0] n41942;
wire     [31:0] n41943;
wire     [31:0] n41944;
wire     [31:0] n41945;
wire     [31:0] n41946;
wire     [31:0] n41947;
wire     [31:0] n41948;
wire     [31:0] n41949;
wire     [31:0] n41950;
wire     [31:0] n41951;
wire     [31:0] n41952;
wire     [31:0] n41953;
wire     [31:0] n41954;
wire     [31:0] n41955;
wire     [31:0] n41956;
wire     [31:0] n41957;
wire     [31:0] n41958;
wire     [31:0] n41959;
wire     [31:0] n41960;
wire     [31:0] n41961;
wire     [31:0] n41962;
wire     [31:0] n41963;
wire     [31:0] n41964;
wire     [31:0] n41965;
wire     [31:0] n41966;
wire     [31:0] n41967;
wire     [31:0] n41968;
wire     [31:0] n41969;
wire     [31:0] n41970;
wire     [31:0] n41971;
wire     [31:0] n41972;
wire     [31:0] n41973;
wire     [31:0] n41974;
wire     [31:0] n41975;
wire     [31:0] n41976;
wire     [31:0] n41977;
wire     [31:0] n41978;
wire     [31:0] n41979;
wire     [31:0] n41980;
wire     [31:0] n41981;
wire     [31:0] n41982;
wire     [31:0] n41983;
wire     [31:0] n41984;
wire     [31:0] n41985;
wire     [31:0] n41986;
wire     [31:0] n41987;
wire     [31:0] n41988;
wire     [31:0] n41989;
wire     [31:0] n41990;
wire     [31:0] n41991;
wire     [31:0] n41992;
wire     [31:0] n41993;
wire     [31:0] n41994;
wire     [31:0] n41995;
wire     [31:0] n41996;
wire     [31:0] n41997;
wire     [31:0] n41998;
wire     [31:0] n41999;
wire     [31:0] n42000;
wire     [31:0] n42001;
wire     [31:0] n42002;
wire     [31:0] n42003;
wire     [31:0] n42004;
wire     [31:0] n42005;
wire     [31:0] n42006;
wire     [31:0] n42007;
wire     [31:0] n42008;
wire     [31:0] n42009;
wire     [31:0] n42010;
wire     [31:0] n42011;
wire     [31:0] n42012;
wire     [31:0] n42013;
wire     [31:0] n42014;
wire     [31:0] n42015;
wire     [31:0] n42016;
wire     [31:0] n42017;
wire     [31:0] n42018;
wire     [31:0] n42019;
wire     [31:0] n42020;
wire     [31:0] n42021;
wire     [31:0] n42022;
wire     [31:0] n42023;
wire     [31:0] n42024;
wire     [31:0] n42025;
wire     [31:0] n42026;
wire     [31:0] n42027;
wire     [31:0] n42028;
wire     [31:0] n42029;
wire     [31:0] n42030;
wire     [31:0] n42031;
wire     [31:0] n42032;
wire     [31:0] n42033;
wire     [31:0] n42034;
wire     [31:0] n42035;
wire     [31:0] n42036;
wire     [31:0] n42037;
wire     [31:0] n42038;
wire     [31:0] n42039;
wire     [31:0] n42040;
wire     [31:0] n42041;
wire     [31:0] n42042;
wire     [31:0] n42043;
wire     [31:0] n42044;
wire     [31:0] n42045;
wire     [31:0] n42046;
wire     [31:0] n42047;
wire     [31:0] n42048;
wire     [31:0] n42049;
wire     [31:0] n42050;
wire     [31:0] n42051;
wire     [31:0] n42052;
wire     [31:0] n42053;
wire     [31:0] n42054;
wire     [31:0] n42055;
wire     [31:0] n42056;
wire     [31:0] n42057;
wire     [31:0] n42058;
wire     [31:0] n42059;
wire     [31:0] n42060;
wire     [31:0] n42061;
wire     [31:0] n42062;
wire     [31:0] n42063;
wire     [31:0] n42064;
wire     [31:0] n42065;
wire     [31:0] n42066;
wire     [31:0] n42067;
wire     [31:0] n42068;
wire     [31:0] n42069;
wire     [31:0] n42070;
wire     [31:0] n42071;
wire     [31:0] n42072;
wire     [31:0] n42073;
wire     [31:0] n42074;
wire     [31:0] n42075;
wire     [31:0] n42076;
wire     [31:0] n42077;
wire     [31:0] n42078;
wire     [31:0] n42079;
wire     [31:0] n42080;
wire     [31:0] n42081;
wire     [31:0] n42082;
wire     [31:0] n42083;
wire     [31:0] n42084;
wire     [31:0] n42085;
wire     [31:0] n42086;
wire     [31:0] n42087;
wire     [31:0] n42088;
wire     [31:0] n42089;
wire     [31:0] n42090;
wire     [31:0] n42091;
wire     [31:0] n42092;
wire     [31:0] n42093;
wire     [31:0] n42094;
wire     [31:0] n42095;
wire     [31:0] n42096;
wire     [31:0] n42097;
wire     [31:0] n42098;
wire     [31:0] n42099;
wire     [31:0] n42100;
wire     [31:0] n42101;
wire     [31:0] n42102;
wire     [31:0] n42103;
wire     [31:0] n42104;
wire     [31:0] n42105;
wire     [31:0] n42106;
wire     [31:0] n42107;
wire     [31:0] n42108;
wire     [31:0] n42109;
wire     [31:0] n42110;
wire     [31:0] n42111;
wire     [31:0] n42112;
wire     [31:0] n42113;
wire     [31:0] n42114;
wire     [31:0] n42115;
wire     [31:0] n42116;
wire     [31:0] n42117;
wire     [31:0] n42118;
wire     [31:0] n42119;
wire     [31:0] n42120;
wire     [31:0] n42121;
wire     [31:0] n42122;
wire     [31:0] n42123;
wire     [31:0] n42124;
wire     [31:0] n42125;
wire     [31:0] n42126;
wire     [31:0] n42127;
wire     [31:0] n42128;
wire     [31:0] n42129;
wire     [31:0] n42130;
wire     [31:0] n42131;
wire     [31:0] n42132;
wire     [31:0] n42133;
wire     [31:0] n42134;
wire     [31:0] n42135;
wire     [31:0] n42136;
wire     [31:0] n42137;
wire     [31:0] n42138;
wire     [31:0] n42139;
wire     [31:0] n42140;
wire     [31:0] n42141;
wire     [31:0] n42142;
wire     [31:0] n42143;
wire     [31:0] n42144;
wire     [31:0] n42145;
wire     [31:0] n42146;
wire     [31:0] n42147;
wire     [31:0] n42148;
wire     [31:0] n42149;
wire     [31:0] n42150;
wire     [31:0] n42151;
wire     [31:0] n42152;
wire     [31:0] n42153;
wire     [31:0] n42154;
wire     [31:0] n42155;
wire     [31:0] n42156;
wire     [31:0] n42157;
wire     [31:0] n42158;
wire     [31:0] n42159;
wire     [31:0] n42160;
wire     [31:0] n42161;
wire     [31:0] n42162;
wire     [31:0] n42163;
wire     [31:0] n42164;
wire     [31:0] n42165;
wire     [31:0] n42166;
wire     [31:0] n42167;
wire     [31:0] n42168;
wire     [31:0] n42169;
wire     [31:0] n42170;
wire     [31:0] n42171;
wire     [31:0] n42172;
wire     [31:0] n42173;
wire     [31:0] n42174;
wire     [31:0] n42175;
wire     [31:0] n42176;
wire     [31:0] n42177;
wire     [31:0] n42178;
wire     [31:0] n42179;
wire     [31:0] n42180;
wire     [31:0] n42181;
wire     [31:0] n42182;
wire     [31:0] n42183;
wire     [31:0] n42184;
wire     [31:0] n42185;
wire     [31:0] n42186;
wire     [31:0] n42187;
wire     [31:0] n42188;
wire     [31:0] n42189;
wire     [31:0] n42190;
wire     [31:0] n42191;
wire     [31:0] n42192;
wire     [31:0] n42193;
wire     [31:0] n42194;
wire     [31:0] n42195;
wire     [31:0] n42196;
wire     [31:0] n42197;
wire     [31:0] n42198;
wire     [31:0] n42199;
wire     [31:0] n42200;
wire     [31:0] n42201;
wire     [31:0] n42202;
wire     [31:0] n42203;
wire     [31:0] n42204;
wire     [31:0] n42205;
wire     [31:0] n42206;
wire     [31:0] n42207;
wire     [31:0] n42208;
wire     [31:0] n42209;
wire     [31:0] n42210;
wire     [31:0] n42211;
wire     [31:0] n42212;
wire     [31:0] n42213;
wire     [31:0] n42214;
wire     [31:0] n42215;
wire     [31:0] n42216;
wire     [31:0] n42217;
wire     [31:0] n42218;
wire     [31:0] n42219;
wire     [31:0] n42220;
wire     [31:0] n42221;
wire     [31:0] n42222;
wire     [31:0] n42223;
wire     [31:0] n42224;
wire     [31:0] n42225;
wire     [31:0] n42226;
wire     [31:0] n42227;
wire     [31:0] n42228;
wire     [31:0] n42229;
wire     [31:0] n42230;
wire     [31:0] n42231;
wire     [31:0] n42232;
wire     [31:0] n42233;
wire     [31:0] n42234;
wire     [31:0] n42235;
wire     [31:0] n42236;
wire     [31:0] n42237;
wire     [31:0] n42238;
wire     [31:0] n42239;
wire     [31:0] n42240;
wire     [31:0] n42241;
wire     [31:0] n42242;
wire     [31:0] n42243;
wire     [31:0] n42244;
wire     [31:0] n42245;
wire     [31:0] n42246;
wire     [31:0] n42247;
wire     [31:0] n42248;
wire     [31:0] n42249;
wire     [31:0] n42250;
wire     [31:0] n42251;
wire     [31:0] n42252;
wire     [31:0] n42253;
wire     [31:0] n42254;
wire     [31:0] n42255;
wire     [31:0] n42256;
wire     [31:0] n42257;
wire     [31:0] n42258;
wire     [31:0] n42259;
wire     [31:0] n42260;
wire     [31:0] n42261;
wire     [31:0] n42262;
wire     [31:0] n42263;
wire     [31:0] n42264;
wire     [31:0] n42265;
wire     [31:0] n42266;
wire     [31:0] n42267;
wire     [31:0] n42268;
wire     [31:0] n42269;
wire     [31:0] n42270;
wire     [31:0] n42271;
wire     [31:0] n42272;
wire     [31:0] n42273;
wire     [31:0] n42274;
wire     [31:0] n42275;
wire     [31:0] n42276;
wire     [31:0] n42277;
wire     [31:0] n42278;
wire     [31:0] n42279;
wire     [31:0] n42280;
wire     [31:0] n42281;
wire     [31:0] n42282;
wire     [31:0] n42283;
wire     [31:0] n42284;
wire     [31:0] n42285;
wire     [31:0] n42286;
wire     [31:0] n42287;
wire     [31:0] n42288;
wire     [31:0] n42289;
wire     [31:0] n42290;
wire     [31:0] n42291;
wire     [31:0] n42292;
wire     [31:0] n42293;
wire     [31:0] n42294;
wire     [31:0] n42295;
wire     [31:0] n42296;
wire     [31:0] n42297;
wire     [31:0] n42298;
wire     [31:0] n42299;
wire     [31:0] n42300;
wire     [31:0] n42301;
wire     [31:0] n42302;
wire     [31:0] n42303;
wire     [31:0] n42304;
wire     [31:0] n42305;
wire     [31:0] n42306;
wire     [31:0] n42307;
wire     [31:0] n42308;
wire     [31:0] n42309;
wire     [31:0] n42310;
wire     [31:0] n42311;
wire     [31:0] n42312;
wire     [31:0] n42313;
wire     [31:0] n42314;
wire     [31:0] n42315;
wire     [31:0] n42316;
wire     [31:0] n42317;
wire     [31:0] n42318;
wire     [31:0] n42319;
wire     [31:0] n42320;
wire     [31:0] n42321;
wire     [31:0] n42322;
wire     [31:0] n42323;
wire     [31:0] n42324;
wire     [31:0] n42325;
wire     [31:0] n42326;
wire     [31:0] n42327;
wire     [31:0] n42328;
wire     [31:0] n42329;
wire     [31:0] n42330;
wire     [31:0] n42331;
wire     [31:0] n42332;
wire     [31:0] n42333;
wire     [31:0] n42334;
wire     [31:0] n42335;
wire     [31:0] n42336;
wire     [31:0] n42337;
wire     [31:0] n42338;
wire     [31:0] n42339;
wire     [31:0] n42340;
wire     [31:0] n42341;
wire     [31:0] n42342;
wire     [31:0] n42343;
wire     [31:0] n42344;
wire     [31:0] n42345;
wire     [31:0] n42346;
wire     [31:0] n42347;
wire     [31:0] n42348;
wire     [31:0] n42349;
wire     [31:0] n42350;
wire     [31:0] n42351;
wire     [31:0] n42352;
wire     [31:0] n42353;
wire     [31:0] n42354;
wire     [31:0] n42355;
wire     [31:0] n42356;
wire     [31:0] n42357;
wire     [31:0] n42358;
wire     [31:0] n42359;
wire     [31:0] n42360;
wire     [31:0] n42361;
wire     [31:0] n42362;
wire     [31:0] n42363;
wire     [31:0] n42364;
wire     [31:0] n42365;
wire     [31:0] n42366;
wire     [31:0] n42367;
wire     [31:0] n42368;
wire     [31:0] n42369;
wire     [31:0] n42370;
wire     [31:0] n42371;
wire     [31:0] n42372;
wire     [31:0] n42373;
wire     [31:0] n42374;
wire     [31:0] n42375;
wire     [31:0] n42376;
wire     [31:0] n42377;
wire     [31:0] n42378;
wire     [31:0] n42379;
wire     [31:0] n42380;
wire     [31:0] n42381;
wire     [31:0] n42382;
wire     [31:0] n42383;
wire     [31:0] n42384;
wire     [31:0] n42385;
wire     [31:0] n42386;
wire     [31:0] n42387;
wire     [31:0] n42388;
wire     [31:0] n42389;
wire     [31:0] n42390;
wire     [31:0] n42391;
wire     [31:0] n42392;
wire     [31:0] n42393;
wire     [31:0] n42394;
wire     [31:0] n42395;
wire     [31:0] n42396;
wire     [31:0] n42397;
wire     [31:0] n42398;
wire     [31:0] n42399;
wire     [31:0] n42400;
wire     [31:0] n42401;
wire     [31:0] n42402;
wire     [31:0] n42403;
wire     [31:0] n42404;
wire     [31:0] n42405;
wire     [31:0] n42406;
wire     [31:0] n42407;
wire     [31:0] n42408;
wire     [31:0] n42409;
wire     [31:0] n42410;
wire     [31:0] n42411;
wire     [31:0] n42412;
wire     [31:0] n42413;
wire     [31:0] n42414;
wire     [31:0] n42415;
wire     [31:0] n42416;
wire     [31:0] n42417;
wire     [31:0] n42418;
wire     [31:0] n42419;
wire     [31:0] n42420;
wire     [31:0] n42421;
wire     [31:0] n42422;
wire     [31:0] n42423;
wire     [31:0] n42424;
wire     [31:0] n42425;
wire     [31:0] n42426;
wire     [31:0] n42427;
wire     [31:0] n42428;
wire     [31:0] n42429;
wire     [31:0] n42430;
wire     [31:0] n42431;
wire     [31:0] n42432;
wire     [31:0] n42433;
wire     [31:0] n42434;
wire     [31:0] n42435;
wire     [31:0] n42436;
wire     [31:0] n42437;
wire     [31:0] n42438;
wire     [31:0] n42439;
wire     [31:0] n42440;
wire     [31:0] n42441;
wire     [31:0] n42442;
wire     [31:0] n42443;
wire     [31:0] n42444;
wire     [31:0] n42445;
wire     [31:0] n42446;
wire     [31:0] n42447;
wire     [31:0] n42448;
wire     [31:0] n42449;
wire     [31:0] n42450;
wire     [31:0] n42451;
wire     [31:0] n42452;
wire     [31:0] n42453;
wire     [31:0] n42454;
wire     [31:0] n42455;
wire     [31:0] n42456;
wire     [31:0] n42457;
wire     [31:0] n42458;
wire     [31:0] n42459;
wire     [31:0] n42460;
wire     [31:0] n42461;
wire     [31:0] n42462;
wire     [31:0] n42463;
wire     [31:0] n42464;
wire     [31:0] n42465;
wire     [31:0] n42466;
wire     [31:0] n42467;
wire     [31:0] n42468;
wire     [31:0] n42469;
wire     [31:0] n42470;
wire     [31:0] n42471;
wire     [31:0] n42472;
wire     [31:0] n42473;
wire     [31:0] n42474;
wire     [31:0] n42475;
wire     [31:0] n42476;
wire     [31:0] n42477;
wire     [31:0] n42478;
wire     [31:0] n42479;
wire     [31:0] n42480;
wire     [31:0] n42481;
wire     [31:0] n42482;
wire     [31:0] n42483;
wire     [31:0] n42484;
wire     [31:0] n42485;
wire     [31:0] n42486;
wire     [31:0] n42487;
wire     [31:0] n42488;
wire     [31:0] n42489;
wire     [31:0] n42490;
wire     [31:0] n42491;
wire     [31:0] n42492;
wire     [31:0] n42493;
wire     [31:0] n42494;
wire     [31:0] n42495;
wire     [31:0] n42496;
wire     [31:0] n42497;
wire     [31:0] n42498;
wire     [31:0] n42499;
wire     [31:0] n42500;
wire     [31:0] n42501;
wire     [31:0] n42502;
wire     [31:0] n42503;
wire     [31:0] n42504;
wire     [31:0] n42505;
wire     [31:0] n42506;
wire     [31:0] n42507;
wire     [31:0] n42508;
wire     [31:0] n42509;
wire     [31:0] n42510;
wire     [31:0] n42511;
wire     [31:0] n42512;
wire     [31:0] n42513;
wire     [31:0] n42514;
wire     [31:0] n42515;
wire     [31:0] n42516;
wire     [31:0] n42517;
wire     [31:0] n42518;
wire     [31:0] n42519;
wire     [31:0] n42520;
wire     [31:0] n42521;
wire     [31:0] n42522;
wire     [31:0] n42523;
wire     [31:0] n42524;
wire     [31:0] n42525;
wire     [31:0] n42526;
wire     [31:0] n42527;
wire     [31:0] n42528;
wire     [31:0] n42529;
wire     [31:0] n42530;
wire     [31:0] n42531;
wire     [31:0] n42532;
wire     [31:0] n42533;
wire     [31:0] n42534;
wire     [31:0] n42535;
wire     [31:0] n42536;
wire     [31:0] n42537;
wire     [31:0] n42538;
wire     [31:0] n42539;
wire     [31:0] n42540;
wire     [31:0] n42541;
wire     [31:0] n42542;
wire     [31:0] n42543;
wire     [31:0] n42544;
wire     [31:0] n42545;
wire     [31:0] n42546;
wire     [31:0] n42547;
wire     [31:0] n42548;
wire     [31:0] n42549;
wire     [31:0] n42550;
wire     [31:0] n42551;
wire     [31:0] n42552;
wire     [31:0] n42553;
wire     [31:0] n42554;
wire     [31:0] n42555;
wire     [31:0] n42556;
wire     [31:0] n42557;
wire     [31:0] n42558;
wire     [31:0] n42559;
wire     [31:0] n42560;
wire     [31:0] n42561;
wire     [31:0] n42562;
wire     [31:0] n42563;
wire     [31:0] n42564;
wire     [31:0] n42565;
wire     [31:0] n42566;
wire     [31:0] n42567;
wire     [31:0] n42568;
wire     [31:0] n42569;
wire     [31:0] n42570;
wire     [31:0] n42571;
wire     [31:0] n42572;
wire     [31:0] n42573;
wire     [31:0] n42574;
wire     [31:0] n42575;
wire     [31:0] n42576;
wire     [31:0] n42577;
wire     [31:0] n42578;
wire     [31:0] n42579;
wire     [31:0] n42580;
wire     [31:0] n42581;
wire     [31:0] n42582;
wire     [31:0] n42583;
wire     [31:0] n42584;
wire     [31:0] n42585;
wire     [31:0] n42586;
wire     [31:0] n42587;
wire     [31:0] n42588;
wire     [31:0] n42589;
wire     [31:0] n42590;
wire     [31:0] n42591;
wire     [31:0] n42592;
wire     [31:0] n42593;
wire     [31:0] n42594;
wire     [31:0] n42595;
wire     [31:0] n42596;
wire     [31:0] n42597;
wire     [31:0] n42598;
wire     [31:0] n42599;
wire     [31:0] n42600;
wire     [31:0] n42601;
wire     [31:0] n42602;
wire     [31:0] n42603;
wire     [31:0] n42604;
wire     [31:0] n42605;
wire     [31:0] n42606;
wire     [31:0] n42607;
wire     [31:0] n42608;
wire     [31:0] n42609;
wire     [31:0] n42610;
wire     [31:0] n42611;
wire     [31:0] n42612;
wire     [31:0] n42613;
wire     [31:0] n42614;
wire     [31:0] n42615;
wire     [31:0] n42616;
wire     [31:0] n42617;
wire     [31:0] n42618;
wire     [31:0] n42619;
wire     [31:0] n42620;
wire     [31:0] n42621;
wire     [31:0] n42622;
wire     [31:0] n42623;
wire     [31:0] n42624;
wire     [31:0] n42625;
wire     [31:0] n42626;
wire     [31:0] n42627;
wire     [31:0] n42628;
wire     [31:0] n42629;
wire     [31:0] n42630;
wire     [31:0] n42631;
wire     [31:0] n42632;
wire     [31:0] n42633;
wire     [31:0] n42634;
wire     [31:0] n42635;
wire     [31:0] n42636;
wire     [31:0] n42637;
wire     [31:0] n42638;
wire     [31:0] n42639;
wire     [31:0] n42640;
wire     [31:0] n42641;
wire     [31:0] n42642;
wire     [31:0] n42643;
wire     [31:0] n42644;
wire     [31:0] n42645;
wire     [31:0] n42646;
wire     [31:0] n42647;
wire     [31:0] n42648;
wire     [31:0] n42649;
wire     [31:0] n42650;
wire     [31:0] n42651;
wire     [31:0] n42652;
wire     [31:0] n42653;
wire     [31:0] n42654;
wire     [31:0] n42655;
wire     [31:0] n42656;
wire     [31:0] n42657;
wire     [31:0] n42658;
wire     [31:0] n42659;
wire     [31:0] n42660;
wire     [31:0] n42661;
wire     [31:0] n42662;
wire     [31:0] n42663;
wire     [31:0] n42664;
wire     [31:0] n42665;
wire     [31:0] n42666;
wire     [31:0] n42667;
wire     [31:0] n42668;
wire     [31:0] n42669;
wire     [31:0] n42670;
wire     [31:0] n42671;
wire     [31:0] n42672;
wire     [31:0] n42673;
wire     [31:0] n42674;
wire     [31:0] n42675;
wire     [31:0] n42676;
wire     [31:0] n42677;
wire     [31:0] n42678;
wire     [31:0] n42679;
wire     [31:0] n42680;
wire     [31:0] n42681;
wire     [31:0] n42682;
wire     [31:0] n42683;
wire     [31:0] n42684;
wire     [31:0] n42685;
wire     [31:0] n42686;
wire     [31:0] n42687;
wire     [31:0] n42688;
wire     [31:0] n42689;
wire     [31:0] n42690;
wire     [31:0] n42691;
wire     [31:0] n42692;
wire     [31:0] n42693;
wire     [31:0] n42694;
wire     [31:0] n42695;
wire     [31:0] n42696;
wire     [31:0] n42697;
wire     [31:0] n42698;
wire     [31:0] n42699;
wire     [31:0] n42700;
wire     [31:0] n42701;
wire     [31:0] n42702;
wire     [31:0] n42703;
wire     [31:0] n42704;
wire     [31:0] n42705;
wire     [31:0] n42706;
wire     [31:0] n42707;
wire     [31:0] n42708;
wire     [31:0] n42709;
wire     [31:0] n42710;
wire     [31:0] n42711;
wire     [31:0] n42712;
wire     [31:0] n42713;
wire     [31:0] n42714;
wire     [31:0] n42715;
wire     [31:0] n42716;
wire     [31:0] n42717;
wire     [31:0] n42718;
wire     [31:0] n42719;
wire     [31:0] n42720;
wire     [31:0] n42721;
wire     [31:0] n42722;
wire     [31:0] n42723;
wire     [31:0] n42724;
wire     [31:0] n42725;
wire     [31:0] n42726;
wire     [31:0] n42727;
wire     [31:0] n42728;
wire     [31:0] n42729;
wire     [31:0] n42730;
wire     [31:0] n42731;
wire     [31:0] n42732;
wire     [31:0] n42733;
wire     [31:0] n42734;
wire     [31:0] n42735;
wire     [31:0] n42736;
wire     [31:0] n42737;
wire     [31:0] n42738;
wire     [31:0] n42739;
wire     [31:0] n42740;
wire     [31:0] n42741;
wire     [31:0] n42742;
wire     [31:0] n42743;
wire     [31:0] n42744;
wire     [31:0] n42745;
wire     [31:0] n42746;
wire     [31:0] n42747;
wire     [31:0] n42748;
wire     [31:0] n42749;
wire     [31:0] n42750;
wire     [31:0] n42751;
wire     [31:0] n42752;
wire     [31:0] n42753;
wire     [31:0] n42754;
wire     [31:0] n42755;
wire     [31:0] n42756;
wire     [31:0] n42757;
wire     [31:0] n42758;
wire     [31:0] n42759;
wire     [31:0] n42760;
wire     [31:0] n42761;
wire     [31:0] n42762;
wire     [31:0] n42763;
wire     [31:0] n42764;
wire     [31:0] n42765;
wire     [31:0] n42766;
wire     [31:0] n42767;
wire     [31:0] n42768;
wire     [31:0] n42769;
wire     [31:0] n42770;
wire     [31:0] n42771;
wire     [31:0] n42772;
wire     [31:0] n42773;
wire     [31:0] n42774;
wire     [31:0] n42775;
wire     [31:0] n42776;
wire     [31:0] n42777;
wire     [31:0] n42778;
wire     [31:0] n42779;
wire     [31:0] n42780;
wire     [31:0] n42781;
wire     [31:0] n42782;
wire     [31:0] n42783;
wire     [31:0] n42784;
wire     [31:0] n42785;
wire     [31:0] n42786;
wire     [31:0] n42787;
wire     [31:0] n42788;
wire     [31:0] n42789;
wire     [31:0] n42790;
wire     [31:0] n42791;
wire     [31:0] n42792;
wire     [31:0] n42793;
wire     [31:0] n42794;
wire     [31:0] n42795;
wire     [31:0] n42796;
wire     [31:0] n42797;
wire     [31:0] n42798;
wire     [31:0] n42799;
wire     [31:0] n42800;
wire     [31:0] n42801;
wire     [31:0] n42802;
wire     [31:0] n42803;
wire     [31:0] n42804;
wire     [31:0] n42805;
wire     [31:0] n42806;
wire     [31:0] n42807;
wire     [31:0] n42808;
wire     [31:0] n42809;
wire     [31:0] n42810;
wire     [31:0] n42811;
wire     [31:0] n42812;
wire     [31:0] n42813;
wire     [31:0] n42814;
wire     [31:0] n42815;
wire     [31:0] n42816;
wire     [31:0] n42817;
wire     [31:0] n42818;
wire     [31:0] n42819;
wire     [31:0] n42820;
wire     [31:0] n42821;
wire     [31:0] n42822;
wire     [31:0] n42823;
wire     [31:0] n42824;
wire     [31:0] n42825;
wire     [31:0] n42826;
wire     [31:0] n42827;
wire     [31:0] n42828;
wire     [31:0] n42829;
wire     [31:0] n42830;
wire     [31:0] n42831;
wire     [31:0] n42832;
wire     [31:0] n42833;
wire     [31:0] n42834;
wire     [31:0] n42835;
wire     [31:0] n42836;
wire     [31:0] n42837;
wire     [31:0] n42838;
wire     [31:0] n42839;
wire     [31:0] n42840;
wire     [31:0] n42841;
wire     [31:0] n42842;
wire     [31:0] n42843;
wire     [31:0] n42844;
wire     [31:0] n42845;
wire     [31:0] n42846;
wire     [31:0] n42847;
wire     [31:0] n42848;
wire     [31:0] n42849;
wire     [31:0] n42850;
wire     [31:0] n42851;
wire     [31:0] n42852;
wire     [31:0] n42853;
wire     [31:0] n42854;
wire     [31:0] n42855;
wire     [31:0] n42856;
wire     [31:0] n42857;
wire     [31:0] n42858;
wire     [31:0] n42859;
wire     [31:0] n42860;
wire     [31:0] n42861;
wire     [31:0] n42862;
wire     [31:0] n42863;
wire     [31:0] n42864;
wire     [31:0] n42865;
wire     [31:0] n42866;
wire     [31:0] n42867;
wire     [31:0] n42868;
wire     [31:0] n42869;
wire     [31:0] n42870;
wire     [31:0] n42871;
wire     [31:0] n42872;
wire     [31:0] n42873;
wire     [31:0] n42874;
wire     [31:0] n42875;
wire     [31:0] n42876;
wire     [31:0] n42877;
wire     [31:0] n42878;
wire     [31:0] n42879;
wire     [31:0] n42880;
wire     [31:0] n42881;
wire     [31:0] n42882;
wire     [31:0] n42883;
wire     [31:0] n42884;
wire     [31:0] n42885;
wire     [31:0] n42886;
wire     [31:0] n42887;
wire     [31:0] n42888;
wire     [31:0] n42889;
wire     [31:0] n42890;
wire     [31:0] n42891;
wire     [31:0] n42892;
wire     [31:0] n42893;
wire     [31:0] n42894;
wire     [31:0] n42895;
wire     [31:0] n42896;
wire     [31:0] n42897;
wire     [31:0] n42898;
wire     [31:0] n42899;
wire     [31:0] n42900;
wire     [31:0] n42901;
wire     [31:0] n42902;
wire     [31:0] n42903;
wire     [31:0] n42904;
wire     [31:0] n42905;
wire     [31:0] n42906;
wire     [31:0] n42907;
wire     [31:0] n42908;
wire     [31:0] n42909;
wire     [31:0] n42910;
wire     [31:0] n42911;
wire     [31:0] n42912;
wire     [31:0] n42913;
wire     [31:0] n42914;
wire     [31:0] n42915;
wire     [31:0] n42916;
wire     [31:0] n42917;
wire     [31:0] n42918;
wire     [31:0] n42919;
wire     [31:0] n42920;
wire     [31:0] n42921;
wire     [31:0] n42922;
wire     [31:0] n42923;
wire     [31:0] n42924;
wire     [31:0] n42925;
wire     [31:0] n42926;
wire     [31:0] n42927;
wire     [31:0] n42928;
wire     [31:0] n42929;
wire     [31:0] n42930;
wire     [31:0] n42931;
wire     [31:0] n42932;
wire     [31:0] n42933;
wire     [31:0] n42934;
wire     [31:0] n42935;
wire     [31:0] n42936;
wire     [31:0] n42937;
wire     [31:0] n42938;
wire     [31:0] n42939;
wire     [31:0] n42940;
wire     [31:0] n42941;
wire     [31:0] n42942;
wire     [31:0] n42943;
wire     [31:0] n42944;
wire     [31:0] n42945;
wire     [31:0] n42946;
wire     [31:0] n42947;
wire     [31:0] n42948;
wire     [31:0] n42949;
wire     [31:0] n42950;
wire     [31:0] n42951;
wire     [31:0] n42952;
wire     [31:0] n42953;
wire     [31:0] n42954;
wire     [31:0] n42955;
wire     [31:0] n42956;
wire     [31:0] n42957;
wire     [31:0] n42958;
wire     [31:0] n42959;
wire     [31:0] n42960;
wire     [31:0] n42961;
wire     [31:0] n42962;
wire     [31:0] n42963;
wire     [31:0] n42964;
wire     [31:0] n42965;
wire     [31:0] n42966;
wire     [31:0] n42967;
wire     [31:0] n42968;
wire     [31:0] n42969;
wire     [31:0] n42970;
wire     [31:0] n42971;
wire     [31:0] n42972;
wire     [31:0] n42973;
wire     [31:0] n42974;
wire     [31:0] n42975;
wire     [31:0] n42976;
wire     [31:0] n42977;
wire     [31:0] n42978;
wire     [31:0] n42979;
wire     [31:0] n42980;
wire     [31:0] n42981;
wire     [31:0] n42982;
wire     [31:0] n42983;
wire     [31:0] n42984;
wire     [31:0] n42985;
wire     [31:0] n42986;
wire     [31:0] n42987;
wire     [31:0] n42988;
wire     [31:0] n42989;
wire     [31:0] n42990;
wire     [31:0] n42991;
wire     [31:0] n42992;
wire     [31:0] n42993;
wire     [31:0] n42994;
wire     [31:0] n42995;
wire     [31:0] n42996;
wire     [31:0] n42997;
wire     [31:0] n42998;
wire     [31:0] n42999;
wire     [31:0] n43000;
wire     [31:0] n43001;
wire     [31:0] n43002;
wire     [31:0] n43003;
wire     [31:0] n43004;
wire     [31:0] n43005;
wire     [31:0] n43006;
wire     [31:0] n43007;
wire     [31:0] n43008;
wire     [31:0] n43009;
wire     [31:0] n43010;
wire     [31:0] n43011;
wire     [31:0] n43012;
wire     [31:0] n43013;
wire     [31:0] n43014;
wire     [31:0] n43015;
wire     [31:0] n43016;
wire     [31:0] n43017;
wire     [31:0] n43018;
wire     [31:0] n43019;
wire     [31:0] n43020;
wire     [31:0] n43021;
wire     [31:0] n43022;
wire     [31:0] n43023;
wire     [31:0] n43024;
wire     [31:0] n43025;
wire     [31:0] n43026;
wire     [31:0] n43027;
wire     [31:0] n43028;
wire     [31:0] n43029;
wire     [31:0] n43030;
wire     [31:0] n43031;
wire     [31:0] n43032;
wire     [31:0] n43033;
wire     [31:0] n43034;
wire     [31:0] n43035;
wire     [31:0] n43036;
wire     [31:0] n43037;
wire     [31:0] n43038;
wire     [31:0] n43039;
wire     [31:0] n43040;
wire     [31:0] n43041;
wire     [31:0] n43042;
wire     [31:0] n43043;
wire     [31:0] n43044;
wire     [31:0] n43045;
wire     [31:0] n43046;
wire     [31:0] n43047;
wire     [31:0] n43048;
wire     [31:0] n43049;
wire     [31:0] n43050;
wire     [31:0] n43051;
wire     [31:0] n43052;
wire     [31:0] n43053;
wire     [31:0] n43054;
wire     [31:0] n43055;
wire     [31:0] n43056;
wire     [31:0] n43057;
wire     [31:0] n43058;
wire     [31:0] n43059;
wire     [31:0] n43060;
wire     [31:0] n43061;
wire     [31:0] n43062;
wire     [31:0] n43063;
wire     [31:0] n43064;
wire     [31:0] n43065;
wire     [31:0] n43066;
wire     [31:0] n43067;
wire     [31:0] n43068;
wire     [31:0] n43069;
wire     [31:0] n43070;
wire     [31:0] n43071;
wire     [31:0] n43072;
wire     [31:0] n43073;
wire     [31:0] n43074;
wire     [31:0] n43075;
wire     [31:0] n43076;
wire     [31:0] n43077;
wire     [31:0] n43078;
wire     [31:0] n43079;
wire     [31:0] n43080;
wire     [31:0] n43081;
wire     [31:0] n43082;
wire     [31:0] n43083;
wire     [31:0] n43084;
wire     [31:0] n43085;
wire     [31:0] n43086;
wire     [31:0] n43087;
wire     [31:0] n43088;
wire     [31:0] n43089;
wire     [31:0] n43090;
wire     [31:0] n43091;
wire     [31:0] n43092;
wire     [31:0] n43093;
wire     [31:0] n43094;
wire     [31:0] n43095;
wire     [31:0] n43096;
wire     [31:0] n43097;
wire     [31:0] n43098;
wire     [31:0] n43099;
wire     [31:0] n43100;
wire     [31:0] n43101;
wire     [31:0] n43102;
wire     [31:0] n43103;
wire     [31:0] n43104;
wire     [31:0] n43105;
wire     [31:0] n43106;
wire     [31:0] n43107;
wire     [31:0] n43108;
wire     [31:0] n43109;
wire     [31:0] n43110;
wire     [31:0] n43111;
wire     [31:0] n43112;
wire     [31:0] n43113;
wire     [31:0] n43114;
wire     [31:0] n43115;
wire     [31:0] n43116;
wire     [31:0] n43117;
wire     [31:0] n43118;
wire     [31:0] n43119;
wire     [31:0] n43120;
wire     [31:0] n43121;
wire     [31:0] n43122;
wire     [31:0] n43123;
wire     [31:0] n43124;
wire     [31:0] n43125;
wire     [31:0] n43126;
wire     [31:0] n43127;
wire     [31:0] n43128;
wire     [31:0] n43129;
wire     [31:0] n43130;
wire     [31:0] n43131;
wire     [31:0] n43132;
wire     [31:0] n43133;
wire     [31:0] n43134;
wire     [31:0] n43135;
wire     [31:0] n43136;
wire     [31:0] n43137;
wire     [31:0] n43138;
wire     [31:0] n43139;
wire     [31:0] n43140;
wire     [31:0] n43141;
wire     [31:0] n43142;
wire     [31:0] n43143;
wire     [31:0] n43144;
wire     [31:0] n43145;
wire     [31:0] n43146;
wire     [31:0] n43147;
wire     [31:0] n43148;
wire     [31:0] n43149;
wire     [31:0] n43150;
wire     [31:0] n43151;
wire     [31:0] n43152;
wire     [31:0] n43153;
wire     [31:0] n43154;
wire     [31:0] n43155;
wire     [31:0] n43156;
wire     [31:0] n43157;
wire     [31:0] n43158;
wire     [31:0] n43159;
wire     [31:0] n43160;
wire     [31:0] n43161;
wire     [31:0] n43162;
wire     [31:0] n43163;
wire     [31:0] n43164;
wire     [31:0] n43165;
wire     [31:0] n43166;
wire     [31:0] n43167;
wire     [31:0] n43168;
wire     [31:0] n43169;
wire     [31:0] n43170;
wire     [31:0] n43171;
wire     [31:0] n43172;
wire     [31:0] n43173;
wire     [31:0] n43174;
wire     [31:0] n43175;
wire     [31:0] n43176;
wire     [31:0] n43177;
wire     [31:0] n43178;
wire     [31:0] n43179;
wire     [31:0] n43180;
wire     [31:0] n43181;
wire     [31:0] n43182;
wire     [31:0] n43183;
wire     [31:0] n43184;
wire     [31:0] n43185;
wire     [31:0] n43186;
wire     [31:0] n43187;
wire     [31:0] n43188;
wire     [31:0] n43189;
wire     [31:0] n43190;
wire     [31:0] n43191;
wire     [31:0] n43192;
wire     [31:0] n43193;
wire     [31:0] n43194;
wire     [31:0] n43195;
wire     [31:0] n43196;
wire     [31:0] n43197;
wire     [31:0] n43198;
wire     [31:0] n43199;
wire     [31:0] n43200;
wire     [31:0] n43201;
wire     [31:0] n43202;
wire     [31:0] n43203;
wire     [31:0] n43204;
wire     [31:0] n43205;
wire     [31:0] n43206;
wire     [31:0] n43207;
wire     [31:0] n43208;
wire     [31:0] n43209;
wire     [31:0] n43210;
wire     [31:0] n43211;
wire     [31:0] n43212;
wire     [31:0] n43213;
wire     [31:0] n43214;
wire     [31:0] n43215;
wire     [31:0] n43216;
wire     [31:0] n43217;
wire     [31:0] n43218;
wire     [31:0] n43219;
wire     [31:0] n43220;
wire     [31:0] n43221;
wire     [31:0] n43222;
wire     [31:0] n43223;
wire     [31:0] n43224;
wire     [31:0] n43225;
wire     [31:0] n43226;
wire     [31:0] n43227;
wire     [31:0] n43228;
wire     [31:0] n43229;
wire     [31:0] n43230;
wire     [31:0] n43231;
wire     [31:0] n43232;
wire     [31:0] n43233;
wire     [31:0] n43234;
wire     [31:0] n43235;
wire     [31:0] n43236;
wire     [31:0] n43237;
wire     [31:0] n43238;
wire     [31:0] n43239;
wire     [31:0] n43240;
wire     [31:0] n43241;
wire     [31:0] n43242;
wire     [31:0] n43243;
wire     [31:0] n43244;
wire     [31:0] n43245;
wire     [31:0] n43246;
wire     [31:0] n43247;
wire     [31:0] n43248;
wire     [31:0] n43249;
wire     [31:0] n43250;
wire     [31:0] n43251;
wire     [31:0] n43252;
wire     [31:0] n43253;
wire     [31:0] n43254;
wire     [31:0] n43255;
wire     [31:0] n43256;
wire     [31:0] n43257;
wire     [31:0] n43258;
wire     [31:0] n43259;
wire     [31:0] n43260;
wire     [31:0] n43261;
wire     [31:0] n43262;
wire     [31:0] n43263;
wire     [31:0] n43264;
wire     [31:0] n43265;
wire     [31:0] n43266;
wire     [31:0] n43267;
wire     [31:0] n43268;
wire     [31:0] n43269;
wire     [31:0] n43270;
wire     [31:0] n43271;
wire     [31:0] n43272;
wire     [31:0] n43273;
wire     [31:0] n43274;
wire     [31:0] n43275;
wire     [31:0] n43276;
wire     [31:0] n43277;
wire     [31:0] n43278;
wire     [31:0] n43279;
wire     [31:0] n43280;
wire     [31:0] n43281;
wire     [31:0] n43282;
wire     [31:0] n43283;
wire     [31:0] n43284;
wire     [31:0] n43285;
wire     [31:0] n43286;
wire     [31:0] n43287;
wire     [31:0] n43288;
wire     [31:0] n43289;
wire     [31:0] n43290;
wire     [31:0] n43291;
wire     [31:0] n43292;
wire     [31:0] n43293;
wire     [31:0] n43294;
wire     [31:0] n43295;
wire     [31:0] n43296;
wire     [31:0] n43297;
wire     [31:0] n43298;
wire     [31:0] n43299;
wire     [31:0] n43300;
wire     [31:0] n43301;
wire     [31:0] n43302;
wire     [31:0] n43303;
wire     [31:0] n43304;
wire     [31:0] n43305;
wire     [31:0] n43306;
wire     [31:0] n43307;
wire     [31:0] n43308;
wire     [31:0] n43309;
wire     [31:0] n43310;
wire     [31:0] n43311;
wire     [31:0] n43312;
wire     [31:0] n43313;
wire     [31:0] n43314;
wire     [31:0] n43315;
wire     [31:0] n43316;
wire     [31:0] n43317;
wire     [31:0] n43318;
wire     [31:0] n43319;
wire     [31:0] n43320;
wire     [31:0] n43321;
wire     [31:0] n43322;
wire     [31:0] n43323;
wire     [31:0] n43324;
wire     [31:0] n43325;
wire     [31:0] n43326;
wire     [31:0] n43327;
wire     [31:0] n43328;
wire     [31:0] n43329;
wire     [31:0] n43330;
wire     [31:0] n43331;
wire     [31:0] n43332;
wire     [31:0] n43333;
wire     [31:0] n43334;
wire     [31:0] n43335;
wire     [31:0] n43336;
wire     [31:0] n43337;
wire     [31:0] n43338;
wire     [31:0] n43339;
wire     [31:0] n43340;
wire     [31:0] n43341;
wire     [31:0] n43342;
wire     [31:0] n43343;
wire     [31:0] n43344;
wire     [31:0] n43345;
wire     [31:0] n43346;
wire     [31:0] n43347;
wire     [31:0] n43348;
wire     [31:0] n43349;
wire     [31:0] n43350;
wire     [31:0] n43351;
wire     [31:0] n43352;
wire     [31:0] n43353;
wire     [31:0] n43354;
wire     [31:0] n43355;
wire     [31:0] n43356;
wire     [31:0] n43357;
wire     [31:0] n43358;
wire     [31:0] n43359;
wire     [31:0] n43360;
wire     [31:0] n43361;
wire     [31:0] n43362;
wire     [31:0] n43363;
wire     [31:0] n43364;
wire     [31:0] n43365;
wire     [31:0] n43366;
wire     [31:0] n43367;
wire     [31:0] n43368;
wire     [31:0] n43369;
wire     [31:0] n43370;
wire     [31:0] n43371;
wire     [31:0] n43372;
wire     [31:0] n43373;
wire     [31:0] n43374;
wire     [31:0] n43375;
wire     [31:0] n43376;
wire     [31:0] n43377;
wire     [31:0] n43378;
wire     [31:0] n43379;
wire     [31:0] n43380;
wire     [31:0] n43381;
wire     [31:0] n43382;
wire     [31:0] n43383;
wire     [31:0] n43384;
wire     [31:0] n43385;
wire     [31:0] n43386;
wire     [31:0] n43387;
wire     [31:0] n43388;
wire     [31:0] n43389;
wire     [31:0] n43390;
wire     [31:0] n43391;
wire     [31:0] n43392;
wire     [31:0] n43393;
wire     [31:0] n43394;
wire     [31:0] n43395;
wire     [31:0] n43396;
wire     [31:0] n43397;
wire     [31:0] n43398;
wire     [31:0] n43399;
wire     [31:0] n43400;
wire     [31:0] n43401;
wire     [31:0] n43402;
wire     [31:0] n43403;
wire     [31:0] n43404;
wire     [31:0] n43405;
wire     [31:0] n43406;
wire     [31:0] n43407;
wire     [31:0] n43408;
wire     [31:0] n43409;
wire     [31:0] n43410;
wire     [31:0] n43411;
wire     [31:0] n43412;
wire     [31:0] n43413;
wire     [31:0] n43414;
wire     [31:0] n43415;
wire     [31:0] n43416;
wire     [31:0] n43417;
wire     [31:0] n43418;
wire     [31:0] n43419;
wire     [31:0] n43420;
wire     [31:0] n43421;
wire     [31:0] n43422;
wire     [31:0] n43423;
wire     [31:0] n43424;
wire     [31:0] n43425;
wire     [31:0] n43426;
wire     [31:0] n43427;
wire     [31:0] n43428;
wire     [31:0] n43429;
wire     [31:0] n43430;
wire     [31:0] n43431;
wire     [31:0] n43432;
wire     [31:0] n43433;
wire     [31:0] n43434;
wire     [31:0] n43435;
wire     [31:0] n43436;
wire     [31:0] n43437;
wire     [31:0] n43438;
wire     [31:0] n43439;
wire     [31:0] n43440;
wire     [31:0] n43441;
wire     [31:0] n43442;
wire     [31:0] n43443;
wire     [31:0] n43444;
wire     [31:0] n43445;
wire     [31:0] n43446;
wire     [31:0] n43447;
wire     [31:0] n43448;
wire     [31:0] n43449;
wire     [31:0] n43450;
wire     [31:0] n43451;
wire     [31:0] n43452;
wire     [31:0] n43453;
wire     [31:0] n43454;
wire     [31:0] n43455;
wire     [31:0] n43456;
wire     [31:0] n43457;
wire     [31:0] n43458;
wire     [31:0] n43459;
wire     [31:0] n43460;
wire     [31:0] n43461;
wire     [31:0] n43462;
wire     [31:0] n43463;
wire     [31:0] n43464;
wire     [31:0] n43465;
wire     [31:0] n43466;
wire     [31:0] n43467;
wire     [31:0] n43468;
wire     [31:0] n43469;
wire     [31:0] n43470;
wire     [31:0] n43471;
wire     [31:0] n43472;
wire     [31:0] n43473;
wire     [31:0] n43474;
wire     [31:0] n43475;
wire     [31:0] n43476;
wire     [31:0] n43477;
wire     [31:0] n43478;
wire     [31:0] n43479;
wire     [31:0] n43480;
wire     [31:0] n43481;
wire     [31:0] n43482;
wire     [31:0] n43483;
wire     [31:0] n43484;
wire     [31:0] n43485;
wire     [31:0] n43486;
wire     [31:0] n43487;
wire     [31:0] n43488;
wire     [31:0] n43489;
wire     [31:0] n43490;
wire     [31:0] n43491;
wire     [31:0] n43492;
wire     [31:0] n43493;
wire     [31:0] n43494;
wire     [31:0] n43495;
wire     [31:0] n43496;
wire     [31:0] n43497;
wire     [31:0] n43498;
wire     [31:0] n43499;
wire     [31:0] n43500;
wire     [31:0] n43501;
wire     [31:0] n43502;
wire     [31:0] n43503;
wire     [31:0] n43504;
wire     [31:0] n43505;
wire     [31:0] n43506;
wire     [31:0] n43507;
wire     [31:0] n43508;
wire     [31:0] n43509;
wire     [31:0] n43510;
wire     [31:0] n43511;
wire     [31:0] n43512;
wire     [31:0] n43513;
wire     [31:0] n43514;
wire     [31:0] n43515;
wire     [31:0] n43516;
wire     [31:0] n43517;
wire     [31:0] n43518;
wire     [31:0] n43519;
wire     [31:0] n43520;
wire     [31:0] n43521;
wire     [31:0] n43522;
wire     [31:0] n43523;
wire     [31:0] n43524;
wire     [31:0] n43525;
wire     [31:0] n43526;
wire     [31:0] n43527;
wire     [31:0] n43528;
wire     [31:0] n43529;
wire     [31:0] n43530;
wire     [31:0] n43531;
wire     [31:0] n43532;
wire     [31:0] n43533;
wire     [31:0] n43534;
wire     [31:0] n43535;
wire     [31:0] n43536;
wire     [31:0] n43537;
wire     [31:0] n43538;
wire     [31:0] n43539;
wire     [31:0] n43540;
wire     [31:0] n43541;
wire     [31:0] n43542;
wire     [31:0] n43543;
wire     [31:0] n43544;
wire     [31:0] n43545;
wire     [31:0] n43546;
wire     [31:0] n43547;
wire     [31:0] n43548;
wire     [31:0] n43549;
wire     [31:0] n43550;
wire     [31:0] n43551;
wire     [31:0] n43552;
wire     [31:0] n43553;
wire     [31:0] n43554;
wire     [31:0] n43555;
wire     [31:0] n43556;
wire     [31:0] n43557;
wire     [31:0] n43558;
wire     [31:0] n43559;
wire     [31:0] n43560;
wire     [31:0] n43561;
wire     [31:0] n43562;
wire     [31:0] n43563;
wire     [31:0] n43564;
wire     [31:0] n43565;
wire     [31:0] n43566;
wire     [31:0] n43567;
wire     [31:0] n43568;
wire     [31:0] n43569;
wire     [31:0] n43570;
wire     [31:0] n43571;
wire     [31:0] n43572;
wire     [31:0] n43573;
wire     [31:0] n43574;
wire     [31:0] n43575;
wire     [31:0] n43576;
wire     [31:0] n43577;
wire     [31:0] n43578;
wire     [31:0] n43579;
wire     [31:0] n43580;
wire     [31:0] n43581;
wire     [31:0] n43582;
wire     [31:0] n43583;
wire     [31:0] n43584;
wire     [31:0] n43585;
wire     [31:0] n43586;
wire     [31:0] n43587;
wire     [31:0] n43588;
wire     [31:0] n43589;
wire     [31:0] n43590;
wire     [31:0] n43591;
wire     [31:0] n43592;
wire     [31:0] n43593;
wire     [31:0] n43594;
wire     [31:0] n43595;
wire     [31:0] n43596;
wire     [31:0] n43597;
wire     [31:0] n43598;
wire     [31:0] n43599;
wire     [31:0] n43600;
wire     [31:0] n43601;
wire     [31:0] n43602;
wire     [31:0] n43603;
wire     [31:0] n43604;
wire     [31:0] n43605;
wire     [31:0] n43606;
wire     [31:0] n43607;
wire     [31:0] n43608;
wire     [31:0] n43609;
wire     [31:0] n43610;
wire     [31:0] n43611;
wire     [31:0] n43612;
wire     [31:0] n43613;
wire     [31:0] n43614;
wire     [31:0] n43615;
wire     [31:0] n43616;
wire     [31:0] n43617;
wire     [31:0] n43618;
wire     [31:0] n43619;
wire     [31:0] n43620;
wire     [31:0] n43621;
wire     [31:0] n43622;
wire     [31:0] n43623;
wire     [31:0] n43624;
wire     [31:0] n43625;
wire     [31:0] n43626;
wire     [31:0] n43627;
wire     [31:0] n43628;
wire     [31:0] n43629;
wire     [31:0] n43630;
wire     [31:0] n43631;
wire     [31:0] n43632;
wire     [31:0] n43633;
wire     [31:0] n43634;
wire     [31:0] n43635;
wire     [31:0] n43636;
wire     [31:0] n43637;
wire     [31:0] n43638;
wire     [31:0] n43639;
wire     [31:0] n43640;
wire     [31:0] n43641;
wire     [31:0] n43642;
wire     [31:0] n43643;
wire     [31:0] n43644;
wire     [31:0] n43645;
wire     [31:0] n43646;
wire     [31:0] n43647;
wire     [31:0] n43648;
wire     [31:0] n43649;
wire     [31:0] n43650;
wire     [31:0] n43651;
wire     [31:0] n43652;
wire     [31:0] n43653;
wire     [31:0] n43654;
wire     [31:0] n43655;
wire     [31:0] n43656;
wire     [31:0] n43657;
wire     [31:0] n43658;
wire     [31:0] n43659;
wire     [31:0] n43660;
wire     [31:0] n43661;
wire     [31:0] n43662;
wire     [31:0] n43663;
wire     [31:0] n43664;
wire     [31:0] n43665;
wire     [31:0] n43666;
wire     [31:0] n43667;
wire     [31:0] n43668;
wire     [31:0] n43669;
wire     [31:0] n43670;
wire     [31:0] n43671;
wire     [31:0] n43672;
wire     [31:0] n43673;
wire     [31:0] n43674;
wire     [31:0] n43675;
wire     [31:0] n43676;
wire     [31:0] n43677;
wire     [31:0] n43678;
wire     [31:0] n43679;
wire     [31:0] n43680;
wire     [31:0] n43681;
wire     [31:0] n43682;
wire     [31:0] n43683;
wire     [31:0] n43684;
wire     [31:0] n43685;
wire     [31:0] n43686;
wire     [31:0] n43687;
wire     [31:0] n43688;
wire     [31:0] n43689;
wire     [31:0] n43690;
wire     [31:0] n43691;
wire     [31:0] n43692;
wire     [31:0] n43693;
wire     [31:0] n43694;
wire     [31:0] n43695;
wire     [31:0] n43696;
wire     [31:0] n43697;
wire     [31:0] n43698;
wire     [31:0] n43699;
wire     [31:0] n43700;
wire     [31:0] n43701;
wire     [31:0] n43702;
wire     [31:0] n43703;
wire     [31:0] n43704;
wire     [31:0] n43705;
wire     [31:0] n43706;
wire     [31:0] n43707;
wire     [31:0] n43708;
wire     [31:0] n43709;
wire     [31:0] n43710;
wire     [31:0] n43711;
wire     [31:0] n43712;
wire     [31:0] n43713;
wire     [31:0] n43714;
wire     [31:0] n43715;
wire     [31:0] n43716;
wire     [31:0] n43717;
wire     [31:0] n43718;
wire     [31:0] n43719;
wire     [31:0] n43720;
wire     [31:0] n43721;
wire     [31:0] n43722;
wire     [31:0] n43723;
wire     [31:0] n43724;
wire     [31:0] n43725;
wire     [31:0] n43726;
wire     [31:0] n43727;
wire     [31:0] n43728;
wire     [31:0] n43729;
wire     [31:0] n43730;
wire     [31:0] n43731;
wire     [31:0] n43732;
wire     [31:0] n43733;
wire     [31:0] n43734;
wire     [31:0] n43735;
wire     [31:0] n43736;
wire     [31:0] n43737;
wire     [31:0] n43738;
wire     [31:0] n43739;
wire     [31:0] n43740;
wire     [31:0] n43741;
wire     [31:0] n43742;
wire     [31:0] n43743;
wire     [31:0] n43744;
wire     [31:0] n43745;
wire     [31:0] n43746;
wire     [31:0] n43747;
wire     [31:0] n43748;
wire     [31:0] n43749;
wire     [31:0] n43750;
wire     [31:0] n43751;
wire     [31:0] n43752;
wire     [31:0] n43753;
wire     [31:0] n43754;
wire     [31:0] n43755;
wire     [31:0] n43756;
wire     [31:0] n43757;
wire     [31:0] n43758;
wire     [31:0] n43759;
wire     [31:0] n43760;
wire     [31:0] n43761;
wire     [31:0] n43762;
wire     [31:0] n43763;
wire     [31:0] n43764;
wire     [31:0] n43765;
wire     [31:0] n43766;
wire     [31:0] n43767;
wire     [31:0] n43768;
wire     [31:0] n43769;
wire     [31:0] n43770;
wire     [31:0] n43771;
wire     [31:0] n43772;
wire     [31:0] n43773;
wire     [31:0] n43774;
wire     [31:0] n43775;
wire     [31:0] n43776;
wire     [31:0] n43777;
wire     [31:0] n43778;
wire     [31:0] n43779;
wire     [31:0] n43780;
wire     [31:0] n43781;
wire     [31:0] n43782;
wire     [31:0] n43783;
wire     [31:0] n43784;
wire     [31:0] n43785;
wire     [31:0] n43786;
wire     [31:0] n43787;
wire     [31:0] n43788;
wire     [31:0] n43789;
wire     [31:0] n43790;
wire     [31:0] n43791;
wire     [31:0] n43792;
wire     [31:0] n43793;
wire     [31:0] n43794;
wire     [31:0] n43795;
wire     [31:0] n43796;
wire     [31:0] n43797;
wire     [31:0] n43798;
wire     [31:0] n43799;
wire     [31:0] n43800;
wire     [31:0] n43801;
wire     [31:0] n43802;
wire     [31:0] n43803;
wire     [31:0] n43804;
wire     [31:0] n43805;
wire     [31:0] n43806;
wire     [31:0] n43807;
wire     [31:0] n43808;
wire     [31:0] n43809;
wire     [31:0] n43810;
wire     [31:0] n43811;
wire     [31:0] n43812;
wire     [31:0] n43813;
wire     [31:0] n43814;
wire     [31:0] n43815;
wire     [31:0] n43816;
wire     [31:0] n43817;
wire     [31:0] n43818;
wire     [31:0] n43819;
wire     [31:0] n43820;
wire     [31:0] n43821;
wire     [31:0] n43822;
wire     [31:0] n43823;
wire     [31:0] n43824;
wire     [31:0] n43825;
wire     [31:0] n43826;
wire     [31:0] n43827;
wire     [31:0] n43828;
wire     [31:0] n43829;
wire     [31:0] n43830;
wire     [31:0] n43831;
wire     [31:0] n43832;
wire     [31:0] n43833;
wire     [31:0] n43834;
wire     [31:0] n43835;
wire     [31:0] n43836;
wire     [31:0] n43837;
wire     [31:0] n43838;
wire     [31:0] n43839;
wire     [31:0] n43840;
wire     [31:0] n43841;
wire     [31:0] n43842;
wire     [31:0] n43843;
wire     [31:0] n43844;
wire     [31:0] n43845;
wire     [31:0] n43846;
wire     [31:0] n43847;
wire     [31:0] n43848;
wire     [31:0] n43849;
wire     [31:0] n43850;
wire     [31:0] n43851;
wire     [31:0] n43852;
wire     [31:0] n43853;
wire     [31:0] n43854;
wire     [31:0] n43855;
wire     [31:0] n43856;
wire     [31:0] n43857;
wire     [31:0] n43858;
wire     [31:0] n43859;
wire     [31:0] n43860;
wire     [31:0] n43861;
wire     [31:0] n43862;
wire     [31:0] n43863;
wire     [31:0] n43864;
wire     [31:0] n43865;
wire     [31:0] n43866;
wire     [31:0] n43867;
wire     [31:0] n43868;
wire     [31:0] n43869;
wire     [31:0] n43870;
wire     [31:0] n43871;
wire     [31:0] n43872;
wire     [31:0] n43873;
wire     [31:0] n43874;
wire     [31:0] n43875;
wire     [31:0] n43876;
wire     [31:0] n43877;
wire     [31:0] n43878;
wire     [31:0] n43879;
wire     [31:0] n43880;
wire     [31:0] n43881;
wire     [31:0] n43882;
wire     [31:0] n43883;
wire     [31:0] n43884;
wire     [31:0] n43885;
wire     [31:0] n43886;
wire     [31:0] n43887;
wire     [31:0] n43888;
wire     [31:0] n43889;
wire     [31:0] n43890;
wire     [31:0] n43891;
wire     [31:0] n43892;
wire     [31:0] n43893;
wire     [31:0] n43894;
wire     [31:0] n43895;
wire     [31:0] n43896;
wire     [31:0] n43897;
wire     [31:0] n43898;
wire     [31:0] n43899;
wire     [31:0] n43900;
wire     [31:0] n43901;
wire     [31:0] n43902;
wire     [31:0] n43903;
wire     [31:0] n43904;
wire     [31:0] n43905;
wire     [31:0] n43906;
wire     [31:0] n43907;
wire     [31:0] n43908;
wire     [31:0] n43909;
wire     [31:0] n43910;
wire     [31:0] n43911;
wire     [31:0] n43912;
wire     [31:0] n43913;
wire     [31:0] n43914;
wire     [31:0] n43915;
wire     [31:0] n43916;
wire     [31:0] n43917;
wire     [31:0] n43918;
wire     [31:0] n43919;
wire     [31:0] n43920;
wire     [31:0] n43921;
wire     [31:0] n43922;
wire     [31:0] n43923;
wire     [31:0] n43924;
wire     [31:0] n43925;
wire     [31:0] n43926;
wire     [31:0] n43927;
wire     [31:0] n43928;
wire     [31:0] n43929;
wire     [31:0] n43930;
wire     [31:0] n43931;
wire     [31:0] n43932;
wire     [31:0] n43933;
wire     [31:0] n43934;
wire     [31:0] n43935;
wire     [31:0] n43936;
wire     [31:0] n43937;
wire     [31:0] n43938;
wire     [31:0] n43939;
wire     [31:0] n43940;
wire     [31:0] n43941;
wire     [31:0] n43942;
wire     [31:0] n43943;
wire     [31:0] n43944;
wire     [31:0] n43945;
wire     [31:0] n43946;
wire     [31:0] n43947;
wire     [31:0] n43948;
wire     [31:0] n43949;
wire     [31:0] n43950;
wire     [31:0] n43951;
wire     [31:0] n43952;
wire     [31:0] n43953;
wire     [31:0] n43954;
wire     [31:0] n43955;
wire     [31:0] n43956;
wire     [31:0] n43957;
wire     [31:0] n43958;
wire     [31:0] n43959;
wire     [31:0] n43960;
wire     [31:0] n43961;
wire     [31:0] n43962;
wire     [31:0] n43963;
wire     [31:0] n43964;
wire     [31:0] n43965;
wire     [31:0] n43966;
wire     [31:0] n43967;
wire     [31:0] n43968;
wire     [31:0] n43969;
wire     [31:0] n43970;
wire     [31:0] n43971;
wire     [31:0] n43972;
wire     [31:0] n43973;
wire     [31:0] n43974;
wire     [31:0] n43975;
wire     [31:0] n43976;
wire     [31:0] n43977;
wire     [31:0] n43978;
wire     [31:0] n43979;
wire     [31:0] n43980;
wire     [31:0] n43981;
wire     [31:0] n43982;
wire     [31:0] n43983;
wire     [31:0] n43984;
wire     [31:0] n43985;
wire     [31:0] n43986;
wire     [31:0] n43987;
wire     [31:0] n43988;
wire     [31:0] n43989;
wire     [31:0] n43990;
wire     [31:0] n43991;
wire     [31:0] n43992;
wire     [31:0] n43993;
wire     [31:0] n43994;
wire     [31:0] n43995;
wire     [31:0] n43996;
wire     [31:0] n43997;
wire     [31:0] n43998;
wire     [31:0] n43999;
wire     [31:0] n44000;
wire     [31:0] n44001;
wire     [31:0] n44002;
wire     [31:0] n44003;
wire     [31:0] n44004;
wire     [31:0] n44005;
wire     [31:0] n44006;
wire     [31:0] n44007;
wire     [31:0] n44008;
wire     [31:0] n44009;
wire     [31:0] n44010;
wire     [31:0] n44011;
wire     [31:0] n44012;
wire     [31:0] n44013;
wire     [31:0] n44014;
wire     [31:0] n44015;
wire     [31:0] n44016;
wire     [31:0] n44017;
wire     [31:0] n44018;
wire     [31:0] n44019;
wire     [31:0] n44020;
wire     [31:0] n44021;
wire     [31:0] n44022;
wire     [31:0] n44023;
wire     [31:0] n44024;
wire     [31:0] n44025;
wire     [31:0] n44026;
wire     [31:0] n44027;
wire     [31:0] n44028;
wire     [31:0] n44029;
wire     [31:0] n44030;
wire     [31:0] n44031;
wire     [31:0] n44032;
wire     [31:0] n44033;
wire     [31:0] n44034;
wire     [31:0] n44035;
wire     [31:0] n44036;
wire     [31:0] n44037;
wire     [31:0] n44038;
wire     [31:0] n44039;
wire     [31:0] n44040;
wire     [31:0] n44041;
wire     [31:0] n44042;
wire     [31:0] n44043;
wire     [31:0] n44044;
wire     [31:0] n44045;
wire     [31:0] n44046;
wire     [31:0] n44047;
wire     [31:0] n44048;
wire     [31:0] n44049;
wire     [31:0] n44050;
wire     [31:0] n44051;
wire     [31:0] n44052;
wire     [31:0] n44053;
wire     [31:0] n44054;
wire     [31:0] n44055;
wire     [31:0] n44056;
wire     [31:0] n44057;
wire     [31:0] n44058;
wire     [31:0] n44059;
wire     [31:0] n44060;
wire     [31:0] n44061;
wire     [31:0] n44062;
wire     [31:0] n44063;
wire     [31:0] n44064;
wire     [31:0] n44065;
wire     [31:0] n44066;
wire     [31:0] n44067;
wire     [31:0] n44068;
wire     [31:0] n44069;
wire     [31:0] n44070;
wire     [31:0] n44071;
wire     [31:0] n44072;
wire     [31:0] n44073;
wire     [31:0] n44074;
wire     [31:0] n44075;
wire     [31:0] n44076;
wire     [31:0] n44077;
wire     [31:0] n44078;
wire     [31:0] n44079;
wire     [31:0] n44080;
wire     [31:0] n44081;
wire     [31:0] n44082;
wire     [31:0] n44083;
wire     [31:0] n44084;
wire     [31:0] n44085;
wire     [31:0] n44086;
wire     [31:0] n44087;
wire     [31:0] n44088;
wire     [31:0] n44089;
wire     [31:0] n44090;
wire     [31:0] n44091;
wire     [31:0] n44092;
wire     [31:0] n44093;
wire     [31:0] n44094;
wire     [31:0] n44095;
wire     [31:0] n44096;
wire     [31:0] n44097;
wire     [31:0] n44098;
wire     [31:0] n44099;
wire     [31:0] n44100;
wire     [31:0] n44101;
wire     [31:0] n44102;
wire     [31:0] n44103;
wire     [31:0] n44104;
wire     [31:0] n44105;
wire     [31:0] n44106;
wire     [31:0] n44107;
wire     [31:0] n44108;
wire     [31:0] n44109;
wire     [31:0] n44110;
wire     [31:0] n44111;
wire     [31:0] n44112;
wire     [31:0] n44113;
wire     [31:0] n44114;
wire     [31:0] n44115;
wire     [31:0] n44116;
wire     [31:0] n44117;
wire     [31:0] n44118;
wire     [31:0] n44119;
wire     [31:0] n44120;
wire     [31:0] n44121;
wire     [31:0] n44122;
wire     [31:0] n44123;
wire     [31:0] n44124;
wire     [31:0] n44125;
wire     [31:0] n44126;
wire     [31:0] n44127;
wire     [31:0] n44128;
wire     [31:0] n44129;
wire     [31:0] n44130;
wire     [31:0] n44131;
wire     [31:0] n44132;
wire     [31:0] n44133;
wire     [31:0] n44134;
wire     [31:0] n44135;
wire     [31:0] n44136;
wire     [31:0] n44137;
wire     [31:0] n44138;
wire     [31:0] n44139;
wire     [31:0] n44140;
wire     [31:0] n44141;
wire     [31:0] n44142;
wire     [31:0] n44143;
wire     [31:0] n44144;
wire     [31:0] n44145;
wire     [31:0] n44146;
wire     [31:0] n44147;
wire     [31:0] n44148;
wire     [31:0] n44149;
wire     [31:0] n44150;
wire     [31:0] n44151;
wire     [31:0] n44152;
wire     [31:0] n44153;
wire     [31:0] n44154;
wire     [31:0] n44155;
wire     [31:0] n44156;
wire     [31:0] n44157;
wire     [31:0] n44158;
wire     [31:0] n44159;
wire     [31:0] n44160;
wire     [31:0] n44161;
wire     [31:0] n44162;
wire     [31:0] n44163;
wire     [31:0] n44164;
wire     [31:0] n44165;
wire     [31:0] n44166;
wire     [31:0] n44167;
wire     [31:0] n44168;
wire     [31:0] n44169;
wire     [31:0] n44170;
wire     [31:0] n44171;
wire     [31:0] n44172;
wire     [31:0] n44173;
wire     [31:0] n44174;
wire     [31:0] n44175;
wire     [31:0] n44176;
wire     [31:0] n44177;
wire     [31:0] n44178;
wire     [31:0] n44179;
wire     [31:0] n44180;
wire     [31:0] n44181;
wire     [31:0] n44182;
wire     [31:0] n44183;
wire     [31:0] n44184;
wire     [31:0] n44185;
wire     [31:0] n44186;
wire     [31:0] n44187;
wire     [31:0] n44188;
wire     [31:0] n44189;
wire     [31:0] n44190;
wire     [31:0] n44191;
wire     [31:0] n44192;
wire     [31:0] n44193;
wire     [31:0] n44194;
wire     [31:0] n44195;
wire     [31:0] n44196;
wire     [31:0] n44197;
wire     [31:0] n44198;
wire     [31:0] n44199;
wire     [31:0] n44200;
wire     [31:0] n44201;
wire     [31:0] n44202;
wire     [31:0] n44203;
wire     [31:0] n44204;
wire     [31:0] n44205;
wire     [31:0] n44206;
wire     [31:0] n44207;
wire     [31:0] n44208;
wire     [31:0] n44209;
wire     [31:0] n44210;
wire     [31:0] n44211;
wire     [31:0] n44212;
wire     [31:0] n44213;
wire     [31:0] n44214;
wire     [31:0] n44215;
wire     [31:0] n44216;
wire     [31:0] n44217;
wire     [31:0] n44218;
wire     [31:0] n44219;
wire     [31:0] n44220;
wire     [31:0] n44221;
wire     [31:0] n44222;
wire     [31:0] n44223;
wire     [31:0] n44224;
wire     [31:0] n44225;
wire     [31:0] n44226;
wire     [31:0] n44227;
wire     [31:0] n44228;
wire     [31:0] n44229;
wire     [31:0] n44230;
wire     [31:0] n44231;
wire     [31:0] n44232;
wire     [31:0] n44233;
wire     [31:0] n44234;
wire     [31:0] n44235;
wire     [31:0] n44236;
wire     [31:0] n44237;
wire     [31:0] n44238;
wire     [31:0] n44239;
wire     [31:0] n44240;
wire     [31:0] n44241;
wire     [31:0] n44242;
wire     [31:0] n44243;
wire     [31:0] n44244;
wire     [31:0] n44245;
wire     [31:0] n44246;
wire     [31:0] n44247;
wire     [31:0] n44248;
wire     [31:0] n44249;
wire     [31:0] n44250;
wire     [31:0] n44251;
wire     [31:0] n44252;
wire     [31:0] n44253;
wire     [31:0] n44254;
wire     [31:0] n44255;
wire     [31:0] n44256;
wire     [31:0] n44257;
wire     [31:0] n44258;
wire     [31:0] n44259;
wire     [31:0] n44260;
wire     [31:0] n44261;
wire     [31:0] n44262;
wire     [31:0] n44263;
wire     [31:0] n44264;
wire     [31:0] n44265;
wire     [31:0] n44266;
wire     [31:0] n44267;
wire     [31:0] n44268;
wire     [31:0] n44269;
wire     [31:0] n44270;
wire     [31:0] n44271;
wire     [31:0] n44272;
wire     [31:0] n44273;
wire     [31:0] n44274;
wire     [31:0] n44275;
wire     [31:0] n44276;
wire     [31:0] n44277;
wire     [31:0] n44278;
wire     [31:0] n44279;
wire     [31:0] n44280;
wire     [31:0] n44281;
wire     [31:0] n44282;
wire     [31:0] n44283;
wire     [31:0] n44284;
wire     [31:0] n44285;
wire     [31:0] n44286;
wire     [31:0] n44287;
wire     [31:0] n44288;
wire     [31:0] n44289;
wire     [31:0] n44290;
wire     [31:0] n44291;
wire     [31:0] n44292;
wire     [31:0] n44293;
wire     [31:0] n44294;
wire     [31:0] n44295;
wire     [31:0] n44296;
wire     [31:0] n44297;
wire     [31:0] n44298;
wire     [31:0] n44299;
wire     [31:0] n44300;
wire     [31:0] n44301;
wire     [31:0] n44302;
wire     [31:0] n44303;
wire     [31:0] n44304;
wire     [31:0] n44305;
wire     [31:0] n44306;
wire     [31:0] n44307;
wire     [31:0] n44308;
wire     [31:0] n44309;
wire     [31:0] n44310;
wire     [31:0] n44311;
wire     [31:0] n44312;
wire     [31:0] n44313;
wire     [31:0] n44314;
wire     [31:0] n44315;
wire     [31:0] n44316;
wire     [31:0] n44317;
wire     [31:0] n44318;
wire     [31:0] n44319;
wire     [31:0] n44320;
wire     [31:0] n44321;
wire     [31:0] n44322;
wire     [31:0] n44323;
wire     [31:0] n44324;
wire     [31:0] n44325;
wire     [31:0] n44326;
wire     [31:0] n44327;
wire     [31:0] n44328;
wire     [31:0] n44329;
wire     [31:0] n44330;
wire     [31:0] n44331;
wire     [31:0] n44332;
wire     [31:0] n44333;
wire     [31:0] n44334;
wire     [31:0] n44335;
wire     [31:0] n44336;
wire     [31:0] n44337;
wire     [31:0] n44338;
wire     [31:0] n44339;
wire     [31:0] n44340;
wire     [31:0] n44341;
wire     [31:0] n44342;
wire     [31:0] n44343;
wire     [31:0] n44344;
wire     [31:0] n44345;
wire     [31:0] n44346;
wire     [31:0] n44347;
wire     [31:0] n44348;
wire     [31:0] n44349;
wire     [31:0] n44350;
wire     [31:0] n44351;
wire     [31:0] n44352;
wire     [31:0] n44353;
wire     [31:0] n44354;
wire     [31:0] n44355;
wire     [31:0] n44356;
wire     [31:0] n44357;
wire     [31:0] n44358;
wire     [31:0] n44359;
wire     [31:0] n44360;
wire     [31:0] n44361;
wire     [31:0] n44362;
wire     [31:0] n44363;
wire     [31:0] n44364;
wire     [31:0] n44365;
wire     [31:0] n44366;
wire     [31:0] n44367;
wire     [31:0] n44368;
wire     [31:0] n44369;
wire     [31:0] n44370;
wire     [31:0] n44371;
wire     [31:0] n44372;
wire     [31:0] n44373;
wire     [31:0] n44374;
wire     [31:0] n44375;
wire     [31:0] n44376;
wire     [31:0] n44377;
wire     [31:0] n44378;
wire     [31:0] n44379;
wire     [31:0] n44380;
wire     [31:0] n44381;
wire     [31:0] n44382;
wire     [31:0] n44383;
wire     [31:0] n44384;
wire     [31:0] n44385;
wire     [31:0] n44386;
wire     [31:0] n44387;
wire     [31:0] n44388;
wire     [31:0] n44389;
wire     [31:0] n44390;
wire     [31:0] n44391;
wire     [31:0] n44392;
wire     [31:0] n44393;
wire     [31:0] n44394;
wire     [31:0] n44395;
wire     [31:0] n44396;
wire     [31:0] n44397;
wire     [31:0] n44398;
wire     [31:0] n44399;
wire     [31:0] n44400;
wire     [31:0] n44401;
wire     [31:0] n44402;
wire     [31:0] n44403;
wire     [31:0] n44404;
wire     [31:0] n44405;
wire     [31:0] n44406;
wire     [31:0] n44407;
wire     [31:0] n44408;
wire     [31:0] n44409;
wire     [31:0] n44410;
wire     [31:0] n44411;
wire     [31:0] n44412;
wire     [31:0] n44413;
wire     [31:0] n44414;
wire     [31:0] n44415;
wire     [31:0] n44416;
wire     [31:0] n44417;
wire     [31:0] n44418;
wire     [31:0] n44419;
wire     [31:0] n44420;
wire     [31:0] n44421;
wire     [31:0] n44422;
wire     [31:0] n44423;
wire     [31:0] n44424;
wire     [31:0] n44425;
wire     [31:0] n44426;
wire     [31:0] n44427;
wire     [31:0] n44428;
wire     [31:0] n44429;
wire     [31:0] n44430;
wire     [31:0] n44431;
wire     [31:0] n44432;
wire     [31:0] n44433;
wire     [31:0] n44434;
wire     [31:0] n44435;
wire     [31:0] n44436;
wire     [31:0] n44437;
wire     [31:0] n44438;
wire     [31:0] n44439;
wire     [31:0] n44440;
wire     [31:0] n44441;
wire     [31:0] n44442;
wire     [31:0] n44443;
wire     [31:0] n44444;
wire     [31:0] n44445;
wire     [31:0] n44446;
wire     [31:0] n44447;
wire     [31:0] n44448;
wire     [31:0] n44449;
wire     [31:0] n44450;
wire     [31:0] n44451;
wire     [31:0] n44452;
wire     [31:0] n44453;
wire     [31:0] n44454;
wire     [31:0] n44455;
wire     [31:0] n44456;
wire     [31:0] n44457;
wire     [31:0] n44458;
wire     [31:0] n44459;
wire     [31:0] n44460;
wire     [31:0] n44461;
wire     [31:0] n44462;
wire     [31:0] n44463;
wire     [31:0] n44464;
wire     [31:0] n44465;
wire     [31:0] n44466;
wire     [31:0] n44467;
wire     [31:0] n44468;
wire     [31:0] n44469;
wire     [31:0] n44470;
wire     [31:0] n44471;
wire     [31:0] n44472;
wire     [31:0] n44473;
wire     [31:0] n44474;
wire     [31:0] n44475;
wire     [31:0] n44476;
wire     [31:0] n44477;
wire     [31:0] n44478;
wire     [31:0] n44479;
wire     [31:0] n44480;
wire     [31:0] n44481;
wire     [31:0] n44482;
wire     [31:0] n44483;
wire     [31:0] n44484;
wire     [31:0] n44485;
wire     [31:0] n44486;
wire     [31:0] n44487;
wire     [31:0] n44488;
wire     [31:0] n44489;
wire     [31:0] n44490;
wire     [31:0] n44491;
wire     [31:0] n44492;
wire     [31:0] n44493;
wire     [31:0] n44494;
wire     [31:0] n44495;
wire     [31:0] n44496;
wire     [31:0] n44497;
wire     [31:0] n44498;
wire     [31:0] n44499;
wire     [31:0] n44500;
wire     [31:0] n44501;
wire     [31:0] n44502;
wire     [31:0] n44503;
wire     [31:0] n44504;
wire     [31:0] n44505;
wire     [31:0] n44506;
wire     [31:0] n44507;
wire     [31:0] n44508;
wire     [31:0] n44509;
wire     [31:0] n44510;
wire     [31:0] n44511;
wire     [31:0] n44512;
wire     [31:0] n44513;
wire     [31:0] n44514;
wire     [31:0] n44515;
wire     [31:0] n44516;
wire     [31:0] n44517;
wire     [31:0] n44518;
wire     [31:0] n44519;
wire     [31:0] n44520;
wire     [31:0] n44521;
wire     [31:0] n44522;
wire     [31:0] n44523;
wire     [31:0] n44524;
wire     [31:0] n44525;
wire     [31:0] n44526;
wire     [31:0] n44527;
wire     [31:0] n44528;
wire     [31:0] n44529;
wire     [31:0] n44530;
wire     [31:0] n44531;
wire     [31:0] n44532;
wire     [31:0] n44533;
wire     [31:0] n44534;
wire     [31:0] n44535;
wire     [31:0] n44536;
wire     [31:0] n44537;
wire     [31:0] n44538;
wire     [31:0] n44539;
wire     [31:0] n44540;
wire     [31:0] n44541;
wire     [31:0] n44542;
wire     [31:0] n44543;
wire     [31:0] n44544;
wire     [31:0] n44545;
wire     [31:0] n44546;
wire     [31:0] n44547;
wire     [31:0] n44548;
wire     [31:0] n44549;
wire     [31:0] n44550;
wire     [31:0] n44551;
wire     [31:0] n44552;
wire     [31:0] n44553;
wire     [31:0] n44554;
wire     [31:0] n44555;
wire     [31:0] n44556;
wire     [31:0] n44557;
wire     [31:0] n44558;
wire     [31:0] n44559;
wire     [31:0] n44560;
wire     [31:0] n44561;
wire     [31:0] n44562;
wire     [31:0] n44563;
wire     [31:0] n44564;
wire     [31:0] n44565;
wire     [31:0] n44566;
wire     [31:0] n44567;
wire     [31:0] n44568;
wire     [31:0] n44569;
wire     [31:0] n44570;
wire     [31:0] n44571;
wire     [31:0] n44572;
wire     [31:0] n44573;
wire     [31:0] n44574;
wire     [31:0] n44575;
wire     [31:0] n44576;
wire     [31:0] n44577;
wire     [31:0] n44578;
wire     [31:0] n44579;
wire     [31:0] n44580;
wire     [31:0] n44581;
wire     [31:0] n44582;
wire     [31:0] n44583;
wire     [31:0] n44584;
wire     [31:0] n44585;
wire     [31:0] n44586;
wire     [31:0] n44587;
wire     [31:0] n44588;
wire     [31:0] n44589;
wire     [31:0] n44590;
wire     [31:0] n44591;
wire     [31:0] n44592;
wire     [31:0] n44593;
wire     [31:0] n44594;
wire     [31:0] n44595;
wire     [31:0] n44596;
wire     [31:0] n44597;
wire     [31:0] n44598;
wire     [31:0] n44599;
wire     [31:0] n44600;
wire     [31:0] n44601;
wire     [31:0] n44602;
wire     [31:0] n44603;
wire     [31:0] n44604;
wire     [31:0] n44605;
wire     [31:0] n44606;
wire     [31:0] n44607;
wire     [31:0] n44608;
wire     [31:0] n44609;
wire     [31:0] n44610;
wire     [31:0] n44611;
wire     [31:0] n44612;
wire     [31:0] n44613;
wire     [31:0] n44614;
wire     [31:0] n44615;
wire     [31:0] n44616;
wire     [31:0] n44617;
wire     [31:0] n44618;
wire     [31:0] n44619;
wire     [31:0] n44620;
wire     [31:0] n44621;
wire     [31:0] n44622;
wire     [31:0] n44623;
wire     [31:0] n44624;
wire     [31:0] n44625;
wire     [31:0] n44626;
wire     [31:0] n44627;
wire     [31:0] n44628;
wire     [31:0] n44629;
wire     [31:0] n44630;
wire     [31:0] n44631;
wire     [31:0] n44632;
wire     [31:0] n44633;
wire     [31:0] n44634;
wire     [31:0] n44635;
wire     [31:0] n44636;
wire     [31:0] n44637;
wire     [31:0] n44638;
wire     [31:0] n44639;
wire     [31:0] n44640;
wire     [31:0] n44641;
wire     [31:0] n44642;
wire     [31:0] n44643;
wire     [31:0] n44644;
wire     [31:0] n44645;
wire     [31:0] n44646;
wire     [31:0] n44647;
wire     [31:0] n44648;
wire     [31:0] n44649;
wire     [31:0] n44650;
wire     [31:0] n44651;
wire     [31:0] n44652;
wire     [31:0] n44653;
wire     [31:0] n44654;
wire     [31:0] n44655;
wire     [31:0] n44656;
wire     [31:0] n44657;
wire     [31:0] n44658;
wire     [31:0] n44659;
wire     [31:0] n44660;
wire     [31:0] n44661;
wire     [31:0] n44662;
wire     [31:0] n44663;
wire     [31:0] n44664;
wire     [31:0] n44665;
wire     [31:0] n44666;
wire     [31:0] n44667;
wire     [31:0] n44668;
wire     [31:0] n44669;
wire     [31:0] n44670;
wire     [31:0] n44671;
wire     [31:0] n44672;
wire     [31:0] n44673;
wire     [31:0] n44674;
wire     [31:0] n44675;
wire     [31:0] n44676;
wire     [31:0] n44677;
wire     [31:0] n44678;
wire     [31:0] n44679;
wire     [31:0] n44680;
wire     [31:0] n44681;
wire     [31:0] n44682;
wire     [31:0] n44683;
wire     [31:0] n44684;
wire     [31:0] n44685;
wire     [31:0] n44686;
wire     [31:0] n44687;
wire     [31:0] n44688;
wire     [31:0] n44689;
wire     [31:0] n44690;
wire     [31:0] n44691;
wire     [31:0] n44692;
wire     [31:0] n44693;
wire     [31:0] n44694;
wire     [31:0] n44695;
wire     [31:0] n44696;
wire     [31:0] n44697;
wire     [31:0] n44698;
wire     [31:0] n44699;
wire     [31:0] n44700;
wire     [31:0] n44701;
wire     [31:0] n44702;
wire     [31:0] n44703;
wire     [31:0] n44704;
wire     [31:0] n44705;
wire     [31:0] n44706;
wire     [31:0] n44707;
wire     [31:0] n44708;
wire     [31:0] n44709;
wire     [31:0] n44710;
wire     [31:0] n44711;
wire     [31:0] n44712;
wire     [31:0] n44713;
wire     [31:0] n44714;
wire     [31:0] n44715;
wire     [31:0] n44716;
wire     [31:0] n44717;
wire     [31:0] n44718;
wire     [31:0] n44719;
wire     [31:0] n44720;
wire     [31:0] n44721;
wire     [31:0] n44722;
wire     [31:0] n44723;
wire     [31:0] n44724;
wire     [31:0] n44725;
wire     [31:0] n44726;
wire     [31:0] n44727;
wire     [31:0] n44728;
wire     [31:0] n44729;
wire     [31:0] n44730;
wire     [31:0] n44731;
wire     [31:0] n44732;
wire     [31:0] n44733;
wire     [31:0] n44734;
wire     [31:0] n44735;
wire     [31:0] n44736;
wire     [31:0] n44737;
wire     [31:0] n44738;
wire     [31:0] n44739;
wire     [31:0] n44740;
wire     [31:0] n44741;
wire     [31:0] n44742;
wire     [31:0] n44743;
wire     [31:0] n44744;
wire     [31:0] n44745;
wire     [31:0] n44746;
wire     [31:0] n44747;
wire     [31:0] n44748;
wire     [31:0] n44749;
wire     [31:0] n44750;
wire     [31:0] n44751;
wire     [31:0] n44752;
wire     [31:0] n44753;
wire     [31:0] n44754;
wire     [31:0] n44755;
wire     [31:0] n44756;
wire     [31:0] n44757;
wire     [31:0] n44758;
wire     [31:0] n44759;
wire     [31:0] n44760;
wire     [31:0] n44761;
wire     [31:0] n44762;
wire     [31:0] n44763;
wire     [31:0] n44764;
wire     [31:0] n44765;
wire     [31:0] n44766;
wire     [31:0] n44767;
wire     [31:0] n44768;
wire     [31:0] n44769;
wire     [31:0] n44770;
wire     [31:0] n44771;
wire     [31:0] n44772;
wire     [31:0] n44773;
wire     [31:0] n44774;
wire     [31:0] n44775;
wire     [31:0] n44776;
wire     [31:0] n44777;
wire     [31:0] n44778;
wire     [31:0] n44779;
wire     [31:0] n44780;
wire     [31:0] n44781;
wire     [31:0] n44782;
wire     [31:0] n44783;
wire     [31:0] n44784;
wire     [31:0] n44785;
wire     [31:0] n44786;
wire     [31:0] n44787;
wire     [31:0] n44788;
wire     [31:0] n44789;
wire     [31:0] n44790;
wire     [31:0] n44791;
wire     [31:0] n44792;
wire     [31:0] n44793;
wire     [31:0] n44794;
wire     [31:0] n44795;
wire     [31:0] n44796;
wire     [31:0] n44797;
wire     [31:0] n44798;
wire     [31:0] n44799;
wire     [31:0] n44800;
wire     [31:0] n44801;
wire     [31:0] n44802;
wire     [31:0] n44803;
wire     [31:0] n44804;
wire     [31:0] n44805;
wire     [31:0] n44806;
wire     [31:0] n44807;
wire     [31:0] n44808;
wire     [31:0] n44809;
wire     [31:0] n44810;
wire     [31:0] n44811;
wire     [31:0] n44812;
wire     [31:0] n44813;
wire     [31:0] n44814;
wire     [31:0] n44815;
wire     [31:0] n44816;
wire     [31:0] n44817;
wire     [31:0] n44818;
wire     [31:0] n44819;
wire     [31:0] n44820;
wire     [31:0] n44821;
wire     [31:0] n44822;
wire     [31:0] n44823;
wire     [31:0] n44824;
wire     [31:0] n44825;
wire     [31:0] n44826;
wire     [31:0] n44827;
wire     [31:0] n44828;
wire     [31:0] n44829;
wire     [31:0] n44830;
wire     [31:0] n44831;
wire     [31:0] n44832;
wire     [31:0] n44833;
wire     [31:0] n44834;
wire     [31:0] n44835;
wire     [31:0] n44836;
wire     [31:0] n44837;
wire     [31:0] n44838;
wire     [31:0] n44839;
wire     [31:0] n44840;
wire     [31:0] n44841;
wire     [31:0] n44842;
wire     [31:0] n44843;
wire     [31:0] n44844;
wire     [31:0] n44845;
wire     [31:0] n44846;
wire     [31:0] n44847;
wire     [31:0] n44848;
wire     [31:0] n44849;
wire     [31:0] n44850;
wire     [31:0] n44851;
wire     [31:0] n44852;
wire     [31:0] n44853;
wire     [31:0] n44854;
wire     [31:0] n44855;
wire     [31:0] n44856;
wire     [31:0] n44857;
wire     [31:0] n44858;
wire     [31:0] n44859;
wire     [31:0] n44860;
wire     [31:0] n44861;
wire     [31:0] n44862;
wire     [31:0] n44863;
wire     [31:0] n44864;
wire     [31:0] n44865;
wire     [31:0] n44866;
wire     [31:0] n44867;
wire     [31:0] n44868;
wire     [31:0] n44869;
wire     [31:0] n44870;
wire     [31:0] n44871;
wire     [31:0] n44872;
wire     [31:0] n44873;
wire     [31:0] n44874;
wire     [31:0] n44875;
wire     [31:0] n44876;
wire     [31:0] n44877;
wire     [31:0] n44878;
wire     [31:0] n44879;
wire     [31:0] n44880;
wire     [31:0] n44881;
wire     [31:0] n44882;
wire     [31:0] n44883;
wire     [31:0] n44884;
wire     [31:0] n44885;
wire     [31:0] n44886;
wire     [31:0] n44887;
wire     [31:0] n44888;
wire     [31:0] n44889;
wire     [31:0] n44890;
wire     [31:0] n44891;
wire     [31:0] n44892;
wire     [31:0] n44893;
wire     [31:0] n44894;
wire     [31:0] n44895;
wire     [31:0] n44896;
wire     [31:0] n44897;
wire     [31:0] n44898;
wire     [31:0] n44899;
wire     [31:0] n44900;
wire     [31:0] n44901;
wire     [31:0] n44902;
wire     [31:0] n44903;
wire     [31:0] n44904;
wire     [31:0] n44905;
wire     [31:0] n44906;
wire     [31:0] n44907;
wire     [31:0] n44908;
wire     [31:0] n44909;
wire     [31:0] n44910;
wire     [31:0] n44911;
wire     [31:0] n44912;
wire     [31:0] n44913;
wire     [31:0] n44914;
wire     [31:0] n44915;
wire     [31:0] n44916;
wire     [31:0] n44917;
wire     [31:0] n44918;
wire     [31:0] n44919;
wire     [31:0] n44920;
wire     [31:0] n44921;
wire     [31:0] n44922;
wire     [31:0] n44923;
wire     [31:0] n44924;
wire     [31:0] n44925;
wire     [31:0] n44926;
wire     [31:0] n44927;
wire     [31:0] n44928;
wire     [31:0] n44929;
wire     [31:0] n44930;
wire     [31:0] n44931;
wire     [31:0] n44932;
wire     [31:0] n44933;
wire     [31:0] n44934;
wire     [31:0] n44935;
wire     [31:0] n44936;
wire     [31:0] n44937;
wire     [31:0] n44938;
wire     [31:0] n44939;
wire     [31:0] n44940;
wire     [31:0] n44941;
wire     [31:0] n44942;
wire     [31:0] n44943;
wire     [31:0] n44944;
wire     [31:0] n44945;
wire     [31:0] n44946;
wire     [31:0] n44947;
wire     [31:0] n44948;
wire     [31:0] n44949;
wire     [31:0] n44950;
wire     [31:0] n44951;
wire     [31:0] n44952;
wire     [31:0] n44953;
wire     [31:0] n44954;
wire     [31:0] n44955;
wire     [31:0] n44956;
wire     [31:0] n44957;
wire     [31:0] n44958;
wire     [31:0] n44959;
wire     [31:0] n44960;
wire     [31:0] n44961;
wire     [31:0] n44962;
wire     [31:0] n44963;
wire     [31:0] n44964;
wire     [31:0] n44965;
wire     [31:0] n44966;
wire     [31:0] n44967;
wire     [31:0] n44968;
wire     [31:0] n44969;
wire     [31:0] n44970;
wire     [31:0] n44971;
wire     [31:0] n44972;
wire     [31:0] n44973;
wire     [31:0] n44974;
wire     [31:0] n44975;
wire     [31:0] n44976;
wire     [31:0] n44977;
wire     [31:0] n44978;
wire     [31:0] n44979;
wire     [31:0] n44980;
wire     [31:0] n44981;
wire     [31:0] n44982;
wire     [31:0] n44983;
wire     [31:0] n44984;
wire     [31:0] n44985;
wire     [31:0] n44986;
wire     [31:0] n44987;
wire     [31:0] n44988;
wire     [31:0] n44989;
wire     [31:0] n44990;
wire     [31:0] n44991;
wire     [31:0] n44992;
wire     [31:0] n44993;
wire     [31:0] n44994;
wire     [31:0] n44995;
wire     [31:0] n44996;
wire     [31:0] n44997;
wire     [31:0] n44998;
wire     [31:0] n44999;
wire     [31:0] n45000;
wire     [31:0] n45001;
wire     [31:0] n45002;
wire     [31:0] n45003;
wire     [31:0] n45004;
wire     [31:0] n45005;
wire     [31:0] n45006;
wire     [31:0] n45007;
wire     [31:0] n45008;
wire     [31:0] n45009;
wire     [31:0] n45010;
wire     [31:0] n45011;
wire     [31:0] n45012;
wire     [31:0] n45013;
wire     [31:0] n45014;
wire     [31:0] n45015;
wire     [31:0] n45016;
wire     [31:0] n45017;
wire     [31:0] n45018;
wire     [31:0] n45019;
wire     [31:0] n45020;
wire     [31:0] n45021;
wire     [31:0] n45022;
wire     [31:0] n45023;
wire     [31:0] n45024;
wire     [31:0] n45025;
wire     [31:0] n45026;
wire     [31:0] n45027;
wire     [31:0] n45028;
wire     [31:0] n45029;
wire     [31:0] n45030;
wire     [31:0] n45031;
wire     [31:0] n45032;
wire     [31:0] n45033;
wire     [31:0] n45034;
wire     [31:0] n45035;
wire     [31:0] n45036;
wire     [31:0] n45037;
wire     [31:0] n45038;
wire     [31:0] n45039;
wire     [31:0] n45040;
wire     [31:0] n45041;
wire     [31:0] n45042;
wire     [31:0] n45043;
wire     [31:0] n45044;
wire     [31:0] n45045;
wire     [31:0] n45046;
wire     [31:0] n45047;
wire     [31:0] n45048;
wire     [31:0] n45049;
wire     [31:0] n45050;
wire     [31:0] n45051;
wire     [31:0] n45052;
wire     [31:0] n45053;
wire     [31:0] n45054;
wire     [31:0] n45055;
wire     [31:0] n45056;
wire     [31:0] n45057;
wire     [31:0] n45058;
wire     [31:0] n45059;
wire     [31:0] n45060;
wire     [31:0] n45061;
wire     [31:0] n45062;
wire     [31:0] n45063;
wire     [31:0] n45064;
wire     [31:0] n45065;
wire     [31:0] n45066;
wire     [31:0] n45067;
wire     [31:0] n45068;
wire     [31:0] n45069;
wire     [31:0] n45070;
wire     [31:0] n45071;
wire     [31:0] n45072;
wire     [31:0] n45073;
wire     [31:0] n45074;
wire     [31:0] n45075;
wire     [31:0] n45076;
wire     [31:0] n45077;
wire     [31:0] n45078;
wire     [31:0] n45079;
wire     [31:0] n45080;
wire     [31:0] n45081;
wire     [31:0] n45082;
wire     [31:0] n45083;
wire     [31:0] n45084;
wire     [31:0] n45085;
wire     [31:0] n45086;
wire     [31:0] n45087;
wire     [31:0] n45088;
wire     [31:0] n45089;
wire     [31:0] n45090;
wire     [31:0] n45091;
wire     [31:0] n45092;
wire     [31:0] n45093;
wire     [31:0] n45094;
wire     [31:0] n45095;
wire     [31:0] n45096;
wire     [31:0] n45097;
wire     [31:0] n45098;
wire     [31:0] n45099;
wire     [31:0] n45100;
wire     [31:0] n45101;
wire     [31:0] n45102;
wire     [31:0] n45103;
wire     [31:0] n45104;
wire     [31:0] n45105;
wire     [31:0] n45106;
wire     [31:0] n45107;
wire     [31:0] n45108;
wire     [31:0] n45109;
wire     [31:0] n45110;
wire     [31:0] n45111;
wire     [31:0] n45112;
wire     [31:0] n45113;
wire     [31:0] n45114;
wire     [31:0] n45115;
wire     [31:0] n45116;
wire     [31:0] n45117;
wire     [31:0] n45118;
wire     [31:0] n45119;
wire     [31:0] n45120;
wire     [31:0] n45121;
wire     [31:0] n45122;
wire     [31:0] n45123;
wire     [31:0] n45124;
wire     [31:0] n45125;
wire     [31:0] n45126;
wire     [31:0] n45127;
wire     [31:0] n45128;
wire     [31:0] n45129;
wire     [31:0] n45130;
wire     [31:0] n45131;
wire     [31:0] n45132;
wire     [31:0] n45133;
wire     [31:0] n45134;
wire     [31:0] n45135;
wire     [31:0] n45136;
wire     [31:0] n45137;
wire     [31:0] n45138;
wire     [31:0] n45139;
wire     [31:0] n45140;
wire     [31:0] n45141;
wire     [31:0] n45142;
wire     [31:0] n45143;
wire     [31:0] n45144;
wire     [31:0] n45145;
wire     [31:0] n45146;
wire     [31:0] n45147;
wire     [31:0] n45148;
wire     [31:0] n45149;
wire     [31:0] n45150;
wire     [31:0] n45151;
wire     [31:0] n45152;
wire     [31:0] n45153;
wire     [31:0] n45154;
wire     [31:0] n45155;
wire     [31:0] n45156;
wire     [31:0] n45157;
wire     [31:0] n45158;
wire     [31:0] n45159;
wire     [31:0] n45160;
wire     [31:0] n45161;
wire     [31:0] n45162;
wire     [31:0] n45163;
wire     [31:0] n45164;
wire     [31:0] n45165;
wire     [31:0] n45166;
wire     [31:0] n45167;
wire     [31:0] n45168;
wire     [31:0] n45169;
wire     [31:0] n45170;
wire     [31:0] n45171;
wire     [31:0] n45172;
wire     [31:0] n45173;
wire     [31:0] n45174;
wire     [31:0] n45175;
wire     [31:0] n45176;
wire     [31:0] n45177;
wire     [31:0] n45178;
wire     [31:0] n45179;
wire     [31:0] n45180;
wire     [31:0] n45181;
wire     [31:0] n45182;
wire     [31:0] n45183;
wire     [31:0] n45184;
wire     [31:0] n45185;
wire     [31:0] n45186;
wire     [31:0] n45187;
wire     [31:0] n45188;
wire     [31:0] n45189;
wire     [31:0] n45190;
wire     [31:0] n45191;
wire     [31:0] n45192;
wire     [31:0] n45193;
wire     [31:0] n45194;
wire     [31:0] n45195;
wire     [31:0] n45196;
wire     [31:0] n45197;
wire     [31:0] n45198;
wire     [31:0] n45199;
wire     [31:0] n45200;
wire     [31:0] n45201;
wire     [31:0] n45202;
wire     [31:0] n45203;
wire     [31:0] n45204;
wire     [31:0] n45205;
wire     [31:0] n45206;
wire     [31:0] n45207;
wire     [31:0] n45208;
wire     [31:0] n45209;
wire     [31:0] n45210;
wire     [31:0] n45211;
wire     [31:0] n45212;
wire     [31:0] n45213;
wire     [31:0] n45214;
wire     [31:0] n45215;
wire     [31:0] n45216;
wire     [31:0] n45217;
wire     [31:0] n45218;
wire     [31:0] n45219;
wire     [31:0] n45220;
wire     [31:0] n45221;
wire     [31:0] n45222;
wire     [31:0] n45223;
wire     [31:0] n45224;
wire     [31:0] n45225;
wire     [31:0] n45226;
wire     [31:0] n45227;
wire     [31:0] n45228;
wire     [31:0] n45229;
wire     [31:0] n45230;
wire     [31:0] n45231;
wire     [31:0] n45232;
wire     [31:0] n45233;
wire     [31:0] n45234;
wire     [31:0] n45235;
wire     [31:0] n45236;
wire     [31:0] n45237;
wire     [31:0] n45238;
wire     [31:0] n45239;
wire     [31:0] n45240;
wire     [31:0] n45241;
wire     [31:0] n45242;
wire     [31:0] n45243;
wire     [31:0] n45244;
wire     [31:0] n45245;
wire     [31:0] n45246;
wire     [31:0] n45247;
wire     [31:0] n45248;
wire     [31:0] n45249;
wire     [31:0] n45250;
wire     [31:0] n45251;
wire     [31:0] n45252;
wire     [31:0] n45253;
wire     [31:0] n45254;
wire     [31:0] n45255;
wire     [31:0] n45256;
wire     [31:0] n45257;
wire     [31:0] n45258;
wire     [31:0] n45259;
wire     [31:0] n45260;
wire     [31:0] n45261;
wire     [31:0] n45262;
wire     [31:0] n45263;
wire     [31:0] n45264;
wire     [31:0] n45265;
wire     [31:0] n45266;
wire     [31:0] n45267;
wire     [31:0] n45268;
wire     [31:0] n45269;
wire     [31:0] n45270;
wire     [31:0] n45271;
wire     [31:0] n45272;
wire     [31:0] n45273;
wire     [31:0] n45274;
wire     [31:0] n45275;
wire     [31:0] n45276;
wire     [31:0] n45277;
wire     [31:0] n45278;
wire     [31:0] n45279;
wire     [31:0] n45280;
wire     [31:0] n45281;
wire     [31:0] n45282;
wire     [31:0] n45283;
wire     [31:0] n45284;
wire     [31:0] n45285;
wire     [31:0] n45286;
wire     [31:0] n45287;
wire     [31:0] n45288;
wire     [31:0] n45289;
wire     [31:0] n45290;
wire     [31:0] n45291;
wire     [31:0] n45292;
wire     [31:0] n45293;
wire     [31:0] n45294;
wire     [31:0] n45295;
wire     [31:0] n45296;
wire     [31:0] n45297;
wire     [31:0] n45298;
wire     [31:0] n45299;
wire     [31:0] n45300;
wire     [31:0] n45301;
wire     [31:0] n45302;
wire     [31:0] n45303;
wire     [31:0] n45304;
wire     [31:0] n45305;
wire     [31:0] n45306;
wire     [31:0] n45307;
wire     [31:0] n45308;
wire     [31:0] n45309;
wire     [31:0] n45310;
wire     [31:0] n45311;
wire     [31:0] n45312;
wire     [31:0] n45313;
wire     [31:0] n45314;
wire     [31:0] n45315;
wire     [31:0] n45316;
wire     [31:0] n45317;
wire     [31:0] n45318;
wire     [31:0] n45319;
wire     [31:0] n45320;
wire     [31:0] n45321;
wire     [31:0] n45322;
wire     [31:0] n45323;
wire     [31:0] n45324;
wire     [31:0] n45325;
wire     [31:0] n45326;
wire     [31:0] n45327;
wire     [31:0] n45328;
wire     [31:0] n45329;
wire     [31:0] n45330;
wire     [31:0] n45331;
wire     [31:0] n45332;
wire     [31:0] n45333;
wire     [31:0] n45334;
wire     [31:0] n45335;
wire     [31:0] n45336;
wire     [31:0] n45337;
wire     [31:0] n45338;
wire     [31:0] n45339;
wire     [31:0] n45340;
wire     [31:0] n45341;
wire     [31:0] n45342;
wire     [31:0] n45343;
wire     [31:0] n45344;
wire     [31:0] n45345;
wire     [31:0] n45346;
wire     [31:0] n45347;
wire     [31:0] n45348;
wire     [31:0] n45349;
wire     [31:0] n45350;
wire     [31:0] n45351;
wire     [31:0] n45352;
wire     [31:0] n45353;
wire     [31:0] n45354;
wire     [31:0] n45355;
wire     [31:0] n45356;
wire     [31:0] n45357;
wire     [31:0] n45358;
wire     [31:0] n45359;
wire     [31:0] n45360;
wire     [31:0] n45361;
wire     [31:0] n45362;
wire     [31:0] n45363;
wire     [31:0] n45364;
wire     [31:0] n45365;
wire     [31:0] n45366;
wire     [31:0] n45367;
wire     [31:0] n45368;
wire     [31:0] n45369;
wire     [31:0] n45370;
wire     [31:0] n45371;
wire     [31:0] n45372;
wire     [31:0] n45373;
wire     [31:0] n45374;
wire     [31:0] n45375;
wire     [31:0] n45376;
wire     [31:0] n45377;
wire     [31:0] n45378;
wire     [31:0] n45379;
wire     [31:0] n45380;
wire     [31:0] n45381;
wire     [31:0] n45382;
wire     [31:0] n45383;
wire     [31:0] n45384;
wire     [31:0] n45385;
wire     [31:0] n45386;
wire     [31:0] n45387;
wire     [31:0] n45388;
wire     [31:0] n45389;
wire     [31:0] n45390;
wire     [31:0] n45391;
wire     [31:0] n45392;
wire     [31:0] n45393;
wire     [31:0] n45394;
wire     [31:0] n45395;
wire     [31:0] n45396;
wire     [31:0] n45397;
wire     [31:0] n45398;
wire     [31:0] n45399;
wire     [31:0] n45400;
wire     [31:0] n45401;
wire     [31:0] n45402;
wire     [31:0] n45403;
wire     [31:0] n45404;
wire     [31:0] n45405;
wire     [31:0] n45406;
wire     [31:0] n45407;
wire     [31:0] n45408;
wire     [31:0] n45409;
wire     [31:0] n45410;
wire     [31:0] n45411;
wire     [31:0] n45412;
wire     [31:0] n45413;
wire     [31:0] n45414;
wire     [31:0] n45415;
wire     [31:0] n45416;
wire     [31:0] n45417;
wire     [31:0] n45418;
wire     [31:0] n45419;
wire     [31:0] n45420;
wire     [31:0] n45421;
wire     [31:0] n45422;
wire     [31:0] n45423;
wire     [31:0] n45424;
wire     [31:0] n45425;
wire     [31:0] n45426;
wire     [31:0] n45427;
wire     [31:0] n45428;
wire     [31:0] n45429;
wire     [31:0] n45430;
wire     [31:0] n45431;
wire     [31:0] n45432;
wire     [31:0] n45433;
wire     [31:0] n45434;
wire     [31:0] n45435;
wire     [31:0] n45436;
wire     [31:0] n45437;
wire     [31:0] n45438;
wire     [31:0] n45439;
wire     [31:0] n45440;
wire     [31:0] n45441;
wire     [31:0] n45442;
wire     [31:0] n45443;
wire     [31:0] n45444;
wire     [31:0] n45445;
wire     [31:0] n45446;
wire     [31:0] n45447;
wire     [31:0] n45448;
wire     [31:0] n45449;
wire     [31:0] n45450;
wire     [31:0] n45451;
wire     [31:0] n45452;
wire     [31:0] n45453;
wire     [31:0] n45454;
wire     [31:0] n45455;
wire     [31:0] n45456;
wire     [31:0] n45457;
wire     [31:0] n45458;
wire     [31:0] n45459;
wire     [31:0] n45460;
wire     [31:0] n45461;
wire     [31:0] n45462;
wire     [31:0] n45463;
wire     [31:0] n45464;
wire     [31:0] n45465;
wire     [31:0] n45466;
wire     [31:0] n45467;
wire     [31:0] n45468;
wire     [31:0] n45469;
wire     [31:0] n45470;
wire     [31:0] n45471;
wire     [31:0] n45472;
wire     [31:0] n45473;
wire     [31:0] n45474;
wire     [31:0] n45475;
wire     [31:0] n45476;
wire     [31:0] n45477;
wire     [31:0] n45478;
wire     [31:0] n45479;
wire     [31:0] n45480;
wire     [31:0] n45481;
wire     [31:0] n45482;
wire     [31:0] n45483;
wire     [31:0] n45484;
wire     [31:0] n45485;
wire     [31:0] n45486;
wire     [31:0] n45487;
wire     [31:0] n45488;
wire     [31:0] n45489;
wire     [31:0] n45490;
wire     [31:0] n45491;
wire     [31:0] n45492;
wire     [31:0] n45493;
wire     [31:0] n45494;
wire     [31:0] n45495;
wire     [31:0] n45496;
wire     [31:0] n45497;
wire     [31:0] n45498;
wire     [31:0] n45499;
wire     [31:0] n45500;
wire     [31:0] n45501;
wire     [31:0] n45502;
wire     [31:0] n45503;
wire     [31:0] n45504;
wire     [31:0] n45505;
wire     [31:0] n45506;
wire     [31:0] n45507;
wire     [31:0] n45508;
wire     [31:0] n45509;
wire     [31:0] n45510;
wire     [31:0] n45511;
wire     [31:0] n45512;
wire     [31:0] n45513;
wire     [31:0] n45514;
wire     [31:0] n45515;
wire     [31:0] n45516;
wire     [31:0] n45517;
wire     [31:0] n45518;
wire     [31:0] n45519;
wire     [31:0] n45520;
wire     [31:0] n45521;
wire     [31:0] n45522;
wire     [31:0] n45523;
wire     [31:0] n45524;
wire     [31:0] n45525;
wire     [31:0] n45526;
wire     [31:0] n45527;
wire     [31:0] n45528;
wire     [31:0] n45529;
wire     [31:0] n45530;
wire     [31:0] n45531;
wire     [31:0] n45532;
wire     [31:0] n45533;
wire     [31:0] n45534;
wire     [31:0] n45535;
wire     [31:0] n45536;
wire     [31:0] n45537;
wire     [31:0] n45538;
wire     [31:0] n45539;
wire     [31:0] n45540;
wire     [31:0] n45541;
wire     [31:0] n45542;
wire     [31:0] n45543;
wire     [31:0] n45544;
wire     [31:0] n45545;
wire     [31:0] n45546;
wire     [31:0] n45547;
wire     [31:0] n45548;
wire     [31:0] n45549;
wire     [31:0] n45550;
wire     [31:0] n45551;
wire     [31:0] n45552;
wire     [31:0] n45553;
wire     [31:0] n45554;
wire     [31:0] n45555;
wire     [31:0] n45556;
wire     [31:0] n45557;
wire     [31:0] n45558;
wire     [31:0] n45559;
wire     [31:0] n45560;
wire     [31:0] n45561;
wire     [31:0] n45562;
wire     [31:0] n45563;
wire     [31:0] n45564;
wire     [31:0] n45565;
wire     [31:0] n45566;
wire     [31:0] n45567;
wire     [31:0] n45568;
wire     [31:0] n45569;
wire     [31:0] n45570;
wire     [31:0] n45571;
wire     [31:0] n45572;
wire     [31:0] n45573;
wire     [31:0] n45574;
wire     [31:0] n45575;
wire     [31:0] n45576;
wire     [31:0] n45577;
wire     [31:0] n45578;
wire     [31:0] n45579;
wire     [31:0] n45580;
wire     [31:0] n45581;
wire     [31:0] n45582;
wire     [31:0] n45583;
wire     [31:0] n45584;
wire     [31:0] n45585;
wire     [31:0] n45586;
wire     [31:0] n45587;
wire     [31:0] n45588;
wire     [31:0] n45589;
wire     [31:0] n45590;
wire     [31:0] n45591;
wire     [31:0] n45592;
wire     [31:0] n45593;
wire     [31:0] n45594;
wire     [31:0] n45595;
wire     [31:0] n45596;
wire     [31:0] n45597;
wire     [31:0] n45598;
wire     [31:0] n45599;
wire     [31:0] n45600;
wire     [31:0] n45601;
wire     [31:0] n45602;
wire     [31:0] n45603;
wire     [31:0] n45604;
wire     [31:0] n45605;
wire     [31:0] n45606;
wire     [31:0] n45607;
wire     [31:0] n45608;
wire     [31:0] n45609;
wire     [31:0] n45610;
wire     [31:0] n45611;
wire     [31:0] n45612;
wire     [31:0] n45613;
wire     [31:0] n45614;
wire     [31:0] n45615;
wire     [31:0] n45616;
wire     [31:0] n45617;
wire     [31:0] n45618;
wire     [31:0] n45619;
wire     [31:0] n45620;
wire     [31:0] n45621;
wire     [31:0] n45622;
wire     [31:0] n45623;
wire     [31:0] n45624;
wire     [31:0] n45625;
wire     [31:0] n45626;
wire     [31:0] n45627;
wire     [31:0] n45628;
wire     [31:0] n45629;
wire     [31:0] n45630;
wire     [31:0] n45631;
wire     [31:0] n45632;
wire     [31:0] n45633;
wire     [31:0] n45634;
wire     [31:0] n45635;
wire     [31:0] n45636;
wire     [31:0] n45637;
wire     [31:0] n45638;
wire     [31:0] n45639;
wire     [31:0] n45640;
wire     [31:0] n45641;
wire     [31:0] n45642;
wire     [31:0] n45643;
wire     [31:0] n45644;
wire     [31:0] n45645;
wire     [31:0] n45646;
wire     [31:0] n45647;
wire     [31:0] n45648;
wire     [31:0] n45649;
wire     [31:0] n45650;
wire     [31:0] n45651;
wire     [31:0] n45652;
wire     [31:0] n45653;
wire     [31:0] n45654;
wire     [31:0] n45655;
wire     [31:0] n45656;
wire     [31:0] n45657;
wire     [31:0] n45658;
wire     [31:0] n45659;
wire     [31:0] n45660;
wire     [31:0] n45661;
wire     [31:0] n45662;
wire     [31:0] n45663;
wire     [31:0] n45664;
wire     [31:0] n45665;
wire     [31:0] n45666;
wire     [31:0] n45667;
wire     [31:0] n45668;
wire     [31:0] n45669;
wire     [31:0] n45670;
wire     [31:0] n45671;
wire     [31:0] n45672;
wire     [31:0] n45673;
wire     [31:0] n45674;
wire     [31:0] n45675;
wire     [31:0] n45676;
wire     [31:0] n45677;
wire     [31:0] n45678;
wire     [31:0] n45679;
wire     [31:0] n45680;
wire     [31:0] n45681;
wire     [31:0] n45682;
wire     [31:0] n45683;
wire     [31:0] n45684;
wire     [31:0] n45685;
wire     [31:0] n45686;
wire     [31:0] n45687;
wire     [31:0] n45688;
wire     [31:0] n45689;
wire     [31:0] n45690;
wire     [31:0] n45691;
wire     [31:0] n45692;
wire     [31:0] n45693;
wire     [31:0] n45694;
wire     [31:0] n45695;
wire     [31:0] n45696;
wire     [31:0] n45697;
wire     [31:0] n45698;
wire     [31:0] n45699;
wire     [31:0] n45700;
wire     [31:0] n45701;
wire     [31:0] n45702;
wire     [31:0] n45703;
wire     [31:0] n45704;
wire     [31:0] n45705;
wire     [31:0] n45706;
wire     [31:0] n45707;
wire     [31:0] n45708;
wire     [31:0] n45709;
wire     [31:0] n45710;
wire     [31:0] n45711;
wire     [31:0] n45712;
wire     [31:0] n45713;
wire     [31:0] n45714;
wire     [31:0] n45715;
wire     [31:0] n45716;
wire     [31:0] n45717;
wire     [31:0] n45718;
wire     [31:0] n45719;
wire     [31:0] n45720;
wire     [31:0] n45721;
wire     [31:0] n45722;
wire     [31:0] n45723;
wire     [31:0] n45724;
wire     [31:0] n45725;
wire     [31:0] n45726;
wire     [31:0] n45727;
wire     [31:0] n45728;
wire     [31:0] n45729;
wire     [31:0] n45730;
wire     [31:0] n45731;
wire     [31:0] n45732;
wire     [31:0] n45733;
wire     [31:0] n45734;
wire     [31:0] n45735;
wire     [31:0] n45736;
wire     [31:0] n45737;
wire     [31:0] n45738;
wire     [31:0] n45739;
wire     [31:0] n45740;
wire     [31:0] n45741;
wire     [31:0] n45742;
wire     [31:0] n45743;
wire     [31:0] n45744;
wire     [31:0] n45745;
wire     [31:0] n45746;
wire     [31:0] n45747;
wire     [31:0] n45748;
wire     [31:0] n45749;
wire     [31:0] n45750;
wire     [31:0] n45751;
wire     [31:0] n45752;
wire     [31:0] n45753;
wire     [31:0] n45754;
wire     [31:0] n45755;
wire     [31:0] n45756;
wire     [31:0] n45757;
wire     [31:0] n45758;
wire     [31:0] n45759;
wire     [31:0] n45760;
wire     [31:0] n45761;
wire     [31:0] n45762;
wire     [31:0] n45763;
wire     [31:0] n45764;
wire     [31:0] n45765;
wire     [31:0] n45766;
wire     [31:0] n45767;
wire     [31:0] n45768;
wire     [31:0] n45769;
wire     [31:0] n45770;
wire     [31:0] n45771;
wire     [31:0] n45772;
wire     [31:0] n45773;
wire     [31:0] n45774;
wire     [31:0] n45775;
wire     [31:0] n45776;
wire     [31:0] n45777;
wire     [31:0] n45778;
wire     [31:0] n45779;
wire     [31:0] n45780;
wire     [31:0] n45781;
wire     [31:0] n45782;
wire     [31:0] n45783;
wire     [31:0] n45784;
wire     [31:0] n45785;
wire     [31:0] n45786;
wire     [31:0] n45787;
wire     [31:0] n45788;
wire     [31:0] n45789;
wire     [31:0] n45790;
wire     [31:0] n45791;
wire     [31:0] n45792;
wire     [31:0] n45793;
wire     [31:0] n45794;
wire     [31:0] n45795;
wire     [31:0] n45796;
wire     [31:0] n45797;
wire     [31:0] n45798;
wire     [31:0] n45799;
wire     [31:0] n45800;
wire     [31:0] n45801;
wire     [31:0] n45802;
wire     [31:0] n45803;
wire     [31:0] n45804;
wire     [31:0] n45805;
wire     [31:0] n45806;
wire     [31:0] n45807;
wire     [31:0] n45808;
wire     [31:0] n45809;
wire     [31:0] n45810;
wire     [31:0] n45811;
wire     [31:0] n45812;
wire     [31:0] n45813;
wire     [31:0] n45814;
wire     [31:0] n45815;
wire     [31:0] n45816;
wire     [31:0] n45817;
wire     [31:0] n45818;
wire     [31:0] n45819;
wire     [31:0] n45820;
wire     [31:0] n45821;
wire     [31:0] n45822;
wire     [31:0] n45823;
wire     [31:0] n45824;
wire     [31:0] n45825;
wire     [31:0] n45826;
wire     [31:0] n45827;
wire     [31:0] n45828;
wire     [31:0] n45829;
wire     [31:0] n45830;
wire     [31:0] n45831;
wire     [31:0] n45832;
wire     [31:0] n45833;
wire     [31:0] n45834;
wire     [31:0] n45835;
wire     [31:0] n45836;
wire     [31:0] n45837;
wire     [31:0] n45838;
wire     [31:0] n45839;
wire     [31:0] n45840;
wire     [31:0] n45841;
wire     [31:0] n45842;
wire     [31:0] n45843;
wire     [31:0] n45844;
wire     [31:0] n45845;
wire     [31:0] n45846;
wire     [31:0] n45847;
wire     [31:0] n45848;
wire     [31:0] n45849;
wire     [31:0] n45850;
wire     [31:0] n45851;
wire     [31:0] n45852;
wire     [31:0] n45853;
wire     [31:0] n45854;
wire     [31:0] n45855;
wire     [31:0] n45856;
wire     [31:0] n45857;
wire     [31:0] n45858;
wire     [31:0] n45859;
wire     [31:0] n45860;
wire     [31:0] n45861;
wire     [31:0] n45862;
wire     [31:0] n45863;
wire     [31:0] n45864;
wire     [31:0] n45865;
wire     [31:0] n45866;
wire     [31:0] n45867;
wire     [31:0] n45868;
wire     [31:0] n45869;
wire     [31:0] n45870;
wire     [31:0] n45871;
wire     [31:0] n45872;
wire     [31:0] n45873;
wire     [31:0] n45874;
wire     [31:0] n45875;
wire     [31:0] n45876;
wire     [31:0] n45877;
wire     [31:0] n45878;
wire     [31:0] n45879;
wire     [31:0] n45880;
wire     [31:0] n45881;
wire     [31:0] n45882;
wire     [31:0] n45883;
wire     [31:0] n45884;
wire     [31:0] n45885;
wire     [31:0] n45886;
wire     [31:0] n45887;
wire     [31:0] n45888;
wire     [31:0] n45889;
wire     [31:0] n45890;
wire     [31:0] n45891;
wire     [31:0] n45892;
wire     [31:0] n45893;
wire     [31:0] n45894;
wire     [31:0] n45895;
wire     [31:0] n45896;
wire     [31:0] n45897;
wire     [31:0] n45898;
wire     [31:0] n45899;
wire     [31:0] n45900;
wire     [31:0] n45901;
wire     [31:0] n45902;
wire     [31:0] n45903;
wire     [31:0] n45904;
wire     [31:0] n45905;
wire     [31:0] n45906;
wire     [31:0] n45907;
wire     [31:0] n45908;
wire     [31:0] n45909;
wire     [31:0] n45910;
wire     [31:0] n45911;
wire     [31:0] n45912;
wire     [31:0] n45913;
wire     [31:0] n45914;
wire     [31:0] n45915;
wire     [31:0] n45916;
wire     [31:0] n45917;
wire     [31:0] n45918;
wire     [31:0] n45919;
wire     [31:0] n45920;
wire     [31:0] n45921;
wire     [31:0] n45922;
wire     [31:0] n45923;
wire     [31:0] n45924;
wire     [31:0] n45925;
wire     [31:0] n45926;
wire     [31:0] n45927;
wire     [31:0] n45928;
wire     [31:0] n45929;
wire     [31:0] n45930;
wire     [31:0] n45931;
wire     [31:0] n45932;
wire     [31:0] n45933;
wire     [31:0] n45934;
wire     [31:0] n45935;
wire     [31:0] n45936;
wire     [31:0] n45937;
wire     [31:0] n45938;
wire     [31:0] n45939;
wire     [31:0] n45940;
wire     [31:0] n45941;
wire     [31:0] n45942;
wire     [31:0] n45943;
wire     [31:0] n45944;
wire     [31:0] n45945;
wire     [31:0] n45946;
wire     [31:0] n45947;
wire     [31:0] n45948;
wire     [31:0] n45949;
wire     [31:0] n45950;
wire     [31:0] n45951;
wire     [31:0] n45952;
wire     [31:0] n45953;
wire     [31:0] n45954;
wire     [31:0] n45955;
wire     [31:0] n45956;
wire     [31:0] n45957;
wire     [31:0] n45958;
wire     [31:0] n45959;
wire     [31:0] n45960;
wire     [31:0] n45961;
wire     [31:0] n45962;
wire     [31:0] n45963;
wire     [31:0] n45964;
wire     [31:0] n45965;
wire     [31:0] n45966;
wire     [31:0] n45967;
wire     [31:0] n45968;
wire     [31:0] n45969;
wire     [31:0] n45970;
wire     [31:0] n45971;
wire     [31:0] n45972;
wire     [31:0] n45973;
wire     [31:0] n45974;
wire     [31:0] n45975;
wire     [31:0] n45976;
wire     [31:0] n45977;
wire     [31:0] n45978;
wire     [31:0] n45979;
wire     [31:0] n45980;
wire     [31:0] n45981;
wire     [31:0] n45982;
wire     [31:0] n45983;
wire     [31:0] n45984;
wire     [31:0] n45985;
wire     [31:0] n45986;
wire     [31:0] n45987;
wire     [31:0] n45988;
wire     [31:0] n45989;
wire     [31:0] n45990;
wire     [31:0] n45991;
wire     [31:0] n45992;
wire     [31:0] n45993;
wire     [31:0] n45994;
wire     [31:0] n45995;
wire     [31:0] n45996;
wire     [31:0] n45997;
wire     [31:0] n45998;
wire     [31:0] n45999;
wire     [31:0] n46000;
wire     [31:0] n46001;
wire     [31:0] n46002;
wire     [31:0] n46003;
wire     [31:0] n46004;
wire     [31:0] n46005;
wire     [31:0] n46006;
wire     [31:0] n46007;
wire     [31:0] n46008;
wire     [31:0] n46009;
wire     [31:0] n46010;
wire     [31:0] n46011;
wire     [31:0] n46012;
wire     [31:0] n46013;
wire     [31:0] n46014;
wire     [31:0] n46015;
wire     [31:0] n46016;
wire     [31:0] n46017;
wire     [31:0] n46018;
wire     [31:0] n46019;
wire     [31:0] n46020;
wire     [31:0] n46021;
wire     [31:0] n46022;
wire     [31:0] n46023;
wire     [31:0] n46024;
wire     [31:0] n46025;
wire     [31:0] n46026;
wire     [31:0] n46027;
wire     [31:0] n46028;
wire     [31:0] n46029;
wire     [31:0] n46030;
wire     [31:0] n46031;
wire     [31:0] n46032;
wire     [31:0] n46033;
wire     [31:0] n46034;
wire     [31:0] n46035;
wire     [31:0] n46036;
wire     [31:0] n46037;
wire     [31:0] n46038;
wire     [31:0] n46039;
wire     [31:0] n46040;
wire     [31:0] n46041;
wire     [31:0] n46042;
wire     [31:0] n46043;
wire     [31:0] n46044;
wire     [31:0] n46045;
wire     [31:0] n46046;
wire     [31:0] n46047;
wire     [31:0] n46048;
wire     [31:0] n46049;
wire     [31:0] n46050;
wire     [31:0] n46051;
wire     [31:0] n46052;
wire     [31:0] n46053;
wire     [31:0] n46054;
wire     [31:0] n46055;
wire     [31:0] n46056;
wire     [31:0] n46057;
wire     [31:0] n46058;
wire     [31:0] n46059;
wire     [31:0] n46060;
wire     [31:0] n46061;
wire     [31:0] n46062;
wire     [31:0] n46063;
wire     [31:0] n46064;
wire     [31:0] n46065;
wire     [31:0] n46066;
wire     [31:0] n46067;
wire     [31:0] n46068;
wire     [31:0] n46069;
wire     [31:0] n46070;
wire     [31:0] n46071;
wire     [31:0] n46072;
wire     [31:0] n46073;
wire     [31:0] n46074;
wire     [31:0] n46075;
wire     [31:0] n46076;
wire     [31:0] n46077;
wire     [31:0] n46078;
wire     [31:0] n46079;
wire     [31:0] n46080;
wire     [31:0] n46081;
wire     [31:0] n46082;
wire     [31:0] n46083;
wire     [31:0] n46084;
wire     [31:0] n46085;
wire     [31:0] n46086;
wire     [31:0] n46087;
wire     [31:0] n46088;
wire     [31:0] n46089;
wire     [31:0] n46090;
wire     [31:0] n46091;
wire     [31:0] n46092;
wire     [31:0] n46093;
wire     [31:0] n46094;
wire     [31:0] n46095;
wire     [31:0] n46096;
wire     [31:0] n46097;
wire     [31:0] n46098;
wire     [31:0] n46099;
wire     [31:0] n46100;
wire     [31:0] n46101;
wire     [31:0] n46102;
wire     [31:0] n46103;
wire     [31:0] n46104;
wire     [31:0] n46105;
wire     [31:0] n46106;
wire     [31:0] n46107;
wire     [31:0] n46108;
wire     [31:0] n46109;
wire     [31:0] n46110;
wire     [31:0] n46111;
wire     [31:0] n46112;
wire     [31:0] n46113;
wire     [31:0] n46114;
wire     [31:0] n46115;
wire     [31:0] n46116;
wire     [31:0] n46117;
wire     [31:0] n46118;
wire     [31:0] n46119;
wire     [31:0] n46120;
wire     [31:0] n46121;
wire     [31:0] n46122;
wire     [31:0] n46123;
wire     [31:0] n46124;
wire     [31:0] n46125;
wire     [31:0] n46126;
wire     [31:0] n46127;
wire     [31:0] n46128;
wire     [31:0] n46129;
wire     [31:0] n46130;
wire     [31:0] n46131;
wire     [31:0] n46132;
wire     [31:0] n46133;
wire     [31:0] n46134;
wire     [31:0] n46135;
wire     [31:0] n46136;
wire     [31:0] n46137;
wire     [31:0] n46138;
wire     [31:0] n46139;
wire     [31:0] n46140;
wire     [31:0] n46141;
wire     [31:0] n46142;
wire     [31:0] n46143;
wire     [31:0] n46144;
wire     [31:0] n46145;
wire     [31:0] n46146;
wire     [31:0] n46147;
wire     [31:0] n46148;
wire     [31:0] n46149;
wire     [31:0] n46150;
wire     [31:0] n46151;
wire     [31:0] n46152;
wire     [31:0] n46153;
wire     [31:0] n46154;
wire     [31:0] n46155;
wire     [31:0] n46156;
wire     [31:0] n46157;
wire     [31:0] n46158;
wire     [31:0] n46159;
wire     [31:0] n46160;
wire     [31:0] n46161;
wire     [31:0] n46162;
wire     [31:0] n46163;
wire     [31:0] n46164;
wire     [31:0] n46165;
wire     [31:0] n46166;
wire     [31:0] n46167;
wire     [31:0] n46168;
wire     [31:0] n46169;
wire     [31:0] n46170;
wire     [31:0] n46171;
wire     [31:0] n46172;
wire     [31:0] n46173;
wire     [31:0] n46174;
wire     [31:0] n46175;
wire     [31:0] n46176;
wire     [31:0] n46177;
wire     [31:0] n46178;
wire     [31:0] n46179;
wire     [31:0] n46180;
wire     [31:0] n46181;
wire     [31:0] n46182;
wire     [31:0] n46183;
wire     [31:0] n46184;
wire     [31:0] n46185;
wire     [31:0] n46186;
wire     [31:0] n46187;
wire     [31:0] n46188;
wire     [31:0] n46189;
wire     [31:0] n46190;
wire     [31:0] n46191;
wire     [31:0] n46192;
wire     [31:0] n46193;
wire     [31:0] n46194;
wire     [31:0] n46195;
wire     [31:0] n46196;
wire     [31:0] n46197;
wire     [31:0] n46198;
wire     [31:0] n46199;
wire     [31:0] n46200;
wire     [31:0] n46201;
wire     [31:0] n46202;
wire     [31:0] n46203;
wire     [31:0] n46204;
wire     [31:0] n46205;
wire     [31:0] n46206;
wire     [31:0] n46207;
wire     [31:0] n46208;
wire     [31:0] n46209;
wire     [31:0] n46210;
wire     [31:0] n46211;
wire     [31:0] n46212;
wire     [31:0] n46213;
wire     [31:0] n46214;
wire     [31:0] n46215;
wire     [31:0] n46216;
wire     [31:0] n46217;
wire     [31:0] n46218;
wire     [31:0] n46219;
wire     [31:0] n46220;
wire     [31:0] n46221;
wire     [31:0] n46222;
wire     [31:0] n46223;
wire     [31:0] n46224;
wire     [31:0] n46225;
wire     [31:0] n46226;
wire     [31:0] n46227;
wire     [31:0] n46228;
wire     [31:0] n46229;
wire     [31:0] n46230;
wire     [31:0] n46231;
wire     [31:0] n46232;
wire     [31:0] n46233;
wire     [31:0] n46234;
wire     [31:0] n46235;
wire     [31:0] n46236;
wire     [31:0] n46237;
wire     [31:0] n46238;
wire     [31:0] n46239;
wire     [31:0] n46240;
wire     [31:0] n46241;
wire     [31:0] n46242;
wire     [31:0] n46243;
wire     [31:0] n46244;
wire     [31:0] n46245;
wire     [31:0] n46246;
wire     [31:0] n46247;
wire     [31:0] n46248;
wire     [31:0] n46249;
wire     [31:0] n46250;
wire     [31:0] n46251;
wire     [31:0] n46252;
wire     [31:0] n46253;
wire     [31:0] n46254;
wire     [31:0] n46255;
wire     [31:0] n46256;
wire     [31:0] n46257;
wire     [31:0] n46258;
wire     [31:0] n46259;
wire     [31:0] n46260;
wire     [31:0] n46261;
wire     [31:0] n46262;
wire     [31:0] n46263;
wire     [31:0] n46264;
wire     [31:0] n46265;
wire     [31:0] n46266;
wire     [31:0] n46267;
wire     [31:0] n46268;
wire     [31:0] n46269;
wire     [31:0] n46270;
wire     [31:0] n46271;
wire     [31:0] n46272;
wire     [31:0] n46273;
wire     [31:0] n46274;
wire     [31:0] n46275;
wire     [31:0] n46276;
wire     [31:0] n46277;
wire     [31:0] n46278;
wire     [31:0] n46279;
wire     [31:0] n46280;
wire     [31:0] n46281;
wire     [31:0] n46282;
wire     [31:0] n46283;
wire     [31:0] n46284;
wire     [31:0] n46285;
wire     [31:0] n46286;
wire     [31:0] n46287;
wire     [31:0] n46288;
wire     [31:0] n46289;
wire     [31:0] n46290;
wire     [31:0] n46291;
wire     [31:0] n46292;
wire     [31:0] n46293;
wire     [31:0] n46294;
wire     [31:0] n46295;
wire     [31:0] n46296;
wire     [31:0] n46297;
wire     [31:0] n46298;
wire     [31:0] n46299;
wire     [31:0] n46300;
wire     [31:0] n46301;
wire     [31:0] n46302;
wire     [31:0] n46303;
wire     [31:0] n46304;
wire     [31:0] n46305;
wire     [31:0] n46306;
wire     [31:0] n46307;
wire     [31:0] n46308;
wire     [31:0] n46309;
wire     [31:0] n46310;
wire     [31:0] n46311;
wire     [31:0] n46312;
wire     [31:0] n46313;
wire     [31:0] n46314;
wire     [31:0] n46315;
wire     [31:0] n46316;
wire     [31:0] n46317;
wire     [31:0] n46318;
wire     [31:0] n46319;
wire     [31:0] n46320;
wire     [31:0] n46321;
wire     [31:0] n46322;
wire     [31:0] n46323;
wire     [31:0] n46324;
wire     [31:0] n46325;
wire     [31:0] n46326;
wire     [31:0] n46327;
wire     [31:0] n46328;
wire     [31:0] n46329;
wire     [31:0] n46330;
wire     [31:0] n46331;
wire     [31:0] n46332;
wire     [31:0] n46333;
wire     [31:0] n46334;
wire     [31:0] n46335;
wire     [31:0] n46336;
wire     [31:0] n46337;
wire     [31:0] n46338;
wire     [31:0] n46339;
wire     [31:0] n46340;
wire     [31:0] n46341;
wire     [31:0] n46342;
wire     [31:0] n46343;
wire     [31:0] n46344;
wire     [31:0] n46345;
wire     [31:0] n46346;
wire     [31:0] n46347;
wire     [31:0] n46348;
wire     [31:0] n46349;
wire     [31:0] n46350;
wire     [31:0] n46351;
wire     [31:0] n46352;
wire     [31:0] n46353;
wire     [31:0] n46354;
wire     [31:0] n46355;
wire     [31:0] n46356;
wire     [31:0] n46357;
wire     [31:0] n46358;
wire     [31:0] n46359;
wire     [31:0] n46360;
wire     [31:0] n46361;
wire     [31:0] n46362;
wire     [31:0] n46363;
wire     [31:0] n46364;
wire     [31:0] n46365;
wire     [31:0] n46366;
wire     [31:0] n46367;
wire     [31:0] n46368;
wire     [31:0] n46369;
wire     [31:0] n46370;
wire     [31:0] n46371;
wire     [31:0] n46372;
wire     [31:0] n46373;
wire     [31:0] n46374;
wire     [31:0] n46375;
wire     [31:0] n46376;
wire     [31:0] n46377;
wire     [31:0] n46378;
wire     [31:0] n46379;
wire     [31:0] n46380;
wire     [31:0] n46381;
wire     [31:0] n46382;
wire     [31:0] n46383;
wire     [31:0] n46384;
wire     [31:0] n46385;
wire     [31:0] n46386;
wire     [31:0] n46387;
wire     [31:0] n46388;
wire     [31:0] n46389;
wire     [31:0] n46390;
wire     [31:0] n46391;
wire     [31:0] n46392;
wire     [31:0] n46393;
wire     [31:0] n46394;
wire     [31:0] n46395;
wire     [31:0] n46396;
wire     [31:0] n46397;
wire     [31:0] n46398;
wire     [31:0] n46399;
wire     [31:0] n46400;
wire     [31:0] n46401;
wire     [31:0] n46402;
wire     [31:0] n46403;
wire     [31:0] n46404;
wire     [31:0] n46405;
wire     [31:0] n46406;
wire     [31:0] n46407;
wire     [31:0] n46408;
wire     [31:0] n46409;
wire     [31:0] n46410;
wire     [31:0] n46411;
wire     [31:0] n46412;
wire     [31:0] n46413;
wire     [31:0] n46414;
wire     [31:0] n46415;
wire     [31:0] n46416;
wire     [31:0] n46417;
wire     [31:0] n46418;
wire     [31:0] n46419;
wire     [31:0] n46420;
wire     [31:0] n46421;
wire     [31:0] n46422;
wire     [31:0] n46423;
wire     [31:0] n46424;
wire     [31:0] n46425;
wire     [31:0] n46426;
wire     [31:0] n46427;
wire     [31:0] n46428;
wire     [31:0] n46429;
wire     [31:0] n46430;
wire     [31:0] n46431;
wire     [31:0] n46432;
wire     [31:0] n46433;
wire     [31:0] n46434;
wire     [31:0] n46435;
wire     [31:0] n46436;
wire     [31:0] n46437;
wire     [31:0] n46438;
wire     [31:0] n46439;
wire     [31:0] n46440;
wire     [31:0] n46441;
wire     [31:0] n46442;
wire     [31:0] n46443;
wire     [31:0] n46444;
wire     [31:0] n46445;
wire     [31:0] n46446;
wire     [31:0] n46447;
wire     [31:0] n46448;
wire     [31:0] n46449;
wire     [31:0] n46450;
wire     [31:0] n46451;
wire     [31:0] n46452;
wire     [31:0] n46453;
wire     [31:0] n46454;
wire     [31:0] n46455;
wire     [31:0] n46456;
wire     [31:0] n46457;
wire     [31:0] n46458;
wire     [31:0] n46459;
wire     [31:0] n46460;
wire     [31:0] n46461;
wire     [31:0] n46462;
wire     [31:0] n46463;
wire     [31:0] n46464;
wire     [31:0] n46465;
wire     [31:0] n46466;
wire     [31:0] n46467;
wire     [31:0] n46468;
wire     [31:0] n46469;
wire     [31:0] n46470;
wire     [31:0] n46471;
wire     [31:0] n46472;
wire     [31:0] n46473;
wire     [31:0] n46474;
wire     [31:0] n46475;
wire     [31:0] n46476;
wire     [31:0] n46477;
wire     [31:0] n46478;
wire     [31:0] n46479;
wire     [31:0] n46480;
wire     [31:0] n46481;
wire     [31:0] n46482;
wire     [31:0] n46483;
wire     [31:0] n46484;
wire     [31:0] n46485;
wire     [31:0] n46486;
wire     [31:0] n46487;
wire     [31:0] n46488;
wire     [31:0] n46489;
wire     [31:0] n46490;
wire     [31:0] n46491;
wire     [31:0] n46492;
wire     [31:0] n46493;
wire     [31:0] n46494;
wire     [31:0] n46495;
wire     [31:0] n46496;
wire     [31:0] n46497;
wire     [31:0] n46498;
wire     [31:0] n46499;
wire     [31:0] n46500;
wire     [31:0] n46501;
wire     [31:0] n46502;
wire     [31:0] n46503;
wire     [31:0] n46504;
wire     [31:0] n46505;
wire     [31:0] n46506;
wire     [31:0] n46507;
wire     [31:0] n46508;
wire     [31:0] n46509;
wire     [31:0] n46510;
wire     [31:0] n46511;
wire     [31:0] n46512;
wire     [31:0] n46513;
wire     [31:0] n46514;
wire     [31:0] n46515;
wire     [31:0] n46516;
wire     [31:0] n46517;
wire     [31:0] n46518;
wire     [31:0] n46519;
wire     [31:0] n46520;
wire     [31:0] n46521;
wire     [31:0] n46522;
wire     [31:0] n46523;
wire     [31:0] n46524;
wire     [31:0] n46525;
wire     [31:0] n46526;
wire     [31:0] n46527;
wire     [31:0] n46528;
wire     [31:0] n46529;
wire     [31:0] n46530;
wire     [31:0] n46531;
wire     [31:0] n46532;
wire     [31:0] n46533;
wire     [31:0] n46534;
wire     [31:0] n46535;
wire     [31:0] n46536;
wire     [31:0] n46537;
wire     [31:0] n46538;
wire     [31:0] n46539;
wire     [31:0] n46540;
wire     [31:0] n46541;
wire     [31:0] n46542;
wire     [31:0] n46543;
wire     [31:0] n46544;
wire     [31:0] n46545;
wire     [31:0] n46546;
wire     [31:0] n46547;
wire     [31:0] n46548;
wire     [31:0] n46549;
wire     [31:0] n46550;
wire     [31:0] n46551;
wire     [31:0] n46552;
wire     [31:0] n46553;
wire     [31:0] n46554;
wire     [31:0] n46555;
wire     [31:0] n46556;
wire     [31:0] n46557;
wire     [31:0] n46558;
wire     [31:0] n46559;
wire     [31:0] n46560;
wire     [31:0] n46561;
wire     [31:0] n46562;
wire     [31:0] n46563;
wire     [31:0] n46564;
wire     [31:0] n46565;
wire     [31:0] n46566;
wire     [31:0] n46567;
wire     [31:0] n46568;
wire     [31:0] n46569;
wire     [31:0] n46570;
wire     [31:0] n46571;
wire     [31:0] n46572;
wire     [31:0] n46573;
wire     [31:0] n46574;
wire     [31:0] n46575;
wire     [31:0] n46576;
wire     [31:0] n46577;
wire     [31:0] n46578;
wire     [31:0] n46579;
wire     [31:0] n46580;
wire     [31:0] n46581;
wire     [31:0] n46582;
wire     [31:0] n46583;
wire     [31:0] n46584;
wire     [31:0] n46585;
wire     [31:0] n46586;
wire     [31:0] n46587;
wire     [31:0] n46588;
wire     [31:0] n46589;
wire     [31:0] n46590;
wire     [31:0] n46591;
wire     [31:0] n46592;
wire     [31:0] n46593;
wire     [31:0] n46594;
wire     [31:0] n46595;
wire     [31:0] n46596;
wire     [31:0] n46597;
wire     [31:0] n46598;
wire     [31:0] n46599;
wire     [31:0] n46600;
wire     [31:0] n46601;
wire     [31:0] n46602;
wire     [31:0] n46603;
wire     [31:0] n46604;
wire     [31:0] n46605;
wire     [31:0] n46606;
wire     [31:0] n46607;
wire     [31:0] n46608;
wire     [31:0] n46609;
wire     [31:0] n46610;
wire     [31:0] n46611;
wire     [31:0] n46612;
wire     [31:0] n46613;
wire     [31:0] n46614;
wire     [31:0] n46615;
wire     [31:0] n46616;
wire     [31:0] n46617;
wire     [31:0] n46618;
wire     [31:0] n46619;
wire     [31:0] n46620;
wire     [31:0] n46621;
wire     [31:0] n46622;
wire     [31:0] n46623;
wire     [31:0] n46624;
wire     [31:0] n46625;
wire     [31:0] n46626;
wire     [31:0] n46627;
wire     [31:0] n46628;
wire     [31:0] n46629;
wire     [31:0] n46630;
wire     [31:0] n46631;
wire     [31:0] n46632;
wire     [31:0] n46633;
wire     [31:0] n46634;
wire     [31:0] n46635;
wire     [31:0] n46636;
wire     [31:0] n46637;
wire     [31:0] n46638;
wire     [31:0] n46639;
wire     [31:0] n46640;
wire     [31:0] n46641;
wire     [31:0] n46642;
wire     [31:0] n46643;
wire     [31:0] n46644;
wire     [31:0] n46645;
wire     [31:0] n46646;
wire     [31:0] n46647;
wire     [31:0] n46648;
wire     [31:0] n46649;
wire     [31:0] n46650;
wire     [31:0] n46651;
wire     [31:0] n46652;
wire     [31:0] n46653;
wire     [31:0] n46654;
wire     [31:0] n46655;
wire     [31:0] n46656;
wire     [31:0] n46657;
wire     [31:0] n46658;
wire     [31:0] n46659;
wire     [31:0] n46660;
wire     [31:0] n46661;
wire     [31:0] n46662;
wire     [31:0] n46663;
wire     [31:0] n46664;
wire     [31:0] n46665;
wire     [31:0] n46666;
wire     [31:0] n46667;
wire     [31:0] n46668;
wire     [31:0] n46669;
wire     [31:0] n46670;
wire     [31:0] n46671;
wire     [31:0] n46672;
wire     [31:0] n46673;
wire     [31:0] n46674;
wire     [31:0] n46675;
wire     [31:0] n46676;
wire     [31:0] n46677;
wire     [31:0] n46678;
wire     [31:0] n46679;
wire     [31:0] n46680;
wire     [31:0] n46681;
wire     [31:0] n46682;
wire     [31:0] n46683;
wire     [31:0] n46684;
wire     [31:0] n46685;
wire     [31:0] n46686;
wire     [31:0] n46687;
wire     [31:0] n46688;
wire     [31:0] n46689;
wire     [31:0] n46690;
wire     [31:0] n46691;
wire     [31:0] n46692;
wire     [31:0] n46693;
wire     [31:0] n46694;
wire     [31:0] n46695;
wire     [31:0] n46696;
wire     [31:0] n46697;
wire     [31:0] n46698;
wire     [31:0] n46699;
wire     [31:0] n46700;
wire     [31:0] n46701;
wire     [31:0] n46702;
wire     [31:0] n46703;
wire     [31:0] n46704;
wire     [31:0] n46705;
wire     [31:0] n46706;
wire     [31:0] n46707;
wire     [31:0] n46708;
wire     [31:0] n46709;
wire     [31:0] n46710;
wire     [31:0] n46711;
wire     [31:0] n46712;
wire     [31:0] n46713;
wire     [31:0] n46714;
wire     [31:0] n46715;
wire     [31:0] n46716;
wire     [31:0] n46717;
wire     [31:0] n46718;
wire     [31:0] n46719;
wire     [31:0] n46720;
wire     [31:0] n46721;
wire     [31:0] n46722;
wire     [31:0] n46723;
wire     [31:0] n46724;
wire     [31:0] n46725;
wire     [31:0] n46726;
wire     [31:0] n46727;
wire     [31:0] n46728;
wire     [31:0] n46729;
wire     [31:0] n46730;
wire     [31:0] n46731;
wire     [31:0] n46732;
wire     [31:0] n46733;
wire     [31:0] n46734;
wire     [31:0] n46735;
wire     [31:0] n46736;
wire     [31:0] n46737;
wire     [31:0] n46738;
wire     [31:0] n46739;
wire     [31:0] n46740;
wire     [31:0] n46741;
wire     [31:0] n46742;
wire     [31:0] n46743;
wire     [31:0] n46744;
wire     [31:0] n46745;
wire     [31:0] n46746;
wire     [31:0] n46747;
wire     [31:0] n46748;
wire     [31:0] n46749;
wire     [31:0] n46750;
wire     [31:0] n46751;
wire     [31:0] n46752;
wire     [31:0] n46753;
wire     [31:0] n46754;
wire     [31:0] n46755;
wire     [31:0] n46756;
wire     [31:0] n46757;
wire     [31:0] n46758;
wire     [31:0] n46759;
wire     [31:0] n46760;
wire     [31:0] n46761;
wire     [31:0] n46762;
wire     [31:0] n46763;
wire     [31:0] n46764;
wire     [31:0] n46765;
wire     [31:0] n46766;
wire     [31:0] n46767;
wire     [31:0] n46768;
wire     [31:0] n46769;
wire     [31:0] n46770;
wire     [31:0] n46771;
wire     [31:0] n46772;
wire     [31:0] n46773;
wire     [31:0] n46774;
wire     [31:0] n46775;
wire     [31:0] n46776;
wire     [31:0] n46777;
wire     [31:0] n46778;
wire     [31:0] n46779;
wire     [31:0] n46780;
wire     [31:0] n46781;
wire     [31:0] n46782;
wire     [31:0] n46783;
wire     [31:0] n46784;
wire     [31:0] n46785;
wire     [31:0] n46786;
wire     [31:0] n46787;
wire     [31:0] n46788;
wire     [31:0] n46789;
wire     [31:0] n46790;
wire     [31:0] n46791;
wire     [31:0] n46792;
wire     [31:0] n46793;
wire     [31:0] n46794;
wire     [31:0] n46795;
wire     [31:0] n46796;
wire     [31:0] n46797;
wire     [31:0] n46798;
wire     [31:0] n46799;
wire     [31:0] n46800;
wire     [31:0] n46801;
wire     [31:0] n46802;
wire     [31:0] n46803;
wire     [31:0] n46804;
wire     [31:0] n46805;
wire     [31:0] n46806;
wire     [31:0] n46807;
wire     [31:0] n46808;
wire     [31:0] n46809;
wire     [31:0] n46810;
wire     [31:0] n46811;
wire     [31:0] n46812;
wire     [31:0] n46813;
wire     [31:0] n46814;
wire     [31:0] n46815;
wire     [31:0] n46816;
wire     [31:0] n46817;
wire     [31:0] n46818;
wire     [31:0] n46819;
wire     [31:0] n46820;
wire     [31:0] n46821;
wire     [31:0] n46822;
wire     [31:0] n46823;
wire     [31:0] n46824;
wire     [31:0] n46825;
wire     [31:0] n46826;
wire     [31:0] n46827;
wire     [31:0] n46828;
wire     [31:0] n46829;
wire     [31:0] n46830;
wire     [31:0] n46831;
wire     [31:0] n46832;
wire     [31:0] n46833;
wire     [31:0] n46834;
wire     [31:0] n46835;
wire     [31:0] n46836;
wire     [31:0] n46837;
wire     [31:0] n46838;
wire     [31:0] n46839;
wire     [31:0] n46840;
wire     [31:0] n46841;
wire     [31:0] n46842;
wire     [31:0] n46843;
wire     [31:0] n46844;
wire     [31:0] n46845;
wire     [31:0] n46846;
wire     [31:0] n46847;
wire     [31:0] n46848;
wire     [31:0] n46849;
wire     [31:0] n46850;
wire     [31:0] n46851;
wire     [31:0] n46852;
wire     [31:0] n46853;
wire     [31:0] n46854;
wire     [31:0] n46855;
wire     [31:0] n46856;
wire     [31:0] n46857;
wire     [31:0] n46858;
wire     [31:0] n46859;
wire     [31:0] n46860;
wire     [31:0] n46861;
wire     [31:0] n46862;
wire     [31:0] n46863;
wire     [31:0] n46864;
wire     [31:0] n46865;
wire     [31:0] n46866;
wire     [31:0] n46867;
wire     [31:0] n46868;
wire     [31:0] n46869;
wire     [31:0] n46870;
wire     [31:0] n46871;
wire     [31:0] n46872;
wire     [31:0] n46873;
wire     [31:0] n46874;
wire     [31:0] n46875;
wire     [31:0] n46876;
wire     [31:0] n46877;
wire     [31:0] n46878;
wire     [31:0] n46879;
wire     [31:0] n46880;
wire     [31:0] n46881;
wire     [31:0] n46882;
wire     [31:0] n46883;
wire     [31:0] n46884;
wire     [31:0] n46885;
wire     [31:0] n46886;
wire     [31:0] n46887;
wire     [31:0] n46888;
wire     [31:0] n46889;
wire     [31:0] n46890;
wire     [31:0] n46891;
wire     [31:0] n46892;
wire     [31:0] n46893;
wire     [31:0] n46894;
wire     [31:0] n46895;
wire     [31:0] n46896;
wire     [31:0] n46897;
wire     [31:0] n46898;
wire     [31:0] n46899;
wire     [31:0] n46900;
wire     [31:0] n46901;
wire     [31:0] n46902;
wire     [31:0] n46903;
wire     [31:0] n46904;
wire     [31:0] n46905;
wire     [31:0] n46906;
wire     [31:0] n46907;
wire     [31:0] n46908;
wire     [31:0] n46909;
wire     [31:0] n46910;
wire     [31:0] n46911;
wire     [31:0] n46912;
wire     [31:0] n46913;
wire     [31:0] n46914;
wire     [31:0] n46915;
wire     [31:0] n46916;
wire     [31:0] n46917;
wire     [31:0] n46918;
wire     [31:0] n46919;
wire     [31:0] n46920;
wire     [31:0] n46921;
wire     [31:0] n46922;
wire     [31:0] n46923;
wire     [31:0] n46924;
wire     [31:0] n46925;
wire     [31:0] n46926;
wire     [31:0] n46927;
wire     [31:0] n46928;
wire     [31:0] n46929;
wire     [31:0] n46930;
wire     [31:0] n46931;
wire     [31:0] n46932;
wire     [31:0] n46933;
wire     [31:0] n46934;
wire     [31:0] n46935;
wire     [31:0] n46936;
wire     [31:0] n46937;
wire     [31:0] n46938;
wire     [31:0] n46939;
wire     [31:0] n46940;
wire     [31:0] n46941;
wire     [31:0] n46942;
wire     [31:0] n46943;
wire     [31:0] n46944;
wire     [31:0] n46945;
wire     [31:0] n46946;
wire     [31:0] n46947;
wire     [31:0] n46948;
wire     [31:0] n46949;
wire     [31:0] n46950;
wire     [31:0] n46951;
wire     [31:0] n46952;
wire     [31:0] n46953;
wire     [31:0] n46954;
wire     [31:0] n46955;
wire     [31:0] n46956;
wire     [31:0] n46957;
wire     [31:0] n46958;
wire     [31:0] n46959;
wire     [31:0] n46960;
wire     [31:0] n46961;
wire     [31:0] n46962;
wire     [31:0] n46963;
wire     [31:0] n46964;
wire     [31:0] n46965;
wire     [31:0] n46966;
wire     [31:0] n46967;
wire     [31:0] n46968;
wire     [31:0] n46969;
wire     [31:0] n46970;
wire     [31:0] n46971;
wire     [31:0] n46972;
wire     [31:0] n46973;
wire     [31:0] n46974;
wire     [31:0] n46975;
wire     [31:0] n46976;
wire     [31:0] n46977;
wire     [31:0] n46978;
wire     [31:0] n46979;
wire     [31:0] n46980;
wire     [31:0] n46981;
wire     [31:0] n46982;
wire     [31:0] n46983;
wire     [31:0] n46984;
wire     [31:0] n46985;
wire     [31:0] n46986;
wire     [31:0] n46987;
wire     [31:0] n46988;
wire     [31:0] n46989;
wire     [31:0] n46990;
wire     [31:0] n46991;
wire     [31:0] n46992;
wire     [31:0] n46993;
wire     [31:0] n46994;
wire     [31:0] n46995;
wire     [31:0] n46996;
wire     [31:0] n46997;
wire     [31:0] n46998;
wire     [31:0] n46999;
wire     [31:0] n47000;
wire     [31:0] n47001;
wire     [31:0] n47002;
wire     [31:0] n47003;
wire     [31:0] n47004;
wire     [31:0] n47005;
wire     [31:0] n47006;
wire     [31:0] n47007;
wire     [31:0] n47008;
wire     [31:0] n47009;
wire     [31:0] n47010;
wire     [31:0] n47011;
wire     [31:0] n47012;
wire     [31:0] n47013;
wire     [31:0] n47014;
wire     [31:0] n47015;
wire     [31:0] n47016;
wire     [31:0] n47017;
wire     [31:0] n47018;
wire     [31:0] n47019;
wire     [31:0] n47020;
wire     [31:0] n47021;
wire     [31:0] n47022;
wire     [31:0] n47023;
wire     [31:0] n47024;
wire     [31:0] n47025;
wire     [31:0] n47026;
wire     [31:0] n47027;
wire     [31:0] n47028;
wire     [31:0] n47029;
wire     [31:0] n47030;
wire     [31:0] n47031;
wire     [31:0] n47032;
wire     [31:0] n47033;
wire     [31:0] n47034;
wire     [31:0] n47035;
wire     [31:0] n47036;
wire     [31:0] n47037;
wire     [31:0] n47038;
wire     [31:0] n47039;
wire     [31:0] n47040;
wire     [31:0] n47041;
wire     [31:0] n47042;
wire     [31:0] n47043;
wire     [31:0] n47044;
wire     [31:0] n47045;
wire     [31:0] n47046;
wire     [31:0] n47047;
wire     [31:0] n47048;
wire     [31:0] n47049;
wire     [31:0] n47050;
wire     [31:0] n47051;
wire     [31:0] n47052;
wire     [31:0] n47053;
wire     [31:0] n47054;
wire     [31:0] n47055;
wire     [31:0] n47056;
wire     [31:0] n47057;
wire     [31:0] n47058;
wire     [31:0] n47059;
wire     [31:0] n47060;
wire     [31:0] n47061;
wire     [31:0] n47062;
wire     [31:0] n47063;
wire     [31:0] n47064;
wire     [31:0] n47065;
wire     [31:0] n47066;
wire     [31:0] n47067;
wire     [31:0] n47068;
wire     [31:0] n47069;
wire     [31:0] n47070;
wire     [31:0] n47071;
wire     [31:0] n47072;
wire     [31:0] n47073;
wire     [31:0] n47074;
wire     [31:0] n47075;
wire     [31:0] n47076;
wire     [31:0] n47077;
wire     [31:0] n47078;
wire     [31:0] n47079;
wire     [31:0] n47080;
wire     [31:0] n47081;
wire     [31:0] n47082;
wire     [31:0] n47083;
wire     [31:0] n47084;
wire     [31:0] n47085;
wire     [31:0] n47086;
wire     [31:0] n47087;
wire     [31:0] n47088;
wire     [31:0] n47089;
wire     [31:0] n47090;
wire     [31:0] n47091;
wire     [31:0] n47092;
wire     [31:0] n47093;
wire     [31:0] n47094;
wire     [31:0] n47095;
wire     [31:0] n47096;
wire     [31:0] n47097;
wire     [31:0] n47098;
wire     [31:0] n47099;
wire     [31:0] n47100;
wire     [31:0] n47101;
wire     [31:0] n47102;
wire     [31:0] n47103;
wire     [31:0] n47104;
wire     [31:0] n47105;
wire     [31:0] n47106;
wire     [31:0] n47107;
wire     [31:0] n47108;
wire     [31:0] n47109;
wire     [31:0] n47110;
wire     [31:0] n47111;
wire     [31:0] n47112;
wire     [31:0] n47113;
wire     [31:0] n47114;
wire     [31:0] n47115;
wire     [31:0] n47116;
wire     [31:0] n47117;
wire     [31:0] n47118;
wire     [31:0] n47119;
wire     [31:0] n47120;
wire     [31:0] n47121;
wire     [31:0] n47122;
wire     [31:0] n47123;
wire     [31:0] n47124;
wire     [31:0] n47125;
wire     [31:0] n47126;
wire     [31:0] n47127;
wire     [31:0] n47128;
wire     [31:0] n47129;
wire     [31:0] n47130;
wire     [31:0] n47131;
wire     [31:0] n47132;
wire     [31:0] n47133;
wire     [31:0] n47134;
wire     [31:0] n47135;
wire     [31:0] n47136;
wire     [31:0] n47137;
wire     [31:0] n47138;
wire     [31:0] n47139;
wire     [31:0] n47140;
wire     [31:0] n47141;
wire     [31:0] n47142;
wire     [31:0] n47143;
wire     [31:0] n47144;
wire     [31:0] n47145;
wire     [31:0] n47146;
wire     [31:0] n47147;
wire     [31:0] n47148;
wire     [31:0] n47149;
wire     [31:0] n47150;
wire     [31:0] n47151;
wire     [31:0] n47152;
wire     [31:0] n47153;
wire     [31:0] n47154;
wire     [31:0] n47155;
wire     [31:0] n47156;
wire     [31:0] n47157;
wire     [31:0] n47158;
wire     [31:0] n47159;
wire     [31:0] n47160;
wire     [31:0] n47161;
wire     [31:0] n47162;
wire     [31:0] n47163;
wire     [31:0] n47164;
wire     [31:0] n47165;
wire     [31:0] n47166;
wire     [31:0] n47167;
wire     [31:0] n47168;
wire     [31:0] n47169;
wire     [31:0] n47170;
wire     [31:0] n47171;
wire     [31:0] n47172;
wire     [31:0] n47173;
wire     [31:0] n47174;
wire     [31:0] n47175;
wire     [31:0] n47176;
wire     [31:0] n47177;
wire     [31:0] n47178;
wire     [31:0] n47179;
wire     [31:0] n47180;
wire     [31:0] n47181;
wire     [31:0] n47182;
wire     [31:0] n47183;
wire     [31:0] n47184;
wire     [31:0] n47185;
wire     [31:0] n47186;
wire     [31:0] n47187;
wire     [31:0] n47188;
wire     [31:0] n47189;
wire     [31:0] n47190;
wire     [31:0] n47191;
wire     [31:0] n47192;
wire     [31:0] n47193;
wire     [31:0] n47194;
wire     [31:0] n47195;
wire     [31:0] n47196;
wire     [31:0] n47197;
wire     [31:0] n47198;
wire     [31:0] n47199;
wire     [31:0] n47200;
wire     [31:0] n47201;
wire     [31:0] n47202;
wire     [31:0] n47203;
wire     [31:0] n47204;
wire     [31:0] n47205;
wire     [31:0] n47206;
wire     [31:0] n47207;
wire     [31:0] n47208;
wire     [31:0] n47209;
wire     [31:0] n47210;
wire     [31:0] n47211;
wire     [31:0] n47212;
wire     [31:0] n47213;
wire     [31:0] n47214;
wire     [31:0] n47215;
wire     [31:0] n47216;
wire     [31:0] n47217;
wire     [31:0] n47218;
wire     [31:0] n47219;
wire     [31:0] n47220;
wire     [31:0] n47221;
wire     [31:0] n47222;
wire     [31:0] n47223;
wire     [31:0] n47224;
wire     [31:0] n47225;
wire     [31:0] n47226;
wire     [31:0] n47227;
wire     [31:0] n47228;
wire     [31:0] n47229;
wire     [31:0] n47230;
wire     [31:0] n47231;
wire     [31:0] n47232;
wire     [31:0] n47233;
wire     [31:0] n47234;
wire     [31:0] n47235;
wire     [31:0] n47236;
wire     [31:0] n47237;
wire     [31:0] n47238;
wire     [31:0] n47239;
wire     [31:0] n47240;
wire     [31:0] n47241;
wire     [31:0] n47242;
wire     [31:0] n47243;
wire     [31:0] n47244;
wire     [31:0] n47245;
wire     [31:0] n47246;
wire     [31:0] n47247;
wire     [31:0] n47248;
wire     [31:0] n47249;
wire     [31:0] n47250;
wire     [31:0] n47251;
wire     [31:0] n47252;
wire     [31:0] n47253;
wire     [31:0] n47254;
wire     [31:0] n47255;
wire     [31:0] n47256;
wire     [31:0] n47257;
wire     [31:0] n47258;
wire     [31:0] n47259;
wire     [31:0] n47260;
wire     [31:0] n47261;
wire     [31:0] n47262;
wire     [31:0] n47263;
wire     [31:0] n47264;
wire     [31:0] n47265;
wire     [31:0] n47266;
wire     [31:0] n47267;
wire     [31:0] n47268;
wire     [31:0] n47269;
wire     [31:0] n47270;
wire     [31:0] n47271;
wire     [31:0] n47272;
wire     [31:0] n47273;
wire     [31:0] n47274;
wire     [31:0] n47275;
wire     [31:0] n47276;
wire     [31:0] n47277;
wire     [31:0] n47278;
wire     [31:0] n47279;
wire     [31:0] n47280;
wire     [31:0] n47281;
wire     [31:0] n47282;
wire     [31:0] n47283;
wire     [31:0] n47284;
wire     [31:0] n47285;
wire     [31:0] n47286;
wire     [31:0] n47287;
wire     [31:0] n47288;
wire     [31:0] n47289;
wire     [31:0] n47290;
wire     [31:0] n47291;
wire     [31:0] n47292;
wire     [31:0] n47293;
wire     [31:0] n47294;
wire     [31:0] n47295;
wire     [31:0] n47296;
wire     [31:0] n47297;
wire     [31:0] n47298;
wire     [31:0] n47299;
wire     [31:0] n47300;
wire     [31:0] n47301;
wire     [31:0] n47302;
wire     [31:0] n47303;
wire     [31:0] n47304;
wire     [31:0] n47305;
wire     [31:0] n47306;
wire     [31:0] n47307;
wire     [31:0] n47308;
wire     [31:0] n47309;
wire     [31:0] n47310;
wire     [31:0] n47311;
wire     [31:0] n47312;
wire     [31:0] n47313;
wire     [31:0] n47314;
wire     [31:0] n47315;
wire     [31:0] n47316;
wire     [31:0] n47317;
wire     [31:0] n47318;
wire     [31:0] n47319;
wire     [31:0] n47320;
wire     [31:0] n47321;
wire     [31:0] n47322;
wire     [31:0] n47323;
wire     [31:0] n47324;
wire     [31:0] n47325;
wire     [31:0] n47326;
wire     [31:0] n47327;
wire     [31:0] n47328;
wire     [31:0] n47329;
wire     [31:0] n47330;
wire     [31:0] n47331;
wire     [31:0] n47332;
wire     [31:0] n47333;
wire     [31:0] n47334;
wire     [31:0] n47335;
wire     [31:0] n47336;
wire     [31:0] n47337;
wire     [31:0] n47338;
wire     [31:0] n47339;
wire     [31:0] n47340;
wire     [31:0] n47341;
wire     [31:0] n47342;
wire     [31:0] n47343;
wire     [31:0] n47344;
wire     [31:0] n47345;
wire     [31:0] n47346;
wire     [31:0] n47347;
wire     [31:0] n47348;
wire     [31:0] n47349;
wire     [31:0] n47350;
wire     [31:0] n47351;
wire     [31:0] n47352;
wire     [31:0] n47353;
wire     [31:0] n47354;
wire     [31:0] n47355;
wire     [31:0] n47356;
wire     [31:0] n47357;
wire     [31:0] n47358;
wire     [31:0] n47359;
wire     [31:0] n47360;
wire     [31:0] n47361;
wire     [31:0] n47362;
wire     [31:0] n47363;
wire     [31:0] n47364;
wire     [31:0] n47365;
wire     [31:0] n47366;
wire     [31:0] n47367;
wire     [31:0] n47368;
wire     [31:0] n47369;
wire     [31:0] n47370;
wire     [31:0] n47371;
wire     [31:0] n47372;
wire     [31:0] n47373;
wire     [31:0] n47374;
wire     [31:0] n47375;
wire     [31:0] n47376;
wire     [31:0] n47377;
wire     [31:0] n47378;
wire     [31:0] n47379;
wire     [31:0] n47380;
wire     [31:0] n47381;
wire     [31:0] n47382;
wire     [31:0] n47383;
wire     [31:0] n47384;
wire     [31:0] n47385;
wire     [31:0] n47386;
wire     [31:0] n47387;
wire     [31:0] n47388;
wire     [31:0] n47389;
wire     [31:0] n47390;
wire     [31:0] n47391;
wire     [31:0] n47392;
wire     [31:0] n47393;
wire     [31:0] n47394;
wire     [31:0] n47395;
wire     [31:0] n47396;
wire     [31:0] n47397;
wire     [31:0] n47398;
wire     [31:0] n47399;
wire     [31:0] n47400;
wire     [31:0] n47401;
wire     [31:0] n47402;
wire     [31:0] n47403;
wire     [31:0] n47404;
wire     [31:0] n47405;
wire     [31:0] n47406;
wire     [31:0] n47407;
wire     [31:0] n47408;
wire     [31:0] n47409;
wire     [31:0] n47410;
wire     [31:0] n47411;
wire     [31:0] n47412;
wire     [31:0] n47413;
wire     [31:0] n47414;
wire     [31:0] n47415;
wire     [31:0] n47416;
wire     [31:0] n47417;
wire     [31:0] n47418;
wire     [31:0] n47419;
wire     [31:0] n47420;
wire     [31:0] n47421;
wire     [31:0] n47422;
wire     [31:0] n47423;
wire     [31:0] n47424;
wire     [31:0] n47425;
wire     [31:0] n47426;
wire     [31:0] n47427;
wire     [31:0] n47428;
wire     [31:0] n47429;
wire     [31:0] n47430;
wire     [31:0] n47431;
wire     [31:0] n47432;
wire     [31:0] n47433;
wire     [31:0] n47434;
wire     [31:0] n47435;
wire     [31:0] n47436;
wire     [31:0] n47437;
wire     [31:0] n47438;
wire     [31:0] n47439;
wire     [31:0] n47440;
wire     [31:0] n47441;
wire     [31:0] n47442;
wire     [31:0] n47443;
wire     [31:0] n47444;
wire     [31:0] n47445;
wire     [31:0] n47446;
wire     [31:0] n47447;
wire     [31:0] n47448;
wire     [31:0] n47449;
wire     [31:0] n47450;
wire     [31:0] n47451;
wire     [31:0] n47452;
wire     [31:0] n47453;
wire     [31:0] n47454;
wire     [31:0] n47455;
wire     [31:0] n47456;
wire     [31:0] n47457;
wire     [31:0] n47458;
wire     [31:0] n47459;
wire     [31:0] n47460;
wire     [31:0] n47461;
wire     [31:0] n47462;
wire     [31:0] n47463;
wire     [31:0] n47464;
wire     [31:0] n47465;
wire     [31:0] n47466;
wire     [31:0] n47467;
wire     [31:0] n47468;
wire     [31:0] n47469;
wire     [31:0] n47470;
wire     [31:0] n47471;
wire     [31:0] n47472;
wire     [31:0] n47473;
wire     [31:0] n47474;
wire     [31:0] n47475;
wire     [31:0] n47476;
wire     [31:0] n47477;
wire     [31:0] n47478;
wire     [31:0] n47479;
wire     [31:0] n47480;
wire     [31:0] n47481;
wire     [31:0] n47482;
wire     [31:0] n47483;
wire     [31:0] n47484;
wire     [31:0] n47485;
wire     [31:0] n47486;
wire     [31:0] n47487;
wire     [31:0] n47488;
wire     [31:0] n47489;
wire     [31:0] n47490;
wire     [31:0] n47491;
wire     [31:0] n47492;
wire     [31:0] n47493;
wire     [31:0] n47494;
wire     [31:0] n47495;
wire     [31:0] n47496;
wire     [31:0] n47497;
wire     [31:0] n47498;
wire     [31:0] n47499;
wire     [31:0] n47500;
wire     [31:0] n47501;
wire     [31:0] n47502;
wire     [31:0] n47503;
wire     [31:0] n47504;
wire     [31:0] n47505;
wire     [31:0] n47506;
wire     [31:0] n47507;
wire     [31:0] n47508;
wire     [31:0] n47509;
wire     [31:0] n47510;
wire     [31:0] n47511;
wire     [31:0] n47512;
wire     [31:0] n47513;
wire     [31:0] n47514;
wire     [31:0] n47515;
wire     [31:0] n47516;
wire     [31:0] n47517;
wire     [31:0] n47518;
wire     [31:0] n47519;
wire     [31:0] n47520;
wire     [31:0] n47521;
wire     [31:0] n47522;
wire     [31:0] n47523;
wire     [31:0] n47524;
wire     [31:0] n47525;
wire     [31:0] n47526;
wire     [31:0] n47527;
wire     [31:0] n47528;
wire     [31:0] n47529;
wire     [31:0] n47530;
wire     [31:0] n47531;
wire     [31:0] n47532;
wire     [31:0] n47533;
wire     [31:0] n47534;
wire     [31:0] n47535;
wire     [31:0] n47536;
wire     [31:0] n47537;
wire     [31:0] n47538;
wire     [31:0] n47539;
wire     [31:0] n47540;
wire     [31:0] n47541;
wire     [31:0] n47542;
wire     [31:0] n47543;
wire     [31:0] n47544;
wire     [31:0] n47545;
wire     [31:0] n47546;
wire     [31:0] n47547;
wire     [31:0] n47548;
wire     [31:0] n47549;
wire     [31:0] n47550;
wire     [31:0] n47551;
wire     [31:0] n47552;
wire     [31:0] n47553;
wire     [31:0] n47554;
wire     [31:0] n47555;
wire     [31:0] n47556;
wire     [31:0] n47557;
wire     [31:0] n47558;
wire     [31:0] n47559;
wire     [31:0] n47560;
wire     [31:0] n47561;
wire     [31:0] n47562;
wire     [31:0] n47563;
wire     [31:0] n47564;
wire     [31:0] n47565;
wire     [31:0] n47566;
wire     [31:0] n47567;
wire     [31:0] n47568;
wire     [31:0] n47569;
wire     [31:0] n47570;
wire     [31:0] n47571;
wire     [31:0] n47572;
wire     [31:0] n47573;
wire     [31:0] n47574;
wire     [31:0] n47575;
wire     [31:0] n47576;
wire     [31:0] n47577;
wire     [31:0] n47578;
wire     [31:0] n47579;
wire     [31:0] n47580;
wire     [31:0] n47581;
wire     [31:0] n47582;
wire     [31:0] n47583;
wire     [31:0] n47584;
wire     [31:0] n47585;
wire     [31:0] n47586;
wire     [31:0] n47587;
wire     [31:0] n47588;
wire     [31:0] n47589;
wire     [31:0] n47590;
wire     [31:0] n47591;
wire     [31:0] n47592;
wire     [31:0] n47593;
wire     [31:0] n47594;
wire     [31:0] n47595;
wire     [31:0] n47596;
wire     [31:0] n47597;
wire     [31:0] n47598;
wire     [31:0] n47599;
wire     [31:0] n47600;
wire     [31:0] n47601;
wire     [31:0] n47602;
wire     [31:0] n47603;
wire     [31:0] n47604;
wire     [31:0] n47605;
wire     [31:0] n47606;
wire     [31:0] n47607;
wire     [31:0] n47608;
wire     [31:0] n47609;
wire     [31:0] n47610;
wire     [31:0] n47611;
wire     [31:0] n47612;
wire     [31:0] n47613;
wire     [31:0] n47614;
wire     [31:0] n47615;
wire     [31:0] n47616;
wire     [31:0] n47617;
wire     [31:0] n47618;
wire     [31:0] n47619;
wire     [31:0] n47620;
wire     [31:0] n47621;
wire     [31:0] n47622;
wire     [31:0] n47623;
wire     [31:0] n47624;
wire     [31:0] n47625;
wire     [31:0] n47626;
wire     [31:0] n47627;
wire     [31:0] n47628;
wire     [31:0] n47629;
wire     [31:0] n47630;
wire     [31:0] n47631;
wire     [31:0] n47632;
wire     [31:0] n47633;
wire     [31:0] n47634;
wire     [31:0] n47635;
wire     [31:0] n47636;
wire     [31:0] n47637;
wire     [31:0] n47638;
wire     [31:0] n47639;
wire     [31:0] n47640;
wire     [31:0] n47641;
wire     [31:0] n47642;
wire     [31:0] n47643;
wire     [31:0] n47644;
wire     [31:0] n47645;
wire     [31:0] n47646;
wire     [31:0] n47647;
wire     [31:0] n47648;
wire     [31:0] n47649;
wire     [31:0] n47650;
wire     [31:0] n47651;
wire     [31:0] n47652;
wire     [31:0] n47653;
wire     [31:0] n47654;
wire     [31:0] n47655;
wire     [31:0] n47656;
wire     [31:0] n47657;
wire     [31:0] n47658;
wire     [31:0] n47659;
wire     [31:0] n47660;
wire     [31:0] n47661;
wire     [31:0] n47662;
wire     [31:0] n47663;
wire     [31:0] n47664;
wire     [31:0] n47665;
wire     [31:0] n47666;
wire     [31:0] n47667;
wire     [31:0] n47668;
wire     [31:0] n47669;
wire     [31:0] n47670;
wire     [31:0] n47671;
wire     [31:0] n47672;
wire     [31:0] n47673;
wire     [31:0] n47674;
wire     [31:0] n47675;
wire     [31:0] n47676;
wire     [31:0] n47677;
wire     [31:0] n47678;
wire     [31:0] n47679;
wire     [31:0] n47680;
wire     [31:0] n47681;
wire     [31:0] n47682;
wire     [31:0] n47683;
wire     [31:0] n47684;
wire     [31:0] n47685;
wire     [31:0] n47686;
wire     [31:0] n47687;
wire     [31:0] n47688;
wire     [31:0] n47689;
wire     [31:0] n47690;
wire     [31:0] n47691;
wire     [31:0] n47692;
wire     [31:0] n47693;
wire     [31:0] n47694;
wire     [31:0] n47695;
wire     [31:0] n47696;
wire     [31:0] n47697;
wire     [31:0] n47698;
wire     [31:0] n47699;
wire     [31:0] n47700;
wire     [31:0] n47701;
wire     [31:0] n47702;
wire     [31:0] n47703;
wire     [31:0] n47704;
wire     [31:0] n47705;
wire     [31:0] n47706;
wire     [31:0] n47707;
wire     [31:0] n47708;
wire     [31:0] n47709;
wire     [31:0] n47710;
wire     [31:0] n47711;
wire     [31:0] n47712;
wire     [31:0] n47713;
wire     [31:0] n47714;
wire     [31:0] n47715;
wire     [31:0] n47716;
wire     [31:0] n47717;
wire     [31:0] n47718;
wire     [31:0] n47719;
wire     [31:0] n47720;
wire     [31:0] n47721;
wire     [31:0] n47722;
wire     [31:0] n47723;
wire     [31:0] n47724;
wire     [31:0] n47725;
wire     [31:0] n47726;
wire     [31:0] n47727;
wire     [31:0] n47728;
wire     [31:0] n47729;
wire     [31:0] n47730;
wire     [31:0] n47731;
wire     [31:0] n47732;
wire     [31:0] n47733;
wire     [31:0] n47734;
wire     [31:0] n47735;
wire     [31:0] n47736;
wire     [31:0] n47737;
wire     [31:0] n47738;
wire     [31:0] n47739;
wire     [31:0] n47740;
wire     [31:0] n47741;
wire     [31:0] n47742;
wire     [31:0] n47743;
wire     [31:0] n47744;
wire     [31:0] n47745;
wire     [31:0] n47746;
wire     [31:0] n47747;
wire     [31:0] n47748;
wire     [31:0] n47749;
wire     [31:0] n47750;
wire     [31:0] n47751;
wire     [31:0] n47752;
wire     [31:0] n47753;
wire     [31:0] n47754;
wire     [31:0] n47755;
wire     [31:0] n47756;
wire     [31:0] n47757;
wire     [31:0] n47758;
wire     [31:0] n47759;
wire     [31:0] n47760;
wire     [31:0] n47761;
wire     [31:0] n47762;
wire     [31:0] n47763;
wire     [31:0] n47764;
wire     [31:0] n47765;
wire     [31:0] n47766;
wire     [31:0] n47767;
wire     [31:0] n47768;
wire     [31:0] n47769;
wire     [31:0] n47770;
wire     [31:0] n47771;
wire     [31:0] n47772;
wire     [31:0] n47773;
wire     [31:0] n47774;
wire     [31:0] n47775;
wire     [31:0] n47776;
wire     [31:0] n47777;
wire     [31:0] n47778;
wire     [31:0] n47779;
wire     [31:0] n47780;
wire     [31:0] n47781;
wire     [31:0] n47782;
wire     [31:0] n47783;
wire     [31:0] n47784;
wire     [31:0] n47785;
wire     [31:0] n47786;
wire     [31:0] n47787;
wire     [31:0] n47788;
wire     [31:0] n47789;
wire     [31:0] n47790;
wire     [31:0] n47791;
wire     [31:0] n47792;
wire     [31:0] n47793;
wire     [31:0] n47794;
wire     [31:0] n47795;
wire     [31:0] n47796;
wire     [31:0] n47797;
wire     [31:0] n47798;
wire     [31:0] n47799;
wire     [31:0] n47800;
wire     [31:0] n47801;
wire     [31:0] n47802;
wire     [31:0] n47803;
wire     [31:0] n47804;
wire     [31:0] n47805;
wire     [31:0] n47806;
wire     [31:0] n47807;
wire     [31:0] n47808;
wire     [31:0] n47809;
wire     [31:0] n47810;
wire     [31:0] n47811;
wire     [31:0] n47812;
wire     [31:0] n47813;
wire     [31:0] n47814;
wire     [31:0] n47815;
wire     [31:0] n47816;
wire     [31:0] n47817;
wire     [31:0] n47818;
wire     [31:0] n47819;
wire     [31:0] n47820;
wire     [31:0] n47821;
wire     [31:0] n47822;
wire     [31:0] n47823;
wire     [31:0] n47824;
wire     [31:0] n47825;
wire     [31:0] n47826;
wire     [31:0] n47827;
wire     [31:0] n47828;
wire     [31:0] n47829;
wire     [31:0] n47830;
wire     [31:0] n47831;
wire     [31:0] n47832;
wire     [31:0] n47833;
wire     [31:0] n47834;
wire     [31:0] n47835;
wire     [31:0] n47836;
wire     [31:0] n47837;
wire     [31:0] n47838;
wire     [31:0] n47839;
wire     [31:0] n47840;
wire     [31:0] n47841;
wire     [31:0] n47842;
wire     [31:0] n47843;
wire     [31:0] n47844;
wire     [31:0] n47845;
wire     [31:0] n47846;
wire     [31:0] n47847;
wire     [31:0] n47848;
wire     [31:0] n47849;
wire     [31:0] n47850;
wire     [31:0] n47851;
wire     [31:0] n47852;
wire     [31:0] n47853;
wire     [31:0] n47854;
wire     [31:0] n47855;
wire     [31:0] n47856;
wire     [31:0] n47857;
wire     [31:0] n47858;
wire     [31:0] n47859;
wire     [31:0] n47860;
wire     [31:0] n47861;
wire     [31:0] n47862;
wire     [31:0] n47863;
wire     [31:0] n47864;
wire     [31:0] n47865;
wire     [31:0] n47866;
wire     [31:0] n47867;
wire     [31:0] n47868;
wire     [31:0] n47869;
wire     [31:0] n47870;
wire     [31:0] n47871;
wire     [31:0] n47872;
wire     [31:0] n47873;
wire     [31:0] n47874;
wire     [31:0] n47875;
wire     [31:0] n47876;
wire     [31:0] n47877;
wire     [31:0] n47878;
wire     [31:0] n47879;
wire     [31:0] n47880;
wire     [31:0] n47881;
wire     [31:0] n47882;
wire     [31:0] n47883;
wire     [31:0] n47884;
wire     [31:0] n47885;
wire     [31:0] n47886;
wire     [31:0] n47887;
wire     [31:0] n47888;
wire     [31:0] n47889;
wire     [31:0] n47890;
wire     [31:0] n47891;
wire     [31:0] n47892;
wire     [31:0] n47893;
wire     [31:0] n47894;
wire     [31:0] n47895;
wire     [31:0] n47896;
wire     [31:0] n47897;
wire     [31:0] n47898;
wire     [31:0] n47899;
wire     [31:0] n47900;
wire     [31:0] n47901;
wire     [31:0] n47902;
wire     [31:0] n47903;
wire     [31:0] n47904;
wire     [31:0] n47905;
wire     [31:0] n47906;
wire     [31:0] n47907;
wire     [31:0] n47908;
wire     [31:0] n47909;
wire     [31:0] n47910;
wire     [31:0] n47911;
wire     [31:0] n47912;
wire     [31:0] n47913;
wire     [31:0] n47914;
wire     [31:0] n47915;
wire     [31:0] n47916;
wire     [31:0] n47917;
wire     [31:0] n47918;
wire     [31:0] n47919;
wire     [31:0] n47920;
wire     [31:0] n47921;
wire     [31:0] n47922;
wire     [31:0] n47923;
wire     [31:0] n47924;
wire     [31:0] n47925;
wire     [31:0] n47926;
wire     [31:0] n47927;
wire     [31:0] n47928;
wire     [31:0] n47929;
wire     [31:0] n47930;
wire     [31:0] n47931;
wire     [31:0] n47932;
wire     [31:0] n47933;
wire     [31:0] n47934;
wire     [31:0] n47935;
wire     [31:0] n47936;
wire     [31:0] n47937;
wire     [31:0] n47938;
wire     [31:0] n47939;
wire     [31:0] n47940;
wire     [31:0] n47941;
wire     [31:0] n47942;
wire     [31:0] n47943;
wire     [31:0] n47944;
wire     [31:0] n47945;
wire     [31:0] n47946;
wire     [31:0] n47947;
wire     [31:0] n47948;
wire     [31:0] n47949;
wire     [31:0] n47950;
wire     [31:0] n47951;
wire     [31:0] n47952;
wire     [31:0] n47953;
wire     [31:0] n47954;
wire     [31:0] n47955;
wire     [31:0] n47956;
wire     [31:0] n47957;
wire     [31:0] n47958;
wire     [31:0] n47959;
wire     [31:0] n47960;
wire     [31:0] n47961;
wire     [31:0] n47962;
wire     [31:0] n47963;
wire     [31:0] n47964;
wire     [31:0] n47965;
wire     [31:0] n47966;
wire     [31:0] n47967;
wire     [31:0] n47968;
wire     [31:0] n47969;
wire     [31:0] n47970;
wire     [31:0] n47971;
wire     [31:0] n47972;
wire     [31:0] n47973;
wire     [31:0] n47974;
wire     [31:0] n47975;
wire     [31:0] n47976;
wire     [31:0] n47977;
wire     [31:0] n47978;
wire     [31:0] n47979;
wire     [31:0] n47980;
wire     [31:0] n47981;
wire     [31:0] n47982;
wire     [31:0] n47983;
wire     [31:0] n47984;
wire     [31:0] n47985;
wire     [31:0] n47986;
wire     [31:0] n47987;
wire     [31:0] n47988;
wire     [31:0] n47989;
wire     [31:0] n47990;
wire     [31:0] n47991;
wire     [31:0] n47992;
wire     [31:0] n47993;
wire     [31:0] n47994;
wire     [31:0] n47995;
wire     [31:0] n47996;
wire     [31:0] n47997;
wire     [31:0] n47998;
wire     [31:0] n47999;
wire     [31:0] n48000;
wire     [31:0] n48001;
wire     [31:0] n48002;
wire     [31:0] n48003;
wire     [31:0] n48004;
wire     [31:0] n48005;
wire     [31:0] n48006;
wire     [31:0] n48007;
wire     [31:0] n48008;
wire     [31:0] n48009;
wire     [31:0] n48010;
wire     [31:0] n48011;
wire     [31:0] n48012;
wire     [31:0] n48013;
wire     [31:0] n48014;
wire     [31:0] n48015;
wire     [31:0] n48016;
wire     [31:0] n48017;
wire     [31:0] n48018;
wire     [31:0] n48019;
wire     [31:0] n48020;
wire     [31:0] n48021;
wire     [31:0] n48022;
wire     [31:0] n48023;
wire     [31:0] n48024;
wire     [31:0] n48025;
wire     [31:0] n48026;
wire     [31:0] n48027;
wire     [31:0] n48028;
wire     [31:0] n48029;
wire     [31:0] n48030;
wire     [31:0] n48031;
wire     [31:0] n48032;
wire     [31:0] n48033;
wire     [31:0] n48034;
wire     [31:0] n48035;
wire     [31:0] n48036;
wire     [31:0] n48037;
wire     [31:0] n48038;
wire     [31:0] n48039;
wire     [31:0] n48040;
wire     [31:0] n48041;
wire     [31:0] n48042;
wire     [31:0] n48043;
wire     [31:0] n48044;
wire     [31:0] n48045;
wire     [31:0] n48046;
wire     [31:0] n48047;
wire     [31:0] n48048;
wire     [31:0] n48049;
wire     [31:0] n48050;
wire     [31:0] n48051;
wire     [31:0] n48052;
wire     [31:0] n48053;
wire     [31:0] n48054;
wire     [31:0] n48055;
wire     [31:0] n48056;
wire     [31:0] n48057;
wire     [31:0] n48058;
wire     [31:0] n48059;
wire     [31:0] n48060;
wire     [31:0] n48061;
wire     [31:0] n48062;
wire     [31:0] n48063;
wire     [31:0] n48064;
wire     [31:0] n48065;
wire     [31:0] n48066;
wire     [31:0] n48067;
wire     [31:0] n48068;
wire     [31:0] n48069;
wire     [31:0] n48070;
wire     [31:0] n48071;
wire     [31:0] n48072;
wire     [31:0] n48073;
wire     [31:0] n48074;
wire     [31:0] n48075;
wire     [31:0] n48076;
wire     [31:0] n48077;
wire     [31:0] n48078;
wire     [31:0] n48079;
wire     [31:0] n48080;
wire     [31:0] n48081;
wire     [31:0] n48082;
wire     [31:0] n48083;
wire     [31:0] n48084;
wire     [31:0] n48085;
wire     [31:0] n48086;
wire     [31:0] n48087;
wire     [31:0] n48088;
wire     [31:0] n48089;
wire     [31:0] n48090;
wire     [31:0] n48091;
wire     [31:0] n48092;
wire     [31:0] n48093;
wire     [31:0] n48094;
wire     [31:0] n48095;
wire     [31:0] n48096;
wire     [31:0] n48097;
wire     [31:0] n48098;
wire     [31:0] n48099;
wire     [31:0] n48100;
wire     [31:0] n48101;
wire     [31:0] n48102;
wire     [31:0] n48103;
wire     [31:0] n48104;
wire     [31:0] n48105;
wire     [31:0] n48106;
wire     [31:0] n48107;
wire     [31:0] n48108;
wire     [31:0] n48109;
wire     [31:0] n48110;
wire     [31:0] n48111;
wire     [31:0] n48112;
wire     [31:0] n48113;
wire     [31:0] n48114;
wire     [31:0] n48115;
wire     [31:0] n48116;
wire     [31:0] n48117;
wire     [31:0] n48118;
wire     [31:0] n48119;
wire     [31:0] n48120;
wire     [31:0] n48121;
wire     [31:0] n48122;
wire     [31:0] n48123;
wire     [31:0] n48124;
wire     [31:0] n48125;
wire     [31:0] n48126;
wire     [31:0] n48127;
wire     [31:0] n48128;
wire     [31:0] n48129;
wire     [31:0] n48130;
wire     [31:0] n48131;
wire     [31:0] n48132;
wire     [31:0] n48133;
wire     [31:0] n48134;
wire     [31:0] n48135;
wire     [31:0] n48136;
wire     [31:0] n48137;
wire     [31:0] n48138;
wire     [31:0] n48139;
wire     [31:0] n48140;
wire     [31:0] n48141;
wire     [31:0] n48142;
wire     [31:0] n48143;
wire     [31:0] n48144;
wire     [31:0] n48145;
wire     [31:0] n48146;
wire     [31:0] n48147;
wire     [31:0] n48148;
wire     [31:0] n48149;
wire     [31:0] n48150;
wire     [31:0] n48151;
wire     [31:0] n48152;
wire     [31:0] n48153;
wire     [31:0] n48154;
wire     [31:0] n48155;
wire     [31:0] n48156;
wire     [31:0] n48157;
wire     [31:0] n48158;
wire     [31:0] n48159;
wire     [31:0] n48160;
wire     [31:0] n48161;
wire     [31:0] n48162;
wire     [31:0] n48163;
wire     [31:0] n48164;
wire     [31:0] n48165;
wire     [31:0] n48166;
wire     [31:0] n48167;
wire     [31:0] n48168;
wire     [31:0] n48169;
wire     [31:0] n48170;
wire     [31:0] n48171;
wire     [31:0] n48172;
wire     [31:0] n48173;
wire     [31:0] n48174;
wire     [31:0] n48175;
wire     [31:0] n48176;
wire     [31:0] n48177;
wire     [31:0] n48178;
wire     [31:0] n48179;
wire     [31:0] n48180;
wire     [31:0] n48181;
wire     [31:0] n48182;
wire     [31:0] n48183;
wire     [31:0] n48184;
wire     [31:0] n48185;
wire     [31:0] n48186;
wire     [31:0] n48187;
wire     [31:0] n48188;
wire     [31:0] n48189;
wire     [31:0] n48190;
wire     [31:0] n48191;
wire     [31:0] n48192;
wire     [31:0] n48193;
wire     [31:0] n48194;
wire     [31:0] n48195;
wire     [31:0] n48196;
wire     [31:0] n48197;
wire     [31:0] n48198;
wire     [31:0] n48199;
wire     [31:0] n48200;
wire     [31:0] n48201;
wire     [31:0] n48202;
wire     [31:0] n48203;
wire     [31:0] n48204;
wire     [31:0] n48205;
wire     [31:0] n48206;
wire     [31:0] n48207;
wire     [31:0] n48208;
wire     [31:0] n48209;
wire     [31:0] n48210;
wire     [31:0] n48211;
wire     [31:0] n48212;
wire     [31:0] n48213;
wire     [31:0] n48214;
wire     [31:0] n48215;
wire     [31:0] n48216;
wire     [31:0] n48217;
wire     [31:0] n48218;
wire     [31:0] n48219;
wire     [31:0] n48220;
wire     [31:0] n48221;
wire     [31:0] n48222;
wire     [31:0] n48223;
wire     [31:0] n48224;
wire     [31:0] n48225;
wire     [31:0] n48226;
wire     [31:0] n48227;
wire     [31:0] n48228;
wire     [31:0] n48229;
wire     [31:0] n48230;
wire     [31:0] n48231;
wire     [31:0] n48232;
wire     [31:0] n48233;
wire     [31:0] n48234;
wire     [31:0] n48235;
wire     [31:0] n48236;
wire     [31:0] n48237;
wire     [31:0] n48238;
wire     [31:0] n48239;
wire     [31:0] n48240;
wire     [31:0] n48241;
wire     [31:0] n48242;
wire     [31:0] n48243;
wire     [31:0] n48244;
wire     [31:0] n48245;
wire     [31:0] n48246;
wire     [31:0] n48247;
wire     [31:0] n48248;
wire     [31:0] n48249;
wire     [31:0] n48250;
wire     [31:0] n48251;
wire     [31:0] n48252;
wire     [31:0] n48253;
wire     [31:0] n48254;
wire     [31:0] n48255;
wire     [31:0] n48256;
wire     [31:0] n48257;
wire     [31:0] n48258;
wire     [31:0] n48259;
wire     [31:0] n48260;
wire     [31:0] n48261;
wire     [31:0] n48262;
wire     [31:0] n48263;
wire     [31:0] n48264;
wire     [31:0] n48265;
wire     [31:0] n48266;
wire     [31:0] n48267;
wire     [31:0] n48268;
wire     [31:0] n48269;
wire     [31:0] n48270;
wire     [31:0] n48271;
wire     [31:0] n48272;
wire     [31:0] n48273;
wire     [31:0] n48274;
wire     [31:0] n48275;
wire     [31:0] n48276;
wire     [31:0] n48277;
wire     [31:0] n48278;
wire     [31:0] n48279;
wire     [31:0] n48280;
wire     [31:0] n48281;
wire     [31:0] n48282;
wire     [31:0] n48283;
wire     [31:0] n48284;
wire     [31:0] n48285;
wire     [31:0] n48286;
wire     [31:0] n48287;
wire     [31:0] n48288;
wire     [31:0] n48289;
wire     [31:0] n48290;
wire     [31:0] n48291;
wire     [31:0] n48292;
wire     [31:0] n48293;
wire     [31:0] n48294;
wire     [31:0] n48295;
wire     [31:0] n48296;
wire     [31:0] n48297;
wire     [31:0] n48298;
wire     [31:0] n48299;
wire     [31:0] n48300;
wire     [31:0] n48301;
wire     [31:0] n48302;
wire     [31:0] n48303;
wire     [31:0] n48304;
wire     [31:0] n48305;
wire     [31:0] n48306;
wire     [31:0] n48307;
wire     [31:0] n48308;
wire     [31:0] n48309;
wire     [31:0] n48310;
wire     [31:0] n48311;
wire     [31:0] n48312;
wire     [31:0] n48313;
wire     [31:0] n48314;
wire     [31:0] n48315;
wire     [31:0] n48316;
wire     [31:0] n48317;
wire     [31:0] n48318;
wire     [31:0] n48319;
wire     [31:0] n48320;
wire     [31:0] n48321;
wire     [31:0] n48322;
wire     [31:0] n48323;
wire     [31:0] n48324;
wire     [31:0] n48325;
wire     [31:0] n48326;
wire     [31:0] n48327;
wire     [31:0] n48328;
wire     [31:0] n48329;
wire     [31:0] n48330;
wire     [31:0] n48331;
wire     [31:0] n48332;
wire     [31:0] n48333;
wire     [31:0] n48334;
wire     [31:0] n48335;
wire     [31:0] n48336;
wire     [31:0] n48337;
wire     [31:0] n48338;
wire     [31:0] n48339;
wire     [31:0] n48340;
wire     [31:0] n48341;
wire     [31:0] n48342;
wire     [31:0] n48343;
wire     [31:0] n48344;
wire     [31:0] n48345;
wire     [31:0] n48346;
wire     [31:0] n48347;
wire     [31:0] n48348;
wire     [31:0] n48349;
wire     [31:0] n48350;
wire     [31:0] n48351;
wire     [31:0] n48352;
wire     [31:0] n48353;
wire     [31:0] n48354;
wire     [31:0] n48355;
wire     [31:0] n48356;
wire     [31:0] n48357;
wire     [31:0] n48358;
wire     [31:0] n48359;
wire     [31:0] n48360;
wire     [31:0] n48361;
wire     [31:0] n48362;
wire     [31:0] n48363;
wire     [31:0] n48364;
wire     [31:0] n48365;
wire     [31:0] n48366;
wire     [31:0] n48367;
wire     [31:0] n48368;
wire     [31:0] n48369;
wire     [31:0] n48370;
wire     [31:0] n48371;
wire     [31:0] n48372;
wire     [31:0] n48373;
wire     [31:0] n48374;
wire     [31:0] n48375;
wire     [31:0] n48376;
wire     [31:0] n48377;
wire     [31:0] n48378;
wire     [31:0] n48379;
wire     [31:0] n48380;
wire     [31:0] n48381;
wire     [31:0] n48382;
wire     [31:0] n48383;
wire     [31:0] n48384;
wire     [31:0] n48385;
wire     [31:0] n48386;
wire     [31:0] n48387;
wire     [31:0] n48388;
wire     [31:0] n48389;
wire     [31:0] n48390;
wire     [31:0] n48391;
wire     [31:0] n48392;
wire     [31:0] n48393;
wire     [31:0] n48394;
wire     [31:0] n48395;
wire     [31:0] n48396;
wire     [31:0] n48397;
wire     [31:0] n48398;
wire     [31:0] n48399;
wire     [31:0] n48400;
wire     [31:0] n48401;
wire     [31:0] n48402;
wire     [31:0] n48403;
wire     [31:0] n48404;
wire     [31:0] n48405;
wire     [31:0] n48406;
wire     [31:0] n48407;
wire     [31:0] n48408;
wire     [31:0] n48409;
wire     [31:0] n48410;
wire     [31:0] n48411;
wire     [31:0] n48412;
wire     [31:0] n48413;
wire     [31:0] n48414;
wire     [31:0] n48415;
wire     [31:0] n48416;
wire     [31:0] n48417;
wire     [31:0] n48418;
wire     [31:0] n48419;
wire     [31:0] n48420;
wire     [31:0] n48421;
wire     [31:0] n48422;
wire     [31:0] n48423;
wire     [31:0] n48424;
wire     [31:0] n48425;
wire     [31:0] n48426;
wire     [31:0] n48427;
wire     [31:0] n48428;
wire     [31:0] n48429;
wire     [31:0] n48430;
wire     [31:0] n48431;
wire     [31:0] n48432;
wire     [31:0] n48433;
wire     [31:0] n48434;
wire     [31:0] n48435;
wire     [31:0] n48436;
wire     [31:0] n48437;
wire     [31:0] n48438;
wire     [31:0] n48439;
wire     [31:0] n48440;
wire     [31:0] n48441;
wire     [31:0] n48442;
wire     [31:0] n48443;
wire     [31:0] n48444;
wire     [31:0] n48445;
wire     [31:0] n48446;
wire     [31:0] n48447;
wire     [31:0] n48448;
wire     [31:0] n48449;
wire     [31:0] n48450;
wire     [31:0] n48451;
wire     [31:0] n48452;
wire     [31:0] n48453;
wire     [31:0] n48454;
wire     [31:0] n48455;
wire     [31:0] n48456;
wire     [31:0] n48457;
wire     [31:0] n48458;
wire     [31:0] n48459;
wire     [31:0] n48460;
wire     [31:0] n48461;
wire     [31:0] n48462;
wire     [31:0] n48463;
wire     [31:0] n48464;
wire     [31:0] n48465;
wire     [31:0] n48466;
wire     [31:0] n48467;
wire     [31:0] n48468;
wire     [31:0] n48469;
wire     [31:0] n48470;
wire     [31:0] n48471;
wire     [31:0] n48472;
wire     [31:0] n48473;
wire     [31:0] n48474;
wire     [31:0] n48475;
wire     [31:0] n48476;
wire     [31:0] n48477;
wire     [31:0] n48478;
wire     [31:0] n48479;
wire     [31:0] n48480;
wire     [31:0] n48481;
wire     [31:0] n48482;
wire     [31:0] n48483;
wire     [31:0] n48484;
wire     [31:0] n48485;
wire     [31:0] n48486;
wire     [31:0] n48487;
wire     [31:0] n48488;
wire     [31:0] n48489;
wire     [31:0] n48490;
wire     [31:0] n48491;
wire     [31:0] n48492;
wire     [31:0] n48493;
wire     [31:0] n48494;
wire     [31:0] n48495;
wire     [31:0] n48496;
wire     [31:0] n48497;
wire     [31:0] n48498;
wire     [31:0] n48499;
wire     [31:0] n48500;
wire     [31:0] n48501;
wire     [31:0] n48502;
wire     [31:0] n48503;
wire     [31:0] n48504;
wire     [31:0] n48505;
wire     [31:0] n48506;
wire     [31:0] n48507;
wire     [31:0] n48508;
wire     [31:0] n48509;
wire     [31:0] n48510;
wire     [31:0] n48511;
wire     [31:0] n48512;
wire     [31:0] n48513;
wire     [31:0] n48514;
wire     [31:0] n48515;
wire     [31:0] n48516;
wire     [31:0] n48517;
wire     [31:0] n48518;
wire     [31:0] n48519;
wire     [31:0] n48520;
wire     [31:0] n48521;
wire     [31:0] n48522;
wire     [31:0] n48523;
wire     [31:0] n48524;
wire     [31:0] n48525;
wire     [31:0] n48526;
wire     [31:0] n48527;
wire     [31:0] n48528;
wire     [31:0] n48529;
wire     [31:0] n48530;
wire     [31:0] n48531;
wire     [31:0] n48532;
wire     [31:0] n48533;
wire     [31:0] n48534;
wire     [31:0] n48535;
wire     [31:0] n48536;
wire     [31:0] n48537;
wire     [31:0] n48538;
wire     [31:0] n48539;
wire     [31:0] n48540;
wire     [31:0] n48541;
wire     [31:0] n48542;
wire     [31:0] n48543;
wire     [31:0] n48544;
wire     [31:0] n48545;
wire     [31:0] n48546;
wire     [31:0] n48547;
wire     [31:0] n48548;
wire     [31:0] n48549;
wire     [31:0] n48550;
wire     [31:0] n48551;
wire     [31:0] n48552;
wire     [31:0] n48553;
wire     [31:0] n48554;
wire     [31:0] n48555;
wire     [31:0] n48556;
wire     [31:0] n48557;
wire     [31:0] n48558;
wire     [31:0] n48559;
wire     [31:0] n48560;
wire     [31:0] n48561;
wire     [31:0] n48562;
wire     [31:0] n48563;
wire     [31:0] n48564;
wire     [31:0] n48565;
wire     [31:0] n48566;
wire     [31:0] n48567;
wire     [31:0] n48568;
wire     [31:0] n48569;
wire     [31:0] n48570;
wire     [31:0] n48571;
wire     [31:0] n48572;
wire     [31:0] n48573;
wire     [31:0] n48574;
wire     [31:0] n48575;
wire     [31:0] n48576;
wire     [31:0] n48577;
wire     [31:0] n48578;
wire     [31:0] n48579;
wire     [31:0] n48580;
wire     [31:0] n48581;
wire     [31:0] n48582;
wire     [31:0] n48583;
wire     [31:0] n48584;
wire     [31:0] n48585;
wire     [31:0] n48586;
wire     [31:0] n48587;
wire     [31:0] n48588;
wire     [31:0] n48589;
wire     [31:0] n48590;
wire     [31:0] n48591;
wire     [31:0] n48592;
wire     [31:0] n48593;
wire     [31:0] n48594;
wire     [31:0] n48595;
wire     [31:0] n48596;
wire     [31:0] n48597;
wire     [31:0] n48598;
wire     [31:0] n48599;
wire     [31:0] n48600;
wire     [31:0] n48601;
wire     [31:0] n48602;
wire     [31:0] n48603;
wire     [31:0] n48604;
wire     [31:0] n48605;
wire     [31:0] n48606;
wire     [31:0] n48607;
wire     [31:0] n48608;
wire     [31:0] n48609;
wire     [31:0] n48610;
wire     [31:0] n48611;
wire     [31:0] n48612;
wire     [31:0] n48613;
wire     [31:0] n48614;
wire     [31:0] n48615;
wire     [31:0] n48616;
wire     [31:0] n48617;
wire     [31:0] n48618;
wire     [31:0] n48619;
wire     [31:0] n48620;
wire     [31:0] n48621;
wire     [31:0] n48622;
wire     [31:0] n48623;
wire     [31:0] n48624;
wire     [31:0] n48625;
wire     [31:0] n48626;
wire     [31:0] n48627;
wire     [31:0] n48628;
wire     [31:0] n48629;
wire     [31:0] n48630;
wire     [31:0] n48631;
wire     [31:0] n48632;
wire     [31:0] n48633;
wire     [31:0] n48634;
wire     [31:0] n48635;
wire     [31:0] n48636;
wire     [31:0] n48637;
wire     [31:0] n48638;
wire     [31:0] n48639;
wire     [31:0] n48640;
wire     [31:0] n48641;
wire     [31:0] n48642;
wire     [31:0] n48643;
wire     [31:0] n48644;
wire     [31:0] n48645;
wire     [31:0] n48646;
wire     [31:0] n48647;
wire     [31:0] n48648;
wire     [31:0] n48649;
wire     [31:0] n48650;
wire     [31:0] n48651;
wire     [31:0] n48652;
wire     [31:0] n48653;
wire     [31:0] n48654;
wire     [31:0] n48655;
wire     [31:0] n48656;
wire     [31:0] n48657;
wire     [31:0] n48658;
wire     [31:0] n48659;
wire     [31:0] n48660;
wire     [31:0] n48661;
wire     [31:0] n48662;
wire     [31:0] n48663;
wire     [31:0] n48664;
wire     [31:0] n48665;
wire     [31:0] n48666;
wire     [31:0] n48667;
wire     [31:0] n48668;
wire     [31:0] n48669;
wire     [31:0] n48670;
wire     [31:0] n48671;
wire     [31:0] n48672;
wire     [31:0] n48673;
wire     [31:0] n48674;
wire     [31:0] n48675;
wire     [31:0] n48676;
wire     [31:0] n48677;
wire     [31:0] n48678;
wire     [31:0] n48679;
wire     [31:0] n48680;
wire     [31:0] n48681;
wire     [31:0] n48682;
wire     [31:0] n48683;
wire     [31:0] n48684;
wire     [31:0] n48685;
wire     [31:0] n48686;
wire     [31:0] n48687;
wire     [31:0] n48688;
wire     [31:0] n48689;
wire     [31:0] n48690;
wire     [31:0] n48691;
wire     [31:0] n48692;
wire     [31:0] n48693;
wire     [31:0] n48694;
wire     [31:0] n48695;
wire     [31:0] n48696;
wire     [31:0] n48697;
wire     [31:0] n48698;
wire     [31:0] n48699;
wire     [31:0] n48700;
wire     [31:0] n48701;
wire     [31:0] n48702;
wire     [31:0] n48703;
wire     [31:0] n48704;
wire     [31:0] n48705;
wire     [31:0] n48706;
wire     [31:0] n48707;
wire     [31:0] n48708;
wire     [31:0] n48709;
wire     [31:0] n48710;
wire     [31:0] n48711;
wire     [31:0] n48712;
wire     [31:0] n48713;
wire     [31:0] n48714;
wire     [31:0] n48715;
wire     [31:0] n48716;
wire     [31:0] n48717;
wire     [31:0] n48718;
wire     [31:0] n48719;
wire     [31:0] n48720;
wire     [31:0] n48721;
wire     [31:0] n48722;
wire     [31:0] n48723;
wire     [31:0] n48724;
wire     [31:0] n48725;
wire     [31:0] n48726;
wire     [31:0] n48727;
wire     [31:0] n48728;
wire     [31:0] n48729;
wire     [31:0] n48730;
wire     [31:0] n48731;
wire     [31:0] n48732;
wire     [31:0] n48733;
wire     [31:0] n48734;
wire     [31:0] n48735;
wire     [31:0] n48736;
wire     [31:0] n48737;
wire     [31:0] n48738;
wire     [31:0] n48739;
wire     [31:0] n48740;
wire     [31:0] n48741;
wire     [31:0] n48742;
wire     [31:0] n48743;
wire     [31:0] n48744;
wire     [31:0] n48745;
wire     [31:0] n48746;
wire     [31:0] n48747;
wire     [31:0] n48748;
wire     [31:0] n48749;
wire     [31:0] n48750;
wire     [31:0] n48751;
wire     [31:0] n48752;
wire     [31:0] n48753;
wire     [31:0] n48754;
wire     [31:0] n48755;
wire     [31:0] n48756;
wire     [31:0] n48757;
wire     [31:0] n48758;
wire     [31:0] n48759;
wire     [31:0] n48760;
wire     [31:0] n48761;
wire     [31:0] n48762;
wire     [31:0] n48763;
wire     [31:0] n48764;
wire     [31:0] n48765;
wire     [31:0] n48766;
wire     [31:0] n48767;
wire     [31:0] n48768;
wire     [31:0] n48769;
wire     [31:0] n48770;
wire     [31:0] n48771;
wire     [31:0] n48772;
wire     [31:0] n48773;
wire     [31:0] n48774;
wire     [31:0] n48775;
wire     [31:0] n48776;
wire     [31:0] n48777;
wire     [31:0] n48778;
wire     [31:0] n48779;
wire     [31:0] n48780;
wire     [31:0] n48781;
wire     [31:0] n48782;
wire     [31:0] n48783;
wire     [31:0] n48784;
wire     [31:0] n48785;
wire     [31:0] n48786;
wire     [31:0] n48787;
wire     [31:0] n48788;
wire     [31:0] n48789;
wire     [31:0] n48790;
wire     [31:0] n48791;
wire     [31:0] n48792;
wire     [31:0] n48793;
wire     [31:0] n48794;
wire     [31:0] n48795;
wire     [31:0] n48796;
wire     [31:0] n48797;
wire     [31:0] n48798;
wire     [31:0] n48799;
wire     [31:0] n48800;
wire     [31:0] n48801;
wire     [31:0] n48802;
wire     [31:0] n48803;
wire     [31:0] n48804;
wire     [31:0] n48805;
wire     [31:0] n48806;
wire     [31:0] n48807;
wire     [31:0] n48808;
wire     [31:0] n48809;
wire     [31:0] n48810;
wire     [31:0] n48811;
wire     [31:0] n48812;
wire     [31:0] n48813;
wire     [31:0] n48814;
wire     [31:0] n48815;
wire     [31:0] n48816;
wire     [31:0] n48817;
wire     [31:0] n48818;
wire     [31:0] n48819;
wire     [31:0] n48820;
wire     [31:0] n48821;
wire     [31:0] n48822;
wire     [31:0] n48823;
wire     [31:0] n48824;
wire     [31:0] n48825;
wire     [31:0] n48826;
wire     [31:0] n48827;
wire     [31:0] n48828;
wire     [31:0] n48829;
wire     [31:0] n48830;
wire     [31:0] n48831;
wire     [31:0] n48832;
wire     [31:0] n48833;
wire     [31:0] n48834;
wire     [31:0] n48835;
wire     [31:0] n48836;
wire     [31:0] n48837;
wire     [31:0] n48838;
wire     [31:0] n48839;
wire     [31:0] n48840;
wire     [31:0] n48841;
wire     [31:0] n48842;
wire     [31:0] n48843;
wire     [31:0] n48844;
wire     [31:0] n48845;
wire     [31:0] n48846;
wire     [31:0] n48847;
wire     [31:0] n48848;
wire     [31:0] n48849;
wire     [31:0] n48850;
wire     [31:0] n48851;
wire     [31:0] n48852;
wire     [31:0] n48853;
wire     [31:0] n48854;
wire     [31:0] n48855;
wire     [31:0] n48856;
wire     [31:0] n48857;
wire     [31:0] n48858;
wire     [31:0] n48859;
wire     [31:0] n48860;
wire     [31:0] n48861;
wire     [31:0] n48862;
wire     [31:0] n48863;
wire     [31:0] n48864;
wire     [31:0] n48865;
wire     [31:0] n48866;
wire     [31:0] n48867;
wire     [31:0] n48868;
wire     [31:0] n48869;
wire     [31:0] n48870;
wire     [31:0] n48871;
wire     [31:0] n48872;
wire     [31:0] n48873;
wire     [31:0] n48874;
wire     [31:0] n48875;
wire     [31:0] n48876;
wire     [31:0] n48877;
wire     [31:0] n48878;
wire     [31:0] n48879;
wire     [31:0] n48880;
wire     [31:0] n48881;
wire     [31:0] n48882;
wire     [31:0] n48883;
wire     [31:0] n48884;
wire     [31:0] n48885;
wire     [31:0] n48886;
wire     [31:0] n48887;
wire     [31:0] n48888;
wire     [31:0] n48889;
wire     [31:0] n48890;
wire     [31:0] n48891;
wire     [31:0] n48892;
wire     [31:0] n48893;
wire     [31:0] n48894;
wire     [31:0] n48895;
wire     [31:0] n48896;
wire     [31:0] n48897;
wire     [31:0] n48898;
wire     [31:0] n48899;
wire     [31:0] n48900;
wire     [31:0] n48901;
wire     [31:0] n48902;
wire     [31:0] n48903;
wire     [31:0] n48904;
wire     [31:0] n48905;
wire     [31:0] n48906;
wire     [31:0] n48907;
wire     [31:0] n48908;
wire     [31:0] n48909;
wire     [31:0] n48910;
wire     [31:0] n48911;
wire     [31:0] n48912;
wire     [31:0] n48913;
wire     [31:0] n48914;
wire     [31:0] n48915;
wire     [31:0] n48916;
wire     [31:0] n48917;
wire     [31:0] n48918;
wire     [31:0] n48919;
wire     [31:0] n48920;
wire     [31:0] n48921;
wire     [31:0] n48922;
wire     [31:0] n48923;
wire     [31:0] n48924;
wire     [31:0] n48925;
wire     [31:0] n48926;
wire     [31:0] n48927;
wire     [31:0] n48928;
wire     [31:0] n48929;
wire     [31:0] n48930;
wire     [31:0] n48931;
wire     [31:0] n48932;
wire     [31:0] n48933;
wire     [31:0] n48934;
wire     [31:0] n48935;
wire     [31:0] n48936;
wire     [31:0] n48937;
wire     [31:0] n48938;
wire     [31:0] n48939;
wire     [31:0] n48940;
wire     [31:0] n48941;
wire     [31:0] n48942;
wire     [31:0] n48943;
wire     [31:0] n48944;
wire     [31:0] n48945;
wire     [31:0] n48946;
wire     [31:0] n48947;
wire     [31:0] n48948;
wire     [31:0] n48949;
wire     [31:0] n48950;
wire     [31:0] n48951;
wire     [31:0] n48952;
wire     [31:0] n48953;
wire     [31:0] n48954;
wire     [31:0] n48955;
wire     [31:0] n48956;
wire     [31:0] n48957;
wire     [31:0] n48958;
wire     [31:0] n48959;
wire     [31:0] n48960;
wire     [31:0] n48961;
wire     [31:0] n48962;
wire     [31:0] n48963;
wire     [31:0] n48964;
wire     [31:0] n48965;
wire     [31:0] n48966;
wire     [31:0] n48967;
wire     [31:0] n48968;
wire     [31:0] n48969;
wire     [31:0] n48970;
wire     [31:0] n48971;
wire     [31:0] n48972;
wire     [31:0] n48973;
wire     [31:0] n48974;
wire     [31:0] n48975;
wire     [31:0] n48976;
wire     [31:0] n48977;
wire     [31:0] n48978;
wire     [31:0] n48979;
wire     [31:0] n48980;
wire     [31:0] n48981;
wire     [31:0] n48982;
wire     [31:0] n48983;
wire     [31:0] n48984;
wire     [31:0] n48985;
wire     [31:0] n48986;
wire     [31:0] n48987;
wire     [31:0] n48988;
wire     [31:0] n48989;
wire     [31:0] n48990;
wire     [31:0] n48991;
wire     [31:0] n48992;
wire     [31:0] n48993;
wire     [31:0] n48994;
wire     [31:0] n48995;
wire     [31:0] n48996;
wire     [31:0] n48997;
wire     [31:0] n48998;
wire     [31:0] n48999;
wire     [31:0] n49000;
wire     [31:0] n49001;
wire     [31:0] n49002;
wire     [31:0] n49003;
wire     [31:0] n49004;
wire     [31:0] n49005;
wire     [31:0] n49006;
wire     [31:0] n49007;
wire     [31:0] n49008;
wire     [31:0] n49009;
wire     [31:0] n49010;
wire     [31:0] n49011;
wire     [31:0] n49012;
wire     [31:0] n49013;
wire     [31:0] n49014;
wire     [31:0] n49015;
wire     [31:0] n49016;
wire     [31:0] n49017;
wire     [31:0] n49018;
wire     [31:0] n49019;
wire     [31:0] n49020;
wire     [31:0] n49021;
wire     [31:0] n49022;
wire     [31:0] n49023;
wire     [31:0] n49024;
wire     [31:0] n49025;
wire     [31:0] n49026;
wire     [31:0] n49027;
wire     [31:0] n49028;
wire     [31:0] n49029;
wire     [31:0] n49030;
wire     [31:0] n49031;
wire     [31:0] n49032;
wire     [31:0] n49033;
wire     [31:0] n49034;
wire     [31:0] n49035;
wire     [31:0] n49036;
wire     [31:0] n49037;
wire     [31:0] n49038;
wire     [31:0] n49039;
wire     [31:0] n49040;
wire     [31:0] n49041;
wire     [31:0] n49042;
wire     [31:0] n49043;
wire     [31:0] n49044;
wire     [31:0] n49045;
wire     [31:0] n49046;
wire     [31:0] n49047;
wire     [31:0] n49048;
wire     [31:0] n49049;
wire     [31:0] n49050;
wire     [31:0] n49051;
wire     [31:0] n49052;
wire     [31:0] n49053;
wire     [31:0] n49054;
wire     [31:0] n49055;
wire     [31:0] n49056;
wire     [31:0] n49057;
wire     [31:0] n49058;
wire     [31:0] n49059;
wire     [31:0] n49060;
wire     [31:0] n49061;
wire     [31:0] n49062;
wire     [31:0] n49063;
wire     [31:0] n49064;
wire     [31:0] n49065;
wire     [31:0] n49066;
wire     [31:0] n49067;
wire     [31:0] n49068;
wire     [31:0] n49069;
wire     [31:0] n49070;
wire     [31:0] n49071;
wire     [31:0] n49072;
wire     [31:0] n49073;
wire     [31:0] n49074;
wire     [31:0] n49075;
wire     [31:0] n49076;
wire     [31:0] n49077;
wire     [31:0] n49078;
wire     [31:0] n49079;
wire     [31:0] n49080;
wire     [31:0] n49081;
wire     [31:0] n49082;
wire     [31:0] n49083;
wire     [31:0] n49084;
wire     [31:0] n49085;
wire     [31:0] n49086;
wire     [31:0] n49087;
wire     [31:0] n49088;
wire     [31:0] n49089;
wire     [31:0] n49090;
wire     [31:0] n49091;
wire     [31:0] n49092;
wire     [31:0] n49093;
wire     [31:0] n49094;
wire     [31:0] n49095;
wire     [31:0] n49096;
wire     [31:0] n49097;
wire     [31:0] n49098;
wire     [31:0] n49099;
wire     [31:0] n49100;
wire     [31:0] n49101;
wire     [31:0] n49102;
wire     [31:0] n49103;
wire     [31:0] n49104;
wire     [31:0] n49105;
wire     [31:0] n49106;
wire     [31:0] n49107;
wire     [31:0] n49108;
wire     [31:0] n49109;
wire     [31:0] n49110;
wire     [31:0] n49111;
wire     [31:0] n49112;
wire     [31:0] n49113;
wire     [31:0] n49114;
wire     [31:0] n49115;
wire     [31:0] n49116;
wire     [31:0] n49117;
wire     [31:0] n49118;
wire     [31:0] n49119;
wire     [31:0] n49120;
wire     [31:0] n49121;
wire     [31:0] n49122;
wire     [31:0] n49123;
wire     [31:0] n49124;
wire     [31:0] n49125;
wire     [31:0] n49126;
wire     [31:0] n49127;
wire     [31:0] n49128;
wire     [31:0] n49129;
wire     [31:0] n49130;
wire     [31:0] n49131;
wire     [31:0] n49132;
wire     [31:0] n49133;
wire     [31:0] n49134;
wire     [31:0] n49135;
wire     [31:0] n49136;
wire     [31:0] n49137;
wire     [31:0] n49138;
wire     [31:0] n49139;
wire     [31:0] n49140;
wire     [31:0] n49141;
wire     [31:0] n49142;
wire     [31:0] n49143;
wire     [31:0] n49144;
wire     [31:0] n49145;
wire     [31:0] n49146;
wire     [31:0] n49147;
wire     [31:0] n49148;
wire     [31:0] n49149;
wire     [31:0] n49150;
wire     [31:0] n49151;
wire     [31:0] n49152;
wire     [31:0] n49153;
wire     [31:0] n49154;
wire     [31:0] n49155;
wire     [31:0] n49156;
wire     [31:0] n49157;
wire     [31:0] n49158;
wire     [31:0] n49159;
wire     [31:0] n49160;
wire     [31:0] n49161;
wire     [31:0] n49162;
wire     [31:0] n49163;
wire     [31:0] n49164;
wire     [31:0] n49165;
wire     [31:0] n49166;
wire     [31:0] n49167;
wire     [31:0] n49168;
wire     [31:0] n49169;
wire     [31:0] n49170;
wire     [31:0] n49171;
wire     [31:0] n49172;
wire     [31:0] n49173;
wire     [31:0] n49174;
wire     [31:0] n49175;
wire     [31:0] n49176;
wire     [31:0] n49177;
wire     [31:0] n49178;
wire     [31:0] n49179;
wire     [31:0] n49180;
wire     [31:0] n49181;
wire     [31:0] n49182;
wire     [31:0] n49183;
wire     [31:0] n49184;
wire     [31:0] n49185;
wire     [31:0] n49186;
wire     [31:0] n49187;
wire     [31:0] n49188;
wire     [31:0] n49189;
wire     [31:0] n49190;
wire     [31:0] n49191;
wire     [31:0] n49192;
wire     [31:0] n49193;
wire     [31:0] n49194;
wire     [31:0] n49195;
wire     [31:0] n49196;
wire     [31:0] n49197;
wire     [31:0] n49198;
wire     [31:0] n49199;
wire     [31:0] n49200;
wire     [31:0] n49201;
wire     [31:0] n49202;
wire     [31:0] n49203;
wire     [31:0] n49204;
wire     [31:0] n49205;
wire     [31:0] n49206;
wire     [31:0] n49207;
wire     [31:0] n49208;
wire     [31:0] n49209;
wire     [31:0] n49210;
wire     [31:0] n49211;
wire     [31:0] n49212;
wire     [31:0] n49213;
wire     [31:0] n49214;
wire     [31:0] n49215;
wire     [31:0] n49216;
wire     [31:0] n49217;
wire     [31:0] n49218;
wire     [31:0] n49219;
wire     [31:0] n49220;
wire     [31:0] n49221;
wire     [31:0] n49222;
wire     [31:0] n49223;
wire     [31:0] n49224;
wire     [31:0] n49225;
wire     [31:0] n49226;
wire     [31:0] n49227;
wire     [31:0] n49228;
wire     [31:0] n49229;
wire     [31:0] n49230;
wire     [31:0] n49231;
wire     [31:0] n49232;
wire     [31:0] n49233;
wire     [31:0] n49234;
wire     [31:0] n49235;
wire     [31:0] n49236;
wire     [31:0] n49237;
wire     [31:0] n49238;
wire     [31:0] n49239;
wire     [31:0] n49240;
wire     [31:0] n49241;
wire     [31:0] n49242;
wire     [31:0] n49243;
wire     [31:0] n49244;
wire     [31:0] n49245;
wire     [31:0] n49246;
wire     [31:0] n49247;
wire     [31:0] n49248;
wire     [31:0] n49249;
wire     [31:0] n49250;
wire     [31:0] n49251;
wire     [31:0] n49252;
wire     [31:0] n49253;
wire     [31:0] n49254;
wire     [31:0] n49255;
wire     [31:0] n49256;
wire     [31:0] n49257;
wire     [31:0] n49258;
wire     [31:0] n49259;
wire     [31:0] n49260;
wire     [31:0] n49261;
wire     [31:0] n49262;
wire     [31:0] n49263;
wire     [31:0] n49264;
wire     [31:0] n49265;
wire     [31:0] n49266;
wire     [31:0] n49267;
wire     [31:0] n49268;
wire     [31:0] n49269;
wire     [31:0] n49270;
wire     [31:0] n49271;
wire     [31:0] n49272;
wire     [31:0] n49273;
wire     [31:0] n49274;
wire     [31:0] n49275;
wire     [31:0] n49276;
wire     [31:0] n49277;
wire     [31:0] n49278;
wire     [31:0] n49279;
wire     [31:0] n49280;
wire     [31:0] n49281;
wire     [31:0] n49282;
wire     [31:0] n49283;
wire     [31:0] n49284;
wire     [31:0] n49285;
wire     [31:0] n49286;
wire     [31:0] n49287;
wire     [31:0] n49288;
wire     [31:0] n49289;
wire     [31:0] n49290;
wire     [31:0] n49291;
wire     [31:0] n49292;
wire     [31:0] n49293;
wire     [31:0] n49294;
wire     [31:0] n49295;
wire     [31:0] n49296;
wire     [31:0] n49297;
wire     [31:0] n49298;
wire     [31:0] n49299;
wire     [31:0] n49300;
wire     [31:0] n49301;
wire     [31:0] n49302;
wire     [31:0] n49303;
wire     [31:0] n49304;
wire     [31:0] n49305;
wire     [31:0] n49306;
wire     [31:0] n49307;
wire     [31:0] n49308;
wire     [31:0] n49309;
wire     [31:0] n49310;
wire     [31:0] n49311;
wire     [31:0] n49312;
wire     [31:0] n49313;
wire     [31:0] n49314;
wire     [31:0] n49315;
wire     [31:0] n49316;
wire     [31:0] n49317;
wire     [31:0] n49318;
wire     [31:0] n49319;
wire     [31:0] n49320;
wire     [31:0] n49321;
wire     [31:0] n49322;
wire     [31:0] n49323;
wire     [31:0] n49324;
wire     [31:0] n49325;
wire     [31:0] n49326;
wire     [31:0] n49327;
wire     [31:0] n49328;
wire     [31:0] n49329;
wire     [31:0] n49330;
wire     [31:0] n49331;
wire     [31:0] n49332;
wire     [31:0] n49333;
wire     [31:0] n49334;
wire     [31:0] n49335;
wire     [31:0] n49336;
wire     [31:0] n49337;
wire     [31:0] n49338;
wire     [31:0] n49339;
wire     [31:0] n49340;
wire     [31:0] n49341;
wire     [31:0] n49342;
wire     [31:0] n49343;
wire     [31:0] n49344;
wire     [31:0] n49345;
wire     [31:0] n49346;
wire     [31:0] n49347;
wire     [31:0] n49348;
wire     [31:0] n49349;
wire     [31:0] n49350;
wire     [31:0] n49351;
wire     [31:0] n49352;
wire     [31:0] n49353;
wire     [31:0] n49354;
wire     [31:0] n49355;
wire     [31:0] n49356;
wire     [31:0] n49357;
wire     [31:0] n49358;
wire     [31:0] n49359;
wire     [31:0] n49360;
wire     [31:0] n49361;
wire     [31:0] n49362;
wire     [31:0] n49363;
wire     [31:0] n49364;
wire     [31:0] n49365;
wire     [31:0] n49366;
wire     [31:0] n49367;
wire     [31:0] n49368;
wire     [31:0] n49369;
wire     [31:0] n49370;
wire     [31:0] n49371;
wire     [31:0] n49372;
wire     [31:0] n49373;
wire     [31:0] n49374;
wire     [31:0] n49375;
wire     [31:0] n49376;
wire     [31:0] n49377;
wire     [31:0] n49378;
wire     [31:0] n49379;
wire     [31:0] n49380;
wire     [31:0] n49381;
wire     [31:0] n49382;
wire     [31:0] n49383;
wire     [31:0] n49384;
wire     [31:0] n49385;
wire     [31:0] n49386;
wire     [31:0] n49387;
wire     [31:0] n49388;
wire     [31:0] n49389;
wire     [31:0] n49390;
wire     [31:0] n49391;
wire     [31:0] n49392;
wire     [31:0] n49393;
wire     [31:0] n49394;
wire     [31:0] n49395;
wire     [31:0] n49396;
wire     [31:0] n49397;
wire     [31:0] n49398;
wire     [31:0] n49399;
wire     [31:0] n49400;
wire     [31:0] n49401;
wire     [31:0] n49402;
wire     [31:0] n49403;
wire     [31:0] n49404;
wire     [31:0] n49405;
wire     [31:0] n49406;
wire     [31:0] n49407;
wire     [31:0] n49408;
wire     [31:0] n49409;
wire     [31:0] n49410;
wire     [31:0] n49411;
wire     [31:0] n49412;
wire     [31:0] n49413;
wire     [31:0] n49414;
wire     [31:0] n49415;
wire     [31:0] n49416;
wire     [31:0] n49417;
wire     [31:0] n49418;
wire     [31:0] n49419;
wire     [31:0] n49420;
wire     [31:0] n49421;
wire     [31:0] n49422;
wire     [31:0] n49423;
wire     [31:0] n49424;
wire     [31:0] n49425;
wire     [31:0] n49426;
wire     [31:0] n49427;
wire     [31:0] n49428;
wire     [31:0] n49429;
wire     [31:0] n49430;
wire     [31:0] n49431;
wire     [31:0] n49432;
wire     [31:0] n49433;
wire     [31:0] n49434;
wire     [31:0] n49435;
wire     [31:0] n49436;
wire     [31:0] n49437;
wire     [31:0] n49438;
wire     [31:0] n49439;
wire     [31:0] n49440;
wire     [31:0] n49441;
wire     [31:0] n49442;
wire     [31:0] n49443;
wire     [31:0] n49444;
wire     [31:0] n49445;
wire     [31:0] n49446;
wire     [31:0] n49447;
wire     [31:0] n49448;
wire     [31:0] n49449;
wire     [31:0] n49450;
wire     [31:0] n49451;
wire     [31:0] n49452;
wire     [31:0] n49453;
wire     [31:0] n49454;
wire     [31:0] n49455;
wire     [31:0] n49456;
wire     [31:0] n49457;
wire     [31:0] n49458;
wire     [31:0] n49459;
wire     [31:0] n49460;
wire     [31:0] n49461;
wire     [31:0] n49462;
wire     [31:0] n49463;
wire     [31:0] n49464;
wire     [31:0] n49465;
wire     [31:0] n49466;
wire     [31:0] n49467;
wire     [31:0] n49468;
wire     [31:0] n49469;
wire     [31:0] n49470;
wire     [31:0] n49471;
wire     [31:0] n49472;
wire     [31:0] n49473;
wire     [31:0] n49474;
wire     [31:0] n49475;
wire     [31:0] n49476;
wire     [31:0] n49477;
wire     [31:0] n49478;
wire     [31:0] n49479;
wire     [31:0] n49480;
wire     [31:0] n49481;
wire     [31:0] n49482;
wire     [31:0] n49483;
wire     [31:0] n49484;
wire     [31:0] n49485;
wire     [31:0] n49486;
wire     [31:0] n49487;
wire     [31:0] n49488;
wire     [31:0] n49489;
wire     [31:0] n49490;
wire     [31:0] n49491;
wire     [31:0] n49492;
wire     [31:0] n49493;
wire     [31:0] n49494;
wire     [31:0] n49495;
wire     [31:0] n49496;
wire     [31:0] n49497;
wire     [31:0] n49498;
wire     [31:0] n49499;
wire     [31:0] n49500;
wire     [31:0] n49501;
wire     [31:0] n49502;
wire     [31:0] n49503;
wire     [31:0] n49504;
wire     [31:0] n49505;
wire     [31:0] n49506;
wire     [31:0] n49507;
wire     [31:0] n49508;
wire     [31:0] n49509;
wire     [31:0] n49510;
wire     [31:0] n49511;
wire     [31:0] n49512;
wire     [31:0] n49513;
wire     [31:0] n49514;
wire     [31:0] n49515;
wire     [31:0] n49516;
wire     [31:0] n49517;
wire     [31:0] n49518;
wire     [31:0] n49519;
wire     [31:0] n49520;
wire     [31:0] n49521;
wire     [31:0] n49522;
wire     [31:0] n49523;
wire     [31:0] n49524;
wire     [31:0] n49525;
wire     [31:0] n49526;
wire     [31:0] n49527;
wire     [31:0] n49528;
wire     [31:0] n49529;
wire     [31:0] n49530;
wire     [31:0] n49531;
wire     [31:0] n49532;
wire     [31:0] n49533;
wire     [31:0] n49534;
wire     [31:0] n49535;
wire     [31:0] n49536;
wire     [31:0] n49537;
wire     [31:0] n49538;
wire     [31:0] n49539;
wire     [31:0] n49540;
wire     [31:0] n49541;
wire     [31:0] n49542;
wire     [31:0] n49543;
wire     [31:0] n49544;
wire     [31:0] n49545;
wire     [31:0] n49546;
wire     [31:0] n49547;
wire     [31:0] n49548;
wire     [31:0] n49549;
wire     [31:0] n49550;
wire     [31:0] n49551;
wire     [31:0] n49552;
wire     [31:0] n49553;
wire     [31:0] n49554;
wire     [31:0] n49555;
wire     [31:0] n49556;
wire     [31:0] n49557;
wire     [31:0] n49558;
wire     [31:0] n49559;
wire     [31:0] n49560;
wire     [31:0] n49561;
wire     [31:0] n49562;
wire     [31:0] n49563;
wire     [31:0] n49564;
wire     [31:0] n49565;
wire     [31:0] n49566;
wire     [31:0] n49567;
wire     [31:0] n49568;
wire     [31:0] n49569;
wire     [31:0] n49570;
wire     [31:0] n49571;
wire     [31:0] n49572;
wire     [31:0] n49573;
wire     [31:0] n49574;
wire     [31:0] n49575;
wire     [31:0] n49576;
wire     [31:0] n49577;
wire     [31:0] n49578;
wire     [31:0] n49579;
wire     [31:0] n49580;
wire     [31:0] n49581;
wire     [31:0] n49582;
wire     [31:0] n49583;
wire     [31:0] n49584;
wire     [31:0] n49585;
wire     [31:0] n49586;
wire     [31:0] n49587;
wire     [31:0] n49588;
wire     [31:0] n49589;
wire     [31:0] n49590;
wire     [31:0] n49591;
wire     [31:0] n49592;
wire     [31:0] n49593;
wire     [31:0] n49594;
wire     [31:0] n49595;
wire     [31:0] n49596;
wire     [31:0] n49597;
wire     [31:0] n49598;
wire     [31:0] n49599;
wire     [31:0] n49600;
wire     [31:0] n49601;
wire     [31:0] n49602;
wire     [31:0] n49603;
wire     [31:0] n49604;
wire     [31:0] n49605;
wire     [31:0] n49606;
wire     [31:0] n49607;
wire     [31:0] n49608;
wire     [31:0] n49609;
wire     [31:0] n49610;
wire     [31:0] n49611;
wire     [31:0] n49612;
wire     [31:0] n49613;
wire     [31:0] n49614;
wire     [31:0] n49615;
wire     [31:0] n49616;
wire     [31:0] n49617;
wire     [31:0] n49618;
wire     [31:0] n49619;
wire     [31:0] n49620;
wire     [31:0] n49621;
wire     [31:0] n49622;
wire     [31:0] n49623;
wire     [31:0] n49624;
wire     [31:0] n49625;
wire     [31:0] n49626;
wire     [31:0] n49627;
wire     [31:0] n49628;
wire     [31:0] n49629;
wire     [31:0] n49630;
wire     [31:0] n49631;
wire     [31:0] n49632;
wire     [31:0] n49633;
wire     [31:0] n49634;
wire     [31:0] n49635;
wire     [31:0] n49636;
wire     [31:0] n49637;
wire     [31:0] n49638;
wire     [31:0] n49639;
wire     [31:0] n49640;
wire     [31:0] n49641;
wire     [31:0] n49642;
wire     [31:0] n49643;
wire     [31:0] n49644;
wire     [31:0] n49645;
wire     [31:0] n49646;
wire     [31:0] n49647;
wire     [31:0] n49648;
wire     [31:0] n49649;
wire     [31:0] n49650;
wire     [31:0] n49651;
wire     [31:0] n49652;
wire     [31:0] n49653;
wire     [31:0] n49654;
wire     [31:0] n49655;
wire     [31:0] n49656;
wire     [31:0] n49657;
wire     [31:0] n49658;
wire     [31:0] n49659;
wire     [31:0] n49660;
wire     [31:0] n49661;
wire     [31:0] n49662;
wire     [31:0] n49663;
wire     [31:0] n49664;
wire     [31:0] n49665;
wire     [31:0] n49666;
wire     [31:0] n49667;
wire     [31:0] n49668;
wire     [31:0] n49669;
wire     [31:0] n49670;
wire     [31:0] n49671;
wire     [31:0] n49672;
wire     [31:0] n49673;
wire     [31:0] n49674;
wire     [31:0] n49675;
wire     [31:0] n49676;
wire     [31:0] n49677;
wire     [31:0] n49678;
wire     [31:0] n49679;
wire     [31:0] n49680;
wire     [31:0] n49681;
wire     [31:0] n49682;
wire     [31:0] n49683;
wire     [31:0] n49684;
wire     [31:0] n49685;
wire     [31:0] n49686;
wire     [31:0] n49687;
wire     [31:0] n49688;
wire     [31:0] n49689;
wire     [31:0] n49690;
wire     [31:0] n49691;
wire     [31:0] n49692;
wire     [31:0] n49693;
wire     [31:0] n49694;
wire     [31:0] n49695;
wire     [31:0] n49696;
wire     [31:0] n49697;
wire     [31:0] n49698;
wire     [31:0] n49699;
wire     [31:0] n49700;
wire     [31:0] n49701;
wire     [31:0] n49702;
wire     [31:0] n49703;
wire     [31:0] n49704;
wire     [31:0] n49705;
wire     [31:0] n49706;
wire     [31:0] n49707;
wire     [31:0] n49708;
wire     [31:0] n49709;
wire     [31:0] n49710;
wire     [31:0] n49711;
wire     [31:0] n49712;
wire     [31:0] n49713;
wire     [31:0] n49714;
wire     [31:0] n49715;
wire     [31:0] n49716;
wire     [31:0] n49717;
wire     [31:0] n49718;
wire     [31:0] n49719;
wire     [31:0] n49720;
wire     [31:0] n49721;
wire     [31:0] n49722;
wire     [31:0] n49723;
wire     [31:0] n49724;
wire     [31:0] n49725;
wire     [31:0] n49726;
wire     [31:0] n49727;
wire     [31:0] n49728;
wire     [31:0] n49729;
wire     [31:0] n49730;
wire     [31:0] n49731;
wire     [31:0] n49732;
wire     [31:0] n49733;
wire     [31:0] n49734;
wire     [31:0] n49735;
wire     [31:0] n49736;
wire     [31:0] n49737;
wire     [31:0] n49738;
wire     [31:0] n49739;
wire     [31:0] n49740;
wire     [31:0] n49741;
wire     [31:0] n49742;
wire     [31:0] n49743;
wire     [31:0] n49744;
wire     [31:0] n49745;
wire     [31:0] n49746;
wire     [31:0] n49747;
wire     [31:0] n49748;
wire     [31:0] n49749;
wire     [31:0] n49750;
wire     [31:0] n49751;
wire     [31:0] n49752;
wire     [31:0] n49753;
wire     [31:0] n49754;
wire     [31:0] n49755;
wire     [31:0] n49756;
wire     [31:0] n49757;
wire     [31:0] n49758;
wire     [31:0] n49759;
wire     [31:0] n49760;
wire     [31:0] n49761;
wire     [31:0] n49762;
wire     [31:0] n49763;
wire     [31:0] n49764;
wire     [31:0] n49765;
wire     [31:0] n49766;
wire     [31:0] n49767;
wire     [31:0] n49768;
wire     [31:0] n49769;
wire     [31:0] n49770;
wire     [31:0] n49771;
wire     [31:0] n49772;
wire     [31:0] n49773;
wire     [31:0] n49774;
wire     [31:0] n49775;
wire     [31:0] n49776;
wire     [31:0] n49777;
wire     [31:0] n49778;
wire     [31:0] n49779;
wire     [31:0] n49780;
wire     [31:0] n49781;
wire     [31:0] n49782;
wire     [31:0] n49783;
wire     [31:0] n49784;
wire     [31:0] n49785;
wire     [31:0] n49786;
wire     [31:0] n49787;
wire     [31:0] n49788;
wire     [31:0] n49789;
wire     [31:0] n49790;
wire     [31:0] n49791;
wire     [31:0] n49792;
wire     [31:0] n49793;
wire     [31:0] n49794;
wire     [31:0] n49795;
wire     [31:0] n49796;
wire     [31:0] n49797;
wire     [31:0] n49798;
wire     [31:0] n49799;
wire     [31:0] n49800;
wire     [31:0] n49801;
wire     [31:0] n49802;
wire     [31:0] n49803;
wire     [31:0] n49804;
wire     [31:0] n49805;
wire     [31:0] n49806;
wire     [31:0] n49807;
wire     [31:0] n49808;
wire     [31:0] n49809;
wire     [31:0] n49810;
wire     [31:0] n49811;
wire     [31:0] n49812;
wire     [31:0] n49813;
wire     [31:0] n49814;
wire     [31:0] n49815;
wire     [31:0] n49816;
wire     [31:0] n49817;
wire     [31:0] n49818;
wire     [31:0] n49819;
wire     [31:0] n49820;
wire     [31:0] n49821;
wire     [31:0] n49822;
wire     [31:0] n49823;
wire     [31:0] n49824;
wire     [31:0] n49825;
wire     [31:0] n49826;
wire     [31:0] n49827;
wire     [31:0] n49828;
wire     [31:0] n49829;
wire     [31:0] n49830;
wire     [31:0] n49831;
wire     [31:0] n49832;
wire     [31:0] n49833;
wire     [31:0] n49834;
wire     [31:0] n49835;
wire     [31:0] n49836;
wire     [31:0] n49837;
wire     [31:0] n49838;
wire     [31:0] n49839;
wire     [31:0] n49840;
wire     [31:0] n49841;
wire     [31:0] n49842;
wire     [31:0] n49843;
wire     [31:0] n49844;
wire     [31:0] n49845;
wire     [31:0] n49846;
wire     [31:0] n49847;
wire     [31:0] n49848;
wire     [31:0] n49849;
wire     [31:0] n49850;
wire     [31:0] n49851;
wire     [31:0] n49852;
wire     [31:0] n49853;
wire     [31:0] n49854;
wire     [31:0] n49855;
wire     [31:0] n49856;
wire     [31:0] n49857;
wire     [31:0] n49858;
wire     [31:0] n49859;
wire     [31:0] n49860;
wire     [31:0] n49861;
wire     [31:0] n49862;
wire     [31:0] n49863;
wire     [31:0] n49864;
wire     [31:0] n49865;
wire     [31:0] n49866;
wire     [31:0] n49867;
wire     [31:0] n49868;
wire     [31:0] n49869;
wire     [31:0] n49870;
wire     [31:0] n49871;
wire     [31:0] n49872;
wire     [31:0] n49873;
wire     [31:0] n49874;
wire     [31:0] n49875;
wire     [31:0] n49876;
wire     [31:0] n49877;
wire     [31:0] n49878;
wire     [31:0] n49879;
wire     [31:0] n49880;
wire     [31:0] n49881;
wire     [31:0] n49882;
wire     [31:0] n49883;
wire     [31:0] n49884;
wire     [31:0] n49885;
wire     [31:0] n49886;
wire     [31:0] n49887;
wire     [31:0] n49888;
wire     [31:0] n49889;
wire     [31:0] n49890;
wire     [31:0] n49891;
wire     [31:0] n49892;
wire     [31:0] n49893;
wire     [31:0] n49894;
wire     [31:0] n49895;
wire     [31:0] n49896;
wire     [31:0] n49897;
wire     [31:0] n49898;
wire     [31:0] n49899;
wire     [31:0] n49900;
wire     [31:0] n49901;
wire     [31:0] n49902;
wire     [31:0] n49903;
wire     [31:0] n49904;
wire     [31:0] n49905;
wire     [31:0] n49906;
wire     [31:0] n49907;
wire     [31:0] n49908;
wire     [31:0] n49909;
wire     [31:0] n49910;
wire     [31:0] n49911;
wire     [31:0] n49912;
wire     [31:0] n49913;
wire     [31:0] n49914;
wire     [31:0] n49915;
wire     [31:0] n49916;
wire     [31:0] n49917;
wire     [31:0] n49918;
wire     [31:0] n49919;
wire     [31:0] n49920;
wire     [31:0] n49921;
wire     [31:0] n49922;
wire     [31:0] n49923;
wire     [31:0] n49924;
wire     [31:0] n49925;
wire     [31:0] n49926;
wire     [31:0] n49927;
wire     [31:0] n49928;
wire     [31:0] n49929;
wire     [31:0] n49930;
wire     [31:0] n49931;
wire     [31:0] n49932;
wire     [31:0] n49933;
wire     [31:0] n49934;
wire     [31:0] n49935;
wire     [31:0] n49936;
wire     [31:0] n49937;
wire     [31:0] n49938;
wire     [31:0] n49939;
wire     [31:0] n49940;
wire     [31:0] n49941;
wire     [31:0] n49942;
wire     [31:0] n49943;
wire     [31:0] n49944;
wire     [31:0] n49945;
wire     [31:0] n49946;
wire     [31:0] n49947;
wire     [31:0] n49948;
wire     [31:0] n49949;
wire     [31:0] n49950;
wire     [31:0] n49951;
wire     [31:0] n49952;
wire     [31:0] n49953;
wire     [31:0] n49954;
wire     [31:0] n49955;
wire     [31:0] n49956;
wire     [31:0] n49957;
wire     [31:0] n49958;
wire     [31:0] n49959;
wire     [31:0] n49960;
wire     [31:0] n49961;
wire     [31:0] n49962;
wire     [31:0] n49963;
wire     [31:0] n49964;
wire     [31:0] n49965;
wire     [31:0] n49966;
wire     [31:0] n49967;
wire     [31:0] n49968;
wire     [31:0] n49969;
wire     [31:0] n49970;
wire     [31:0] n49971;
wire     [31:0] n49972;
wire     [31:0] n49973;
wire     [31:0] n49974;
wire     [31:0] n49975;
wire     [31:0] n49976;
wire     [31:0] n49977;
wire     [31:0] n49978;
wire     [31:0] n49979;
wire     [31:0] n49980;
wire     [31:0] n49981;
wire     [31:0] n49982;
wire     [31:0] n49983;
wire     [31:0] n49984;
wire     [31:0] n49985;
wire     [31:0] n49986;
wire     [31:0] n49987;
wire     [31:0] n49988;
wire     [31:0] n49989;
wire     [31:0] n49990;
wire     [31:0] n49991;
wire     [31:0] n49992;
wire     [31:0] n49993;
wire     [31:0] n49994;
wire     [31:0] n49995;
wire     [31:0] n49996;
wire     [31:0] n49997;
wire     [31:0] n49998;
wire     [31:0] n49999;
wire     [31:0] n50000;
wire     [31:0] n50001;
wire     [31:0] n50002;
wire     [31:0] n50003;
wire     [31:0] n50004;
wire     [31:0] n50005;
wire     [31:0] n50006;
wire     [31:0] n50007;
wire     [31:0] n50008;
wire     [31:0] n50009;
wire     [31:0] n50010;
wire     [31:0] n50011;
wire     [31:0] n50012;
wire     [31:0] n50013;
wire     [31:0] n50014;
wire     [31:0] n50015;
wire     [31:0] n50016;
wire     [31:0] n50017;
wire     [31:0] n50018;
wire     [31:0] n50019;
wire     [31:0] n50020;
wire     [31:0] n50021;
wire     [31:0] n50022;
wire     [31:0] n50023;
wire     [31:0] n50024;
wire     [31:0] n50025;
wire     [31:0] n50026;
wire     [31:0] n50027;
wire     [31:0] n50028;
wire     [31:0] n50029;
wire     [31:0] n50030;
wire     [31:0] n50031;
wire     [31:0] n50032;
wire     [31:0] n50033;
wire     [31:0] n50034;
wire     [31:0] n50035;
wire     [31:0] n50036;
wire     [31:0] n50037;
wire     [31:0] n50038;
wire     [31:0] n50039;
wire     [31:0] n50040;
wire     [31:0] n50041;
wire     [31:0] n50042;
wire     [31:0] n50043;
wire     [31:0] n50044;
wire     [31:0] n50045;
wire     [31:0] n50046;
wire     [31:0] n50047;
wire     [31:0] n50048;
wire     [31:0] n50049;
wire     [31:0] n50050;
wire     [31:0] n50051;
wire     [31:0] n50052;
wire     [31:0] n50053;
wire     [31:0] n50054;
wire     [31:0] n50055;
wire     [31:0] n50056;
wire     [31:0] n50057;
wire     [31:0] n50058;
wire     [31:0] n50059;
wire     [31:0] n50060;
wire     [31:0] n50061;
wire     [31:0] n50062;
wire     [31:0] n50063;
wire     [31:0] n50064;
wire     [31:0] n50065;
wire     [31:0] n50066;
wire     [31:0] n50067;
wire     [31:0] n50068;
wire     [31:0] n50069;
wire     [31:0] n50070;
wire     [31:0] n50071;
wire     [31:0] n50072;
wire     [31:0] n50073;
wire     [31:0] n50074;
wire     [31:0] n50075;
wire     [31:0] n50076;
wire     [31:0] n50077;
wire     [31:0] n50078;
wire     [31:0] n50079;
wire     [31:0] n50080;
wire     [31:0] n50081;
wire     [31:0] n50082;
wire     [31:0] n50083;
wire     [31:0] n50084;
wire     [31:0] n50085;
wire     [31:0] n50086;
wire     [31:0] n50087;
wire     [31:0] n50088;
wire     [31:0] n50089;
wire     [31:0] n50090;
wire     [31:0] n50091;
wire     [31:0] n50092;
wire     [31:0] n50093;
wire     [31:0] n50094;
wire     [31:0] n50095;
wire     [31:0] n50096;
wire     [31:0] n50097;
wire     [31:0] n50098;
wire     [31:0] n50099;
wire     [31:0] n50100;
wire     [31:0] n50101;
wire     [31:0] n50102;
wire     [31:0] n50103;
wire     [31:0] n50104;
wire     [31:0] n50105;
wire     [31:0] n50106;
wire     [31:0] n50107;
wire     [31:0] n50108;
wire     [31:0] n50109;
wire     [31:0] n50110;
wire     [31:0] n50111;
wire     [31:0] n50112;
wire     [31:0] n50113;
wire     [31:0] n50114;
wire     [31:0] n50115;
wire     [31:0] n50116;
wire     [31:0] n50117;
wire     [31:0] n50118;
wire     [31:0] n50119;
wire     [31:0] n50120;
wire     [31:0] n50121;
wire     [31:0] n50122;
wire     [31:0] n50123;
wire     [31:0] n50124;
wire     [31:0] n50125;
wire     [31:0] n50126;
wire     [31:0] n50127;
wire     [31:0] n50128;
wire     [31:0] n50129;
wire     [31:0] n50130;
wire     [31:0] n50131;
wire     [31:0] n50132;
wire     [31:0] n50133;
wire     [31:0] n50134;
wire     [31:0] n50135;
wire     [31:0] n50136;
wire     [31:0] n50137;
wire     [31:0] n50138;
wire     [31:0] n50139;
wire     [31:0] n50140;
wire     [31:0] n50141;
wire     [31:0] n50142;
wire     [31:0] n50143;
wire     [31:0] n50144;
wire     [31:0] n50145;
wire     [31:0] n50146;
wire     [31:0] n50147;
wire     [31:0] n50148;
wire     [31:0] n50149;
wire     [31:0] n50150;
wire     [31:0] n50151;
wire     [31:0] n50152;
wire     [31:0] n50153;
wire     [31:0] n50154;
wire     [31:0] n50155;
wire     [31:0] n50156;
wire     [31:0] n50157;
wire     [31:0] n50158;
wire     [31:0] n50159;
wire     [31:0] n50160;
wire     [31:0] n50161;
wire     [31:0] n50162;
wire     [31:0] n50163;
wire     [31:0] n50164;
wire     [31:0] n50165;
wire     [31:0] n50166;
wire     [31:0] n50167;
wire     [31:0] n50168;
wire     [31:0] n50169;
wire     [31:0] n50170;
wire     [31:0] n50171;
wire     [31:0] n50172;
wire     [31:0] n50173;
wire     [31:0] n50174;
wire     [31:0] n50175;
wire     [31:0] n50176;
wire     [31:0] n50177;
wire     [31:0] n50178;
wire     [31:0] n50179;
wire     [31:0] n50180;
wire     [31:0] n50181;
wire     [31:0] n50182;
wire     [31:0] n50183;
wire     [31:0] n50184;
wire     [31:0] n50185;
wire     [31:0] n50186;
wire     [31:0] n50187;
wire     [31:0] n50188;
wire     [31:0] n50189;
wire     [31:0] n50190;
wire     [31:0] n50191;
wire     [31:0] n50192;
wire     [31:0] n50193;
wire     [31:0] n50194;
wire     [31:0] n50195;
wire     [31:0] n50196;
wire     [31:0] n50197;
wire     [31:0] n50198;
wire     [31:0] n50199;
wire     [31:0] n50200;
wire     [31:0] n50201;
wire     [31:0] n50202;
wire     [31:0] n50203;
wire     [31:0] n50204;
wire     [31:0] n50205;
wire     [31:0] n50206;
wire     [31:0] n50207;
wire     [31:0] n50208;
wire     [31:0] n50209;
wire     [31:0] n50210;
wire     [31:0] n50211;
wire     [31:0] n50212;
wire     [31:0] n50213;
wire     [31:0] n50214;
wire     [31:0] n50215;
wire     [31:0] n50216;
wire     [31:0] n50217;
wire     [31:0] n50218;
wire     [31:0] n50219;
wire     [31:0] n50220;
wire     [31:0] n50221;
wire     [31:0] n50222;
wire     [31:0] n50223;
wire     [31:0] n50224;
wire     [31:0] n50225;
wire     [31:0] n50226;
wire     [31:0] n50227;
wire     [31:0] n50228;
wire     [31:0] n50229;
wire     [31:0] n50230;
wire     [31:0] n50231;
wire     [31:0] n50232;
wire     [31:0] n50233;
wire     [31:0] n50234;
wire     [31:0] n50235;
wire     [31:0] n50236;
wire     [31:0] n50237;
wire     [31:0] n50238;
wire     [31:0] n50239;
wire     [31:0] n50240;
wire     [31:0] n50241;
wire     [31:0] n50242;
wire     [31:0] n50243;
wire     [31:0] n50244;
wire     [31:0] n50245;
wire     [31:0] n50246;
wire     [31:0] n50247;
wire     [31:0] n50248;
wire     [31:0] n50249;
wire     [31:0] n50250;
wire     [31:0] n50251;
wire     [31:0] n50252;
wire     [31:0] n50253;
wire     [31:0] n50254;
wire     [31:0] n50255;
wire     [31:0] n50256;
wire     [31:0] n50257;
wire     [31:0] n50258;
wire     [31:0] n50259;
wire     [31:0] n50260;
wire     [31:0] n50261;
wire     [31:0] n50262;
wire     [31:0] n50263;
wire     [31:0] n50264;
wire     [31:0] n50265;
wire     [31:0] n50266;
wire     [31:0] n50267;
wire     [31:0] n50268;
wire     [31:0] n50269;
wire     [31:0] n50270;
wire     [31:0] n50271;
wire     [31:0] n50272;
wire     [31:0] n50273;
wire     [31:0] n50274;
wire     [31:0] n50275;
wire     [31:0] n50276;
wire     [31:0] n50277;
wire     [31:0] n50278;
wire     [31:0] n50279;
wire     [31:0] n50280;
wire     [31:0] n50281;
wire     [31:0] n50282;
wire     [31:0] n50283;
wire     [31:0] n50284;
wire     [31:0] n50285;
wire     [31:0] n50286;
wire     [31:0] n50287;
wire     [31:0] n50288;
wire     [31:0] n50289;
wire     [31:0] n50290;
wire     [31:0] n50291;
wire     [31:0] n50292;
wire     [31:0] n50293;
wire     [31:0] n50294;
wire     [31:0] n50295;
wire     [31:0] n50296;
wire     [31:0] n50297;
wire     [31:0] n50298;
wire     [31:0] n50299;
wire     [31:0] n50300;
wire     [31:0] n50301;
wire     [31:0] n50302;
wire     [31:0] n50303;
wire     [31:0] n50304;
wire     [31:0] n50305;
wire     [31:0] n50306;
wire     [31:0] n50307;
wire     [31:0] n50308;
wire     [31:0] n50309;
wire     [31:0] n50310;
wire     [31:0] n50311;
wire     [31:0] n50312;
wire     [31:0] n50313;
wire     [31:0] n50314;
wire     [31:0] n50315;
wire     [31:0] n50316;
wire     [31:0] n50317;
wire     [31:0] n50318;
wire     [31:0] n50319;
wire     [31:0] n50320;
wire     [31:0] n50321;
wire     [31:0] n50322;
wire     [31:0] n50323;
wire     [31:0] n50324;
wire     [31:0] n50325;
wire     [31:0] n50326;
wire     [31:0] n50327;
wire     [31:0] n50328;
wire     [31:0] n50329;
wire     [31:0] n50330;
wire     [31:0] n50331;
wire     [31:0] n50332;
wire     [31:0] n50333;
wire     [31:0] n50334;
wire     [31:0] n50335;
wire     [31:0] n50336;
wire     [31:0] n50337;
wire     [31:0] n50338;
wire     [31:0] n50339;
wire     [31:0] n50340;
wire     [31:0] n50341;
wire     [31:0] n50342;
wire     [31:0] n50343;
wire     [31:0] n50344;
wire     [31:0] n50345;
wire     [31:0] n50346;
wire     [31:0] n50347;
wire     [31:0] n50348;
wire     [31:0] n50349;
wire     [31:0] n50350;
wire     [31:0] n50351;
wire     [31:0] n50352;
wire     [31:0] n50353;
wire     [31:0] n50354;
wire     [31:0] n50355;
wire     [31:0] n50356;
wire     [31:0] n50357;
wire     [31:0] n50358;
wire     [31:0] n50359;
wire     [31:0] n50360;
wire     [31:0] n50361;
wire     [31:0] n50362;
wire     [31:0] n50363;
wire     [31:0] n50364;
wire     [31:0] n50365;
wire     [31:0] n50366;
wire     [31:0] n50367;
wire     [31:0] n50368;
wire     [31:0] n50369;
wire     [31:0] n50370;
wire     [31:0] n50371;
wire     [31:0] n50372;
wire     [31:0] n50373;
wire     [31:0] n50374;
wire     [31:0] n50375;
wire     [31:0] n50376;
wire     [31:0] n50377;
wire     [31:0] n50378;
wire     [31:0] n50379;
wire     [31:0] n50380;
wire     [31:0] n50381;
wire     [31:0] n50382;
wire     [31:0] n50383;
wire     [31:0] n50384;
wire     [31:0] n50385;
wire     [31:0] n50386;
wire     [31:0] n50387;
wire     [31:0] n50388;
wire     [31:0] n50389;
wire     [31:0] n50390;
wire     [31:0] n50391;
wire     [31:0] n50392;
wire     [31:0] n50393;
wire     [31:0] n50394;
wire     [31:0] n50395;
wire     [31:0] n50396;
wire     [31:0] n50397;
wire     [31:0] n50398;
wire     [31:0] n50399;
wire     [31:0] n50400;
wire     [31:0] n50401;
wire     [31:0] n50402;
wire     [31:0] n50403;
wire     [31:0] n50404;
wire     [31:0] n50405;
wire     [31:0] n50406;
wire     [31:0] n50407;
wire     [31:0] n50408;
wire     [31:0] n50409;
wire     [31:0] n50410;
wire     [31:0] n50411;
wire     [31:0] n50412;
wire     [31:0] n50413;
wire     [31:0] n50414;
wire     [31:0] n50415;
wire     [31:0] n50416;
wire     [31:0] n50417;
wire     [31:0] n50418;
wire     [31:0] n50419;
wire     [31:0] n50420;
wire     [31:0] n50421;
wire     [31:0] n50422;
wire     [31:0] n50423;
wire     [31:0] n50424;
wire     [31:0] n50425;
wire     [31:0] n50426;
wire     [31:0] n50427;
wire     [31:0] n50428;
wire     [31:0] n50429;
wire     [31:0] n50430;
wire     [31:0] n50431;
wire     [31:0] n50432;
wire     [31:0] n50433;
wire     [31:0] n50434;
wire     [31:0] n50435;
wire     [31:0] n50436;
wire     [31:0] n50437;
wire     [31:0] n50438;
wire     [31:0] n50439;
wire     [31:0] n50440;
wire     [31:0] n50441;
wire     [31:0] n50442;
wire     [31:0] n50443;
wire     [31:0] n50444;
wire     [31:0] n50445;
wire     [31:0] n50446;
wire     [31:0] n50447;
wire     [31:0] n50448;
wire     [31:0] n50449;
wire     [31:0] n50450;
wire     [31:0] n50451;
wire     [31:0] n50452;
wire     [31:0] n50453;
wire     [31:0] n50454;
wire     [31:0] n50455;
wire     [31:0] n50456;
wire     [31:0] n50457;
wire     [31:0] n50458;
wire     [31:0] n50459;
wire     [31:0] n50460;
wire     [31:0] n50461;
wire     [31:0] n50462;
wire     [31:0] n50463;
wire     [31:0] n50464;
wire     [31:0] n50465;
wire     [31:0] n50466;
wire     [31:0] n50467;
wire     [31:0] n50468;
wire     [31:0] n50469;
wire     [31:0] n50470;
wire     [31:0] n50471;
wire     [31:0] n50472;
wire     [31:0] n50473;
wire     [31:0] n50474;
wire     [31:0] n50475;
wire     [31:0] n50476;
wire     [31:0] n50477;
wire     [31:0] n50478;
wire     [31:0] n50479;
wire     [31:0] n50480;
wire     [31:0] n50481;
wire     [31:0] n50482;
wire     [31:0] n50483;
wire     [31:0] n50484;
wire     [31:0] n50485;
wire     [31:0] n50486;
wire     [31:0] n50487;
wire     [31:0] n50488;
wire     [31:0] n50489;
wire     [31:0] n50490;
wire     [31:0] n50491;
wire     [31:0] n50492;
wire     [31:0] n50493;
wire     [31:0] n50494;
wire     [31:0] n50495;
wire     [31:0] n50496;
wire     [31:0] n50497;
wire     [31:0] n50498;
wire     [31:0] n50499;
wire     [31:0] n50500;
wire     [31:0] n50501;
wire     [31:0] n50502;
wire     [31:0] n50503;
wire     [31:0] n50504;
wire     [31:0] n50505;
wire     [31:0] n50506;
wire     [31:0] n50507;
wire     [31:0] n50508;
wire     [31:0] n50509;
wire     [31:0] n50510;
wire     [31:0] n50511;
wire     [31:0] n50512;
wire     [31:0] n50513;
wire     [31:0] n50514;
wire     [31:0] n50515;
wire     [31:0] n50516;
wire     [31:0] n50517;
wire     [31:0] n50518;
wire     [31:0] n50519;
wire     [31:0] n50520;
wire     [31:0] n50521;
wire     [31:0] n50522;
wire     [31:0] n50523;
wire     [31:0] n50524;
wire     [31:0] n50525;
wire     [31:0] n50526;
wire     [31:0] n50527;
wire     [31:0] n50528;
wire     [31:0] n50529;
wire     [31:0] n50530;
wire     [31:0] n50531;
wire     [31:0] n50532;
wire     [31:0] n50533;
wire     [31:0] n50534;
wire     [31:0] n50535;
wire     [31:0] n50536;
wire     [31:0] n50537;
wire     [31:0] n50538;
wire     [31:0] n50539;
wire     [31:0] n50540;
wire     [31:0] n50541;
wire     [31:0] n50542;
wire     [31:0] n50543;
wire     [31:0] n50544;
wire     [31:0] n50545;
wire     [31:0] n50546;
wire     [31:0] n50547;
wire     [31:0] n50548;
wire     [31:0] n50549;
wire     [31:0] n50550;
wire     [31:0] n50551;
wire     [31:0] n50552;
wire     [31:0] n50553;
wire     [31:0] n50554;
wire     [31:0] n50555;
wire     [31:0] n50556;
wire     [31:0] n50557;
wire     [31:0] n50558;
wire     [31:0] n50559;
wire     [31:0] n50560;
wire     [31:0] n50561;
wire     [31:0] n50562;
wire     [31:0] n50563;
wire     [31:0] n50564;
wire     [31:0] n50565;
wire     [31:0] n50566;
wire     [31:0] n50567;
wire     [31:0] n50568;
wire     [31:0] n50569;
wire     [31:0] n50570;
wire     [31:0] n50571;
wire     [31:0] n50572;
wire     [31:0] n50573;
wire     [31:0] n50574;
wire     [31:0] n50575;
wire     [31:0] n50576;
wire     [31:0] n50577;
wire     [31:0] n50578;
wire     [31:0] n50579;
wire     [31:0] n50580;
wire     [31:0] n50581;
wire     [31:0] n50582;
wire     [31:0] n50583;
wire     [31:0] n50584;
wire     [31:0] n50585;
wire     [31:0] n50586;
wire     [31:0] n50587;
wire     [31:0] n50588;
wire     [31:0] n50589;
wire     [31:0] n50590;
wire     [31:0] n50591;
wire     [31:0] n50592;
wire     [31:0] n50593;
wire     [31:0] n50594;
wire     [31:0] n50595;
wire     [31:0] n50596;
wire     [31:0] n50597;
wire     [31:0] n50598;
wire     [31:0] n50599;
wire     [31:0] n50600;
wire     [31:0] n50601;
wire     [31:0] n50602;
wire     [31:0] n50603;
wire     [31:0] n50604;
wire     [31:0] n50605;
wire     [31:0] n50606;
wire     [31:0] n50607;
wire     [31:0] n50608;
wire     [31:0] n50609;
wire     [31:0] n50610;
wire     [31:0] n50611;
wire     [31:0] n50612;
wire     [31:0] n50613;
wire     [31:0] n50614;
wire     [31:0] n50615;
wire     [31:0] n50616;
wire     [31:0] n50617;
wire     [31:0] n50618;
wire     [31:0] n50619;
wire     [31:0] n50620;
wire     [31:0] n50621;
wire     [31:0] n50622;
wire     [31:0] n50623;
wire     [31:0] n50624;
wire     [31:0] n50625;
wire     [31:0] n50626;
wire     [31:0] n50627;
wire     [31:0] n50628;
wire     [31:0] n50629;
wire     [31:0] n50630;
wire     [31:0] n50631;
wire     [31:0] n50632;
wire     [31:0] n50633;
wire     [31:0] n50634;
wire     [31:0] n50635;
wire     [31:0] n50636;
wire     [31:0] n50637;
wire     [31:0] n50638;
wire     [31:0] n50639;
wire     [31:0] n50640;
wire     [31:0] n50641;
wire     [31:0] n50642;
wire     [31:0] n50643;
wire     [31:0] n50644;
wire     [31:0] n50645;
wire     [31:0] n50646;
wire     [31:0] n50647;
wire     [31:0] n50648;
wire     [31:0] n50649;
wire     [31:0] n50650;
wire     [31:0] n50651;
wire     [31:0] n50652;
wire     [31:0] n50653;
wire     [31:0] n50654;
wire     [31:0] n50655;
wire     [31:0] n50656;
wire     [31:0] n50657;
wire     [31:0] n50658;
wire     [31:0] n50659;
wire     [31:0] n50660;
wire     [31:0] n50661;
wire     [31:0] n50662;
wire     [31:0] n50663;
wire     [31:0] n50664;
wire     [31:0] n50665;
wire     [31:0] n50666;
wire     [31:0] n50667;
wire     [31:0] n50668;
wire     [31:0] n50669;
wire     [31:0] n50670;
wire     [31:0] n50671;
wire     [31:0] n50672;
wire     [31:0] n50673;
wire     [31:0] n50674;
wire     [31:0] n50675;
wire     [31:0] n50676;
wire     [31:0] n50677;
wire     [31:0] n50678;
wire     [31:0] n50679;
wire     [31:0] n50680;
wire     [31:0] n50681;
wire     [31:0] n50682;
wire     [31:0] n50683;
wire     [31:0] n50684;
wire     [31:0] n50685;
wire     [31:0] n50686;
wire     [31:0] n50687;
wire     [31:0] n50688;
wire     [31:0] n50689;
wire     [31:0] n50690;
wire     [31:0] n50691;
wire     [31:0] n50692;
wire     [31:0] n50693;
wire     [31:0] n50694;
wire     [31:0] n50695;
wire     [31:0] n50696;
wire     [31:0] n50697;
wire     [31:0] n50698;
wire     [31:0] n50699;
wire     [31:0] n50700;
wire     [31:0] n50701;
wire     [31:0] n50702;
wire     [31:0] n50703;
wire     [31:0] n50704;
wire     [31:0] n50705;
wire     [31:0] n50706;
wire     [31:0] n50707;
wire     [31:0] n50708;
wire     [31:0] n50709;
wire     [31:0] n50710;
wire     [31:0] n50711;
wire     [31:0] n50712;
wire     [31:0] n50713;
wire     [31:0] n50714;
wire     [31:0] n50715;
wire     [31:0] n50716;
wire     [31:0] n50717;
wire     [31:0] n50718;
wire     [31:0] n50719;
wire     [31:0] n50720;
wire     [31:0] n50721;
wire     [31:0] n50722;
wire     [31:0] n50723;
wire     [31:0] n50724;
wire     [31:0] n50725;
wire     [31:0] n50726;
wire     [31:0] n50727;
wire     [31:0] n50728;
wire     [31:0] n50729;
wire     [31:0] n50730;
wire     [31:0] n50731;
wire     [31:0] n50732;
wire     [31:0] n50733;
wire     [31:0] n50734;
wire     [31:0] n50735;
wire     [31:0] n50736;
wire     [31:0] n50737;
wire     [31:0] n50738;
wire     [31:0] n50739;
wire     [31:0] n50740;
wire     [31:0] n50741;
wire     [31:0] n50742;
wire     [31:0] n50743;
wire     [31:0] n50744;
wire     [31:0] n50745;
wire     [31:0] n50746;
wire     [31:0] n50747;
wire     [31:0] n50748;
wire     [31:0] n50749;
wire     [31:0] n50750;
wire     [31:0] n50751;
wire     [31:0] n50752;
wire     [31:0] n50753;
wire     [31:0] n50754;
wire     [31:0] n50755;
wire     [31:0] n50756;
wire     [31:0] n50757;
wire     [31:0] n50758;
wire     [31:0] n50759;
wire     [31:0] n50760;
wire     [31:0] n50761;
wire     [31:0] n50762;
wire     [31:0] n50763;
wire     [31:0] n50764;
wire     [31:0] n50765;
wire     [31:0] n50766;
wire     [31:0] n50767;
wire     [31:0] n50768;
wire     [31:0] n50769;
wire     [31:0] n50770;
wire     [31:0] n50771;
wire     [31:0] n50772;
wire     [31:0] n50773;
wire     [31:0] n50774;
wire     [31:0] n50775;
wire     [31:0] n50776;
wire     [31:0] n50777;
wire     [31:0] n50778;
wire     [31:0] n50779;
wire     [31:0] n50780;
wire     [31:0] n50781;
wire     [31:0] n50782;
wire     [31:0] n50783;
wire     [31:0] n50784;
wire     [31:0] n50785;
wire     [31:0] n50786;
wire     [31:0] n50787;
wire     [31:0] n50788;
wire     [31:0] n50789;
wire     [31:0] n50790;
wire     [31:0] n50791;
wire     [31:0] n50792;
wire     [31:0] n50793;
wire     [31:0] n50794;
wire     [31:0] n50795;
wire     [31:0] n50796;
wire     [31:0] n50797;
wire     [31:0] n50798;
wire     [31:0] n50799;
wire     [31:0] n50800;
wire     [31:0] n50801;
wire     [31:0] n50802;
wire     [31:0] n50803;
wire     [31:0] n50804;
wire     [31:0] n50805;
wire     [31:0] n50806;
wire     [31:0] n50807;
wire     [31:0] n50808;
wire     [31:0] n50809;
wire     [31:0] n50810;
wire     [31:0] n50811;
wire     [31:0] n50812;
wire     [31:0] n50813;
wire     [31:0] n50814;
wire     [31:0] n50815;
wire     [31:0] n50816;
wire     [31:0] n50817;
wire     [31:0] n50818;
wire     [31:0] n50819;
wire     [31:0] n50820;
wire     [31:0] n50821;
wire     [31:0] n50822;
wire     [31:0] n50823;
wire     [31:0] n50824;
wire     [31:0] n50825;
wire     [31:0] n50826;
wire     [31:0] n50827;
wire     [31:0] n50828;
wire     [31:0] n50829;
wire     [31:0] n50830;
wire     [31:0] n50831;
wire     [31:0] n50832;
wire     [31:0] n50833;
wire     [31:0] n50834;
wire     [31:0] n50835;
wire     [31:0] n50836;
wire     [31:0] n50837;
wire     [31:0] n50838;
wire     [31:0] n50839;
wire     [31:0] n50840;
wire     [31:0] n50841;
wire     [31:0] n50842;
wire     [31:0] n50843;
wire     [31:0] n50844;
wire     [31:0] n50845;
wire     [31:0] n50846;
wire     [31:0] n50847;
wire     [31:0] n50848;
wire     [31:0] n50849;
wire     [31:0] n50850;
wire     [31:0] n50851;
wire     [31:0] n50852;
wire     [31:0] n50853;
wire     [31:0] n50854;
wire     [31:0] n50855;
wire     [31:0] n50856;
wire     [31:0] n50857;
wire     [31:0] n50858;
wire     [31:0] n50859;
wire     [31:0] n50860;
wire     [31:0] n50861;
wire     [31:0] n50862;
wire     [31:0] n50863;
wire     [31:0] n50864;
wire     [31:0] n50865;
wire     [31:0] n50866;
wire     [31:0] n50867;
wire     [31:0] n50868;
wire     [31:0] n50869;
wire     [31:0] n50870;
wire     [31:0] n50871;
wire     [31:0] n50872;
wire     [31:0] n50873;
wire     [31:0] n50874;
wire     [31:0] n50875;
wire     [31:0] n50876;
wire     [31:0] n50877;
wire     [31:0] n50878;
wire     [31:0] n50879;
wire     [31:0] n50880;
wire     [31:0] n50881;
wire     [31:0] n50882;
wire     [31:0] n50883;
wire     [31:0] n50884;
wire     [31:0] n50885;
wire     [31:0] n50886;
wire     [31:0] n50887;
wire     [31:0] n50888;
wire     [31:0] n50889;
wire     [31:0] n50890;
wire     [31:0] n50891;
wire     [31:0] n50892;
wire     [31:0] n50893;
wire     [31:0] n50894;
wire     [31:0] n50895;
wire     [31:0] n50896;
wire     [31:0] n50897;
wire     [31:0] n50898;
wire     [31:0] n50899;
wire     [31:0] n50900;
wire     [31:0] n50901;
wire     [31:0] n50902;
wire     [31:0] n50903;
wire     [31:0] n50904;
wire     [31:0] n50905;
wire     [31:0] n50906;
wire     [31:0] n50907;
wire     [31:0] n50908;
wire     [31:0] n50909;
wire     [31:0] n50910;
wire     [31:0] n50911;
wire     [31:0] n50912;
wire     [31:0] n50913;
wire     [31:0] n50914;
wire     [31:0] n50915;
wire     [31:0] n50916;
wire     [31:0] n50917;
wire     [31:0] n50918;
wire     [31:0] n50919;
wire     [31:0] n50920;
wire     [31:0] n50921;
wire     [31:0] n50922;
wire     [31:0] n50923;
wire     [31:0] n50924;
wire     [31:0] n50925;
wire     [31:0] n50926;
wire     [31:0] n50927;
wire     [31:0] n50928;
wire     [31:0] n50929;
wire     [31:0] n50930;
wire     [31:0] n50931;
wire     [31:0] n50932;
wire     [31:0] n50933;
wire     [31:0] n50934;
wire     [31:0] n50935;
wire     [31:0] n50936;
wire     [31:0] n50937;
wire     [31:0] n50938;
wire     [31:0] n50939;
wire     [31:0] n50940;
wire     [31:0] n50941;
wire     [31:0] n50942;
wire     [31:0] n50943;
wire     [31:0] n50944;
wire     [31:0] n50945;
wire     [31:0] n50946;
wire     [31:0] n50947;
wire     [31:0] n50948;
wire     [31:0] n50949;
wire     [31:0] n50950;
wire     [31:0] n50951;
wire     [31:0] n50952;
wire     [31:0] n50953;
wire     [31:0] n50954;
wire     [31:0] n50955;
wire     [31:0] n50956;
wire     [31:0] n50957;
wire     [31:0] n50958;
wire     [31:0] n50959;
wire     [31:0] n50960;
wire     [31:0] n50961;
wire     [31:0] n50962;
wire     [31:0] n50963;
wire     [31:0] n50964;
wire     [31:0] n50965;
wire     [31:0] n50966;
wire     [31:0] n50967;
wire     [31:0] n50968;
wire     [31:0] n50969;
wire     [31:0] n50970;
wire     [31:0] n50971;
wire     [31:0] n50972;
wire     [31:0] n50973;
wire     [31:0] n50974;
wire     [31:0] n50975;
wire     [31:0] n50976;
wire     [31:0] n50977;
wire     [31:0] n50978;
wire     [31:0] n50979;
wire     [31:0] n50980;
wire     [31:0] n50981;
wire     [31:0] n50982;
wire     [31:0] n50983;
wire     [31:0] n50984;
wire     [31:0] n50985;
wire     [31:0] n50986;
wire     [31:0] n50987;
wire     [31:0] n50988;
wire     [31:0] n50989;
wire     [31:0] n50990;
wire     [31:0] n50991;
wire     [31:0] n50992;
wire     [31:0] n50993;
wire     [31:0] n50994;
wire     [31:0] n50995;
wire     [31:0] n50996;
wire     [31:0] n50997;
wire     [31:0] n50998;
wire     [31:0] n50999;
wire     [31:0] n51000;
wire     [31:0] n51001;
wire     [31:0] n51002;
wire     [31:0] n51003;
wire     [31:0] n51004;
wire     [31:0] n51005;
wire     [31:0] n51006;
wire     [31:0] n51007;
wire     [31:0] n51008;
wire     [31:0] n51009;
wire     [31:0] n51010;
wire     [31:0] n51011;
wire     [31:0] n51012;
wire     [31:0] n51013;
wire     [31:0] n51014;
wire     [31:0] n51015;
wire     [31:0] n51016;
wire     [31:0] n51017;
wire     [31:0] n51018;
wire     [31:0] n51019;
wire     [31:0] n51020;
wire     [31:0] n51021;
wire     [31:0] n51022;
wire     [31:0] n51023;
wire     [31:0] n51024;
wire     [31:0] n51025;
wire     [31:0] n51026;
wire     [31:0] n51027;
wire     [31:0] n51028;
wire     [31:0] n51029;
wire     [31:0] n51030;
wire     [31:0] n51031;
wire     [31:0] n51032;
wire     [31:0] n51033;
wire     [31:0] n51034;
wire     [31:0] n51035;
wire     [31:0] n51036;
wire     [31:0] n51037;
wire     [31:0] n51038;
wire     [31:0] n51039;
wire     [31:0] n51040;
wire     [31:0] n51041;
wire     [31:0] n51042;
wire     [31:0] n51043;
wire     [31:0] n51044;
wire     [31:0] n51045;
wire     [31:0] n51046;
wire     [31:0] n51047;
wire     [31:0] n51048;
wire     [31:0] n51049;
wire     [31:0] n51050;
wire     [31:0] n51051;
wire     [31:0] n51052;
wire     [31:0] n51053;
wire     [31:0] n51054;
wire     [31:0] n51055;
wire     [31:0] n51056;
wire     [31:0] n51057;
wire     [31:0] n51058;
wire     [31:0] n51059;
wire     [31:0] n51060;
wire     [31:0] n51061;
wire     [31:0] n51062;
wire     [31:0] n51063;
wire     [31:0] n51064;
wire     [31:0] n51065;
wire     [31:0] n51066;
wire     [31:0] n51067;
wire     [31:0] n51068;
wire     [31:0] n51069;
wire     [31:0] n51070;
wire     [31:0] n51071;
wire     [31:0] n51072;
wire     [31:0] n51073;
wire     [31:0] n51074;
wire     [31:0] n51075;
wire     [31:0] n51076;
wire     [31:0] n51077;
wire     [31:0] n51078;
wire     [31:0] n51079;
wire     [31:0] n51080;
wire     [31:0] n51081;
wire     [31:0] n51082;
wire     [31:0] n51083;
wire     [31:0] n51084;
wire     [31:0] n51085;
wire     [31:0] n51086;
wire     [31:0] n51087;
wire     [31:0] n51088;
wire     [31:0] n51089;
wire     [31:0] n51090;
wire     [31:0] n51091;
wire     [31:0] n51092;
wire     [31:0] n51093;
wire     [31:0] n51094;
wire     [31:0] n51095;
wire     [31:0] n51096;
wire     [31:0] n51097;
wire     [31:0] n51098;
wire     [31:0] n51099;
wire     [31:0] n51100;
wire     [31:0] n51101;
wire     [31:0] n51102;
wire     [31:0] n51103;
wire     [31:0] n51104;
wire     [31:0] n51105;
wire     [31:0] n51106;
wire     [31:0] n51107;
wire     [31:0] n51108;
wire     [31:0] n51109;
wire     [31:0] n51110;
wire     [31:0] n51111;
wire     [31:0] n51112;
wire     [31:0] n51113;
wire     [31:0] n51114;
wire     [31:0] n51115;
wire     [31:0] n51116;
wire     [31:0] n51117;
wire     [31:0] n51118;
wire     [31:0] n51119;
wire     [31:0] n51120;
wire     [31:0] n51121;
wire     [31:0] n51122;
wire     [31:0] n51123;
wire     [31:0] n51124;
wire     [31:0] n51125;
wire     [31:0] n51126;
wire     [31:0] n51127;
wire     [31:0] n51128;
wire     [31:0] n51129;
wire     [31:0] n51130;
wire     [31:0] n51131;
wire     [31:0] n51132;
wire     [31:0] n51133;
wire     [31:0] n51134;
wire     [31:0] n51135;
wire     [31:0] n51136;
wire     [31:0] n51137;
wire     [31:0] n51138;
wire     [31:0] n51139;
wire     [31:0] n51140;
wire     [31:0] n51141;
wire     [31:0] n51142;
wire     [31:0] n51143;
wire     [31:0] n51144;
wire     [31:0] n51145;
wire     [31:0] n51146;
wire     [31:0] n51147;
wire     [31:0] n51148;
wire     [31:0] n51149;
wire     [31:0] n51150;
wire     [31:0] n51151;
wire     [31:0] n51152;
wire     [31:0] n51153;
wire     [31:0] n51154;
wire     [31:0] n51155;
wire     [31:0] n51156;
wire     [31:0] n51157;
wire     [31:0] n51158;
wire     [31:0] n51159;
wire     [31:0] n51160;
wire     [31:0] n51161;
wire     [31:0] n51162;
wire     [31:0] n51163;
wire     [31:0] n51164;
wire     [31:0] n51165;
wire     [31:0] n51166;
wire     [31:0] n51167;
wire     [31:0] n51168;
wire     [31:0] n51169;
wire     [31:0] n51170;
wire     [31:0] n51171;
wire     [31:0] n51172;
wire     [31:0] n51173;
wire     [31:0] n51174;
wire     [31:0] n51175;
wire     [31:0] n51176;
wire     [31:0] n51177;
wire     [31:0] n51178;
wire     [31:0] n51179;
wire     [31:0] n51180;
wire     [31:0] n51181;
wire     [31:0] n51182;
wire     [31:0] n51183;
wire     [31:0] n51184;
wire     [31:0] n51185;
wire     [31:0] n51186;
wire     [31:0] n51187;
wire     [31:0] n51188;
wire     [31:0] n51189;
wire     [31:0] n51190;
wire     [31:0] n51191;
wire     [31:0] n51192;
wire     [31:0] n51193;
wire     [31:0] n51194;
wire     [31:0] n51195;
wire     [31:0] n51196;
wire     [31:0] n51197;
wire     [31:0] n51198;
wire     [31:0] n51199;
wire     [31:0] n51200;
wire     [31:0] n51201;
wire     [31:0] n51202;
wire     [31:0] n51203;
wire     [31:0] n51204;
wire     [31:0] n51205;
wire     [31:0] n51206;
wire     [31:0] n51207;
wire     [31:0] n51208;
wire     [31:0] n51209;
wire     [31:0] n51210;
wire     [31:0] n51211;
wire     [31:0] n51212;
wire     [31:0] n51213;
wire     [31:0] n51214;
wire     [31:0] n51215;
wire     [31:0] n51216;
wire     [31:0] n51217;
wire     [31:0] n51218;
wire     [31:0] n51219;
wire     [31:0] n51220;
wire     [31:0] n51221;
wire     [31:0] n51222;
reg     [31:0] mem;
wire clk;
wire rst;
wire step;
assign n0 = pc[31:2] ;
assign n1 =  {2'd0 , n0}  ;
assign imem_raddr_ila = n1  ;
assign n2 = imem_rdata_ila  ;
//assign n2 =  (  mem [ n1 ] )  ;
assign n3 = n2[9:5] ;
assign n4 =  ( n3 ) == ( 5'd0 )  ;
assign n5 = n2[31:29] ;
assign n6 =  ( n5 ) == ( 3'd6 )  ;
assign n7 = n2[28:26] ;
assign n8 =  ( n7 ) == ( 3'd0 )  ;
assign n9 = n2[25:20] ;
assign n10 =  ( n9 ) == ( 6'd5 )  ;
assign n11 = n2[4:0] ;
assign n12 =  ( n11 ) == ( 5'd31 )  ;
assign n13 =  ( n11 ) == ( 5'd30 )  ;
assign n14 =  ( n11 ) == ( 5'd29 )  ;
assign n15 =  ( n11 ) == ( 5'd28 )  ;
assign n16 =  ( n11 ) == ( 5'd27 )  ;
assign n17 =  ( n11 ) == ( 5'd26 )  ;
assign n18 =  ( n11 ) == ( 5'd25 )  ;
assign n19 =  ( n11 ) == ( 5'd24 )  ;
assign n20 =  ( n11 ) == ( 5'd23 )  ;
assign n21 =  ( n11 ) == ( 5'd22 )  ;
assign n22 =  ( n11 ) == ( 5'd21 )  ;
assign n23 =  ( n11 ) == ( 5'd20 )  ;
assign n24 =  ( n11 ) == ( 5'd19 )  ;
assign n25 =  ( n11 ) == ( 5'd18 )  ;
assign n26 =  ( n11 ) == ( 5'd17 )  ;
assign n27 =  ( n11 ) == ( 5'd16 )  ;
assign n28 =  ( n11 ) == ( 5'd15 )  ;
assign n29 =  ( n11 ) == ( 5'd14 )  ;
assign n30 =  ( n11 ) == ( 5'd13 )  ;
assign n31 =  ( n11 ) == ( 5'd12 )  ;
assign n32 =  ( n11 ) == ( 5'd11 )  ;
assign n33 =  ( n11 ) == ( 5'd10 )  ;
assign n34 =  ( n11 ) == ( 5'd9 )  ;
assign n35 =  ( n11 ) == ( 5'd8 )  ;
assign n36 =  ( n11 ) == ( 5'd7 )  ;
assign n37 =  ( n11 ) == ( 5'd6 )  ;
assign n38 =  ( n11 ) == ( 5'd5 )  ;
assign n39 =  ( n11 ) == ( 5'd4 )  ;
assign n40 =  ( n11 ) == ( 5'd3 )  ;
assign n41 =  ( n11 ) == ( 5'd2 )  ;
assign n42 =  ( n11 ) == ( 5'd1 )  ;
assign n43 =  ( n11 ) == ( 5'd0 )  ;
assign n44 =  ( n43 ) ? ( SREG_0 ) : ( SREG_0 ) ;
assign n45 =  ( n42 ) ? ( SREG_1 ) : ( n44 ) ;
assign n46 =  ( n41 ) ? ( SREG_2 ) : ( n45 ) ;
assign n47 =  ( n40 ) ? ( SREG_3 ) : ( n46 ) ;
assign n48 =  ( n39 ) ? ( SREG_4 ) : ( n47 ) ;
assign n49 =  ( n38 ) ? ( SREG_5 ) : ( n48 ) ;
assign n50 =  ( n37 ) ? ( SREG_6 ) : ( n49 ) ;
assign n51 =  ( n36 ) ? ( SREG_7 ) : ( n50 ) ;
assign n52 =  ( n35 ) ? ( SREG_8 ) : ( n51 ) ;
assign n53 =  ( n34 ) ? ( SREG_9 ) : ( n52 ) ;
assign n54 =  ( n33 ) ? ( SREG_10 ) : ( n53 ) ;
assign n55 =  ( n32 ) ? ( SREG_11 ) : ( n54 ) ;
assign n56 =  ( n31 ) ? ( SREG_12 ) : ( n55 ) ;
assign n57 =  ( n30 ) ? ( SREG_13 ) : ( n56 ) ;
assign n58 =  ( n29 ) ? ( SREG_14 ) : ( n57 ) ;
assign n59 =  ( n28 ) ? ( SREG_15 ) : ( n58 ) ;
assign n60 =  ( n27 ) ? ( SREG_16 ) : ( n59 ) ;
assign n61 =  ( n26 ) ? ( SREG_17 ) : ( n60 ) ;
assign n62 =  ( n25 ) ? ( SREG_18 ) : ( n61 ) ;
assign n63 =  ( n24 ) ? ( SREG_19 ) : ( n62 ) ;
assign n64 =  ( n23 ) ? ( SREG_20 ) : ( n63 ) ;
assign n65 =  ( n22 ) ? ( SREG_21 ) : ( n64 ) ;
assign n66 =  ( n21 ) ? ( SREG_22 ) : ( n65 ) ;
assign n67 =  ( n20 ) ? ( SREG_23 ) : ( n66 ) ;
assign n68 =  ( n19 ) ? ( SREG_24 ) : ( n67 ) ;
assign n69 =  ( n18 ) ? ( SREG_25 ) : ( n68 ) ;
assign n70 =  ( n17 ) ? ( SREG_26 ) : ( n69 ) ;
assign n71 =  ( n16 ) ? ( SREG_27 ) : ( n70 ) ;
assign n72 =  ( n15 ) ? ( SREG_28 ) : ( n71 ) ;
assign n73 =  ( n14 ) ? ( SREG_29 ) : ( n72 ) ;
assign n74 =  ( n13 ) ? ( SREG_30 ) : ( n73 ) ;
assign n75 =  ( n12 ) ? ( SREG_31 ) : ( n74 ) ;
assign n76 = n2[19:15] ;
assign n77 =  ( n76 ) == ( 5'd31 )  ;
assign n78 =  ( n76 ) == ( 5'd30 )  ;
assign n79 =  ( n76 ) == ( 5'd29 )  ;
assign n80 =  ( n76 ) == ( 5'd28 )  ;
assign n81 =  ( n76 ) == ( 5'd27 )  ;
assign n82 =  ( n76 ) == ( 5'd26 )  ;
assign n83 =  ( n76 ) == ( 5'd25 )  ;
assign n84 =  ( n76 ) == ( 5'd24 )  ;
assign n85 =  ( n76 ) == ( 5'd23 )  ;
assign n86 =  ( n76 ) == ( 5'd22 )  ;
assign n87 =  ( n76 ) == ( 5'd21 )  ;
assign n88 =  ( n76 ) == ( 5'd20 )  ;
assign n89 =  ( n76 ) == ( 5'd19 )  ;
assign n90 =  ( n76 ) == ( 5'd18 )  ;
assign n91 =  ( n76 ) == ( 5'd17 )  ;
assign n92 =  ( n76 ) == ( 5'd16 )  ;
assign n93 =  ( n76 ) == ( 5'd15 )  ;
assign n94 =  ( n76 ) == ( 5'd14 )  ;
assign n95 =  ( n76 ) == ( 5'd13 )  ;
assign n96 =  ( n76 ) == ( 5'd12 )  ;
assign n97 =  ( n76 ) == ( 5'd11 )  ;
assign n98 =  ( n76 ) == ( 5'd10 )  ;
assign n99 =  ( n76 ) == ( 5'd9 )  ;
assign n100 =  ( n76 ) == ( 5'd8 )  ;
assign n101 =  ( n76 ) == ( 5'd7 )  ;
assign n102 =  ( n76 ) == ( 5'd6 )  ;
assign n103 =  ( n76 ) == ( 5'd5 )  ;
assign n104 =  ( n76 ) == ( 5'd4 )  ;
assign n105 =  ( n76 ) == ( 5'd3 )  ;
assign n106 =  ( n76 ) == ( 5'd2 )  ;
assign n107 =  ( n76 ) == ( 5'd1 )  ;
assign n108 =  ( n76 ) == ( 5'd0 )  ;
assign n109 =  ( n108 ) ? ( SREG_0 ) : ( SREG_0 ) ;
assign n110 =  ( n107 ) ? ( SREG_1 ) : ( n109 ) ;
assign n111 =  ( n106 ) ? ( SREG_2 ) : ( n110 ) ;
assign n112 =  ( n105 ) ? ( SREG_3 ) : ( n111 ) ;
assign n113 =  ( n104 ) ? ( SREG_4 ) : ( n112 ) ;
assign n114 =  ( n103 ) ? ( SREG_5 ) : ( n113 ) ;
assign n115 =  ( n102 ) ? ( SREG_6 ) : ( n114 ) ;
assign n116 =  ( n101 ) ? ( SREG_7 ) : ( n115 ) ;
assign n117 =  ( n100 ) ? ( SREG_8 ) : ( n116 ) ;
assign n118 =  ( n99 ) ? ( SREG_9 ) : ( n117 ) ;
assign n119 =  ( n98 ) ? ( SREG_10 ) : ( n118 ) ;
assign n120 =  ( n97 ) ? ( SREG_11 ) : ( n119 ) ;
assign n121 =  ( n96 ) ? ( SREG_12 ) : ( n120 ) ;
assign n122 =  ( n95 ) ? ( SREG_13 ) : ( n121 ) ;
assign n123 =  ( n94 ) ? ( SREG_14 ) : ( n122 ) ;
assign n124 =  ( n93 ) ? ( SREG_15 ) : ( n123 ) ;
assign n125 =  ( n92 ) ? ( SREG_16 ) : ( n124 ) ;
assign n126 =  ( n91 ) ? ( SREG_17 ) : ( n125 ) ;
assign n127 =  ( n90 ) ? ( SREG_18 ) : ( n126 ) ;
assign n128 =  ( n89 ) ? ( SREG_19 ) : ( n127 ) ;
assign n129 =  ( n88 ) ? ( SREG_20 ) : ( n128 ) ;
assign n130 =  ( n87 ) ? ( SREG_21 ) : ( n129 ) ;
assign n131 =  ( n86 ) ? ( SREG_22 ) : ( n130 ) ;
assign n132 =  ( n85 ) ? ( SREG_23 ) : ( n131 ) ;
assign n133 =  ( n84 ) ? ( SREG_24 ) : ( n132 ) ;
assign n134 =  ( n83 ) ? ( SREG_25 ) : ( n133 ) ;
assign n135 =  ( n82 ) ? ( SREG_26 ) : ( n134 ) ;
assign n136 =  ( n81 ) ? ( SREG_27 ) : ( n135 ) ;
assign n137 =  ( n80 ) ? ( SREG_28 ) : ( n136 ) ;
assign n138 =  ( n79 ) ? ( SREG_29 ) : ( n137 ) ;
assign n139 =  ( n78 ) ? ( SREG_30 ) : ( n138 ) ;
assign n140 =  ( n77 ) ? ( SREG_31 ) : ( n139 ) ;
assign n141 =  ( n75 ) + ( n140 )  ;
assign n142 =  ( n9 ) == ( 6'd6 )  ;
assign n143 =  ( n75 ) - ( n140 )  ;
assign n144 =  ( n9 ) == ( 6'd1 )  ;
assign n145 =  ( n75 ) & ( n140 )  ;
assign n146 =  ( n9 ) == ( 6'd0 )  ;
assign n147 =  ( n75 ) | ( n140 )  ;
assign n148 =  ( n9 ) == ( 6'd31 )  ;
assign n149 =  ( ( n75 ) * ( n140 ))  ;
assign n150 =  ( n148 ) ? ( n149 ) : ( SREG_0 ) ;
assign n151 =  ( n146 ) ? ( n147 ) : ( n150 ) ;
assign n152 =  ( n144 ) ? ( n145 ) : ( n151 ) ;
assign n153 =  ( n142 ) ? ( n143 ) : ( n152 ) ;
assign n154 =  ( n10 ) ? ( n141 ) : ( n153 ) ;
assign n155 =  ( n8 ) ? ( n154 ) : ( SREG_0 ) ;
assign n156 = n2[31:31] ;
assign n157 =  ( n156 ) == ( 1'd0 )  ;
assign n158 = n2[30:29] ;
assign n159 =  ( n158 ) == ( 2'd0 )  ;
assign n160 = n2[28:24] ;
assign n161 =  {1'd0 , n160}  ;
assign n162 =  ( n161 ) == ( 6'd5 )  ;
assign n163 = n2[23:10] ;
assign n164 =  {18'd0 , n163}  ;
assign n165 =  ( n75 ) + ( n164 )  ;
assign n166 =  ( n161 ) == ( 6'd6 )  ;
assign n167 =  ( n75 ) - ( n164 )  ;
assign n168 =  ( n161 ) == ( 6'd1 )  ;
assign n169 =  ( n75 ) & ( n164 )  ;
assign n170 =  ( n161 ) == ( 6'd0 )  ;
assign n171 =  ( n75 ) | ( n164 )  ;
assign n172 =  ( n161 ) == ( 6'd31 )  ;
assign n173 =  ( n172 ) ? ( n149 ) : ( SREG_0 ) ;
assign n174 =  ( n170 ) ? ( n171 ) : ( n173 ) ;
assign n175 =  ( n168 ) ? ( n169 ) : ( n174 ) ;
assign n176 =  ( n166 ) ? ( n167 ) : ( n175 ) ;
assign n177 =  ( n162 ) ? ( n165 ) : ( n176 ) ;
assign n178 =  ( n158 ) == ( 2'd2 )  ;
assign n179 = n2[23:15] ;
assign n180 =  {23'd0 , n179}  ;
assign n181 =  ( n75 ) + ( n180 )  ;
assign n182 =  ( n75 ) - ( n180 )  ;
assign n183 =  ( n75 ) & ( n180 )  ;
assign n184 =  ( n75 ) | ( n180 )  ;
assign n185 =  ( n170 ) ? ( n184 ) : ( n173 ) ;
assign n186 =  ( n168 ) ? ( n183 ) : ( n185 ) ;
assign n187 =  ( n166 ) ? ( n182 ) : ( n186 ) ;
assign n188 =  ( n162 ) ? ( n181 ) : ( n187 ) ;
assign n189 =  ( n178 ) ? ( n188 ) : ( SREG_0 ) ;
assign n190 =  ( n159 ) ? ( n177 ) : ( n189 ) ;
assign n191 = n2[29:29] ;
assign n192 =  ( n191 ) == ( 1'd1 )  ;
assign n193 =  ( n192 ) ? ( SREG_0 ) : ( SREG_0 ) ;
assign n194 =  ( n157 ) ? ( n190 ) : ( n193 ) ;
assign n195 =  ( n6 ) ? ( n155 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( n195 ) : ( SREG_0 ) ;
assign n197 =  ( n3 ) == ( 5'd1 )  ;
assign n198 =  ( n148 ) ? ( n149 ) : ( SREG_1 ) ;
assign n199 =  ( n146 ) ? ( n147 ) : ( n198 ) ;
assign n200 =  ( n144 ) ? ( n145 ) : ( n199 ) ;
assign n201 =  ( n142 ) ? ( n143 ) : ( n200 ) ;
assign n202 =  ( n10 ) ? ( n141 ) : ( n201 ) ;
assign n203 =  ( n8 ) ? ( n202 ) : ( SREG_1 ) ;
assign n204 =  ( n172 ) ? ( n149 ) : ( SREG_1 ) ;
assign n205 =  ( n170 ) ? ( n171 ) : ( n204 ) ;
assign n206 =  ( n168 ) ? ( n169 ) : ( n205 ) ;
assign n207 =  ( n166 ) ? ( n167 ) : ( n206 ) ;
assign n208 =  ( n162 ) ? ( n165 ) : ( n207 ) ;
assign n209 =  ( n170 ) ? ( n184 ) : ( n204 ) ;
assign n210 =  ( n168 ) ? ( n183 ) : ( n209 ) ;
assign n211 =  ( n166 ) ? ( n182 ) : ( n210 ) ;
assign n212 =  ( n162 ) ? ( n181 ) : ( n211 ) ;
assign n213 =  ( n178 ) ? ( n212 ) : ( SREG_1 ) ;
assign n214 =  ( n159 ) ? ( n208 ) : ( n213 ) ;
assign n215 =  ( n192 ) ? ( SREG_1 ) : ( SREG_1 ) ;
assign n216 =  ( n157 ) ? ( n214 ) : ( n215 ) ;
assign n217 =  ( n6 ) ? ( n203 ) : ( n216 ) ;
assign n218 =  ( n197 ) ? ( n217 ) : ( SREG_1 ) ;
assign n219 =  ( n3 ) == ( 5'd10 )  ;
assign n220 =  ( n148 ) ? ( n149 ) : ( SREG_10 ) ;
assign n221 =  ( n146 ) ? ( n147 ) : ( n220 ) ;
assign n222 =  ( n144 ) ? ( n145 ) : ( n221 ) ;
assign n223 =  ( n142 ) ? ( n143 ) : ( n222 ) ;
assign n224 =  ( n10 ) ? ( n141 ) : ( n223 ) ;
assign n225 =  ( n8 ) ? ( n224 ) : ( SREG_10 ) ;
assign n226 =  ( n172 ) ? ( n149 ) : ( SREG_10 ) ;
assign n227 =  ( n170 ) ? ( n171 ) : ( n226 ) ;
assign n228 =  ( n168 ) ? ( n169 ) : ( n227 ) ;
assign n229 =  ( n166 ) ? ( n167 ) : ( n228 ) ;
assign n230 =  ( n162 ) ? ( n165 ) : ( n229 ) ;
assign n231 =  ( n170 ) ? ( n184 ) : ( n226 ) ;
assign n232 =  ( n168 ) ? ( n183 ) : ( n231 ) ;
assign n233 =  ( n166 ) ? ( n182 ) : ( n232 ) ;
assign n234 =  ( n162 ) ? ( n181 ) : ( n233 ) ;
assign n235 =  ( n178 ) ? ( n234 ) : ( SREG_10 ) ;
assign n236 =  ( n159 ) ? ( n230 ) : ( n235 ) ;
assign n237 =  ( n192 ) ? ( SREG_10 ) : ( SREG_10 ) ;
assign n238 =  ( n157 ) ? ( n236 ) : ( n237 ) ;
assign n239 =  ( n6 ) ? ( n225 ) : ( n238 ) ;
assign n240 =  ( n219 ) ? ( n239 ) : ( SREG_10 ) ;
assign n241 =  ( n3 ) == ( 5'd11 )  ;
assign n242 =  ( n148 ) ? ( n149 ) : ( SREG_11 ) ;
assign n243 =  ( n146 ) ? ( n147 ) : ( n242 ) ;
assign n244 =  ( n144 ) ? ( n145 ) : ( n243 ) ;
assign n245 =  ( n142 ) ? ( n143 ) : ( n244 ) ;
assign n246 =  ( n10 ) ? ( n141 ) : ( n245 ) ;
assign n247 =  ( n8 ) ? ( n246 ) : ( SREG_11 ) ;
assign n248 =  ( n172 ) ? ( n149 ) : ( SREG_11 ) ;
assign n249 =  ( n170 ) ? ( n171 ) : ( n248 ) ;
assign n250 =  ( n168 ) ? ( n169 ) : ( n249 ) ;
assign n251 =  ( n166 ) ? ( n167 ) : ( n250 ) ;
assign n252 =  ( n162 ) ? ( n165 ) : ( n251 ) ;
assign n253 =  ( n170 ) ? ( n184 ) : ( n248 ) ;
assign n254 =  ( n168 ) ? ( n183 ) : ( n253 ) ;
assign n255 =  ( n166 ) ? ( n182 ) : ( n254 ) ;
assign n256 =  ( n162 ) ? ( n181 ) : ( n255 ) ;
assign n257 =  ( n178 ) ? ( n256 ) : ( SREG_11 ) ;
assign n258 =  ( n159 ) ? ( n252 ) : ( n257 ) ;
assign n259 =  ( n192 ) ? ( SREG_11 ) : ( SREG_11 ) ;
assign n260 =  ( n157 ) ? ( n258 ) : ( n259 ) ;
assign n261 =  ( n6 ) ? ( n247 ) : ( n260 ) ;
assign n262 =  ( n241 ) ? ( n261 ) : ( SREG_11 ) ;
assign n263 =  ( n3 ) == ( 5'd12 )  ;
assign n264 =  ( n148 ) ? ( n149 ) : ( SREG_12 ) ;
assign n265 =  ( n146 ) ? ( n147 ) : ( n264 ) ;
assign n266 =  ( n144 ) ? ( n145 ) : ( n265 ) ;
assign n267 =  ( n142 ) ? ( n143 ) : ( n266 ) ;
assign n268 =  ( n10 ) ? ( n141 ) : ( n267 ) ;
assign n269 =  ( n8 ) ? ( n268 ) : ( SREG_12 ) ;
assign n270 =  ( n172 ) ? ( n149 ) : ( SREG_12 ) ;
assign n271 =  ( n170 ) ? ( n171 ) : ( n270 ) ;
assign n272 =  ( n168 ) ? ( n169 ) : ( n271 ) ;
assign n273 =  ( n166 ) ? ( n167 ) : ( n272 ) ;
assign n274 =  ( n162 ) ? ( n165 ) : ( n273 ) ;
assign n275 =  ( n170 ) ? ( n184 ) : ( n270 ) ;
assign n276 =  ( n168 ) ? ( n183 ) : ( n275 ) ;
assign n277 =  ( n166 ) ? ( n182 ) : ( n276 ) ;
assign n278 =  ( n162 ) ? ( n181 ) : ( n277 ) ;
assign n279 =  ( n178 ) ? ( n278 ) : ( SREG_12 ) ;
assign n280 =  ( n159 ) ? ( n274 ) : ( n279 ) ;
assign n281 =  ( n192 ) ? ( SREG_12 ) : ( SREG_12 ) ;
assign n282 =  ( n157 ) ? ( n280 ) : ( n281 ) ;
assign n283 =  ( n6 ) ? ( n269 ) : ( n282 ) ;
assign n284 =  ( n263 ) ? ( n283 ) : ( SREG_12 ) ;
assign n285 =  ( n3 ) == ( 5'd13 )  ;
assign n286 =  ( n148 ) ? ( n149 ) : ( SREG_13 ) ;
assign n287 =  ( n146 ) ? ( n147 ) : ( n286 ) ;
assign n288 =  ( n144 ) ? ( n145 ) : ( n287 ) ;
assign n289 =  ( n142 ) ? ( n143 ) : ( n288 ) ;
assign n290 =  ( n10 ) ? ( n141 ) : ( n289 ) ;
assign n291 =  ( n8 ) ? ( n290 ) : ( SREG_13 ) ;
assign n292 =  ( n172 ) ? ( n149 ) : ( SREG_13 ) ;
assign n293 =  ( n170 ) ? ( n171 ) : ( n292 ) ;
assign n294 =  ( n168 ) ? ( n169 ) : ( n293 ) ;
assign n295 =  ( n166 ) ? ( n167 ) : ( n294 ) ;
assign n296 =  ( n162 ) ? ( n165 ) : ( n295 ) ;
assign n297 =  ( n170 ) ? ( n184 ) : ( n292 ) ;
assign n298 =  ( n168 ) ? ( n183 ) : ( n297 ) ;
assign n299 =  ( n166 ) ? ( n182 ) : ( n298 ) ;
assign n300 =  ( n162 ) ? ( n181 ) : ( n299 ) ;
assign n301 =  ( n178 ) ? ( n300 ) : ( SREG_13 ) ;
assign n302 =  ( n159 ) ? ( n296 ) : ( n301 ) ;
assign n303 =  ( n192 ) ? ( SREG_13 ) : ( SREG_13 ) ;
assign n304 =  ( n157 ) ? ( n302 ) : ( n303 ) ;
assign n305 =  ( n6 ) ? ( n291 ) : ( n304 ) ;
assign n306 =  ( n285 ) ? ( n305 ) : ( SREG_13 ) ;
assign n307 =  ( n3 ) == ( 5'd14 )  ;
assign n308 =  ( n148 ) ? ( n149 ) : ( SREG_14 ) ;
assign n309 =  ( n146 ) ? ( n147 ) : ( n308 ) ;
assign n310 =  ( n144 ) ? ( n145 ) : ( n309 ) ;
assign n311 =  ( n142 ) ? ( n143 ) : ( n310 ) ;
assign n312 =  ( n10 ) ? ( n141 ) : ( n311 ) ;
assign n313 =  ( n8 ) ? ( n312 ) : ( SREG_14 ) ;
assign n314 =  ( n172 ) ? ( n149 ) : ( SREG_14 ) ;
assign n315 =  ( n170 ) ? ( n171 ) : ( n314 ) ;
assign n316 =  ( n168 ) ? ( n169 ) : ( n315 ) ;
assign n317 =  ( n166 ) ? ( n167 ) : ( n316 ) ;
assign n318 =  ( n162 ) ? ( n165 ) : ( n317 ) ;
assign n319 =  ( n170 ) ? ( n184 ) : ( n314 ) ;
assign n320 =  ( n168 ) ? ( n183 ) : ( n319 ) ;
assign n321 =  ( n166 ) ? ( n182 ) : ( n320 ) ;
assign n322 =  ( n162 ) ? ( n181 ) : ( n321 ) ;
assign n323 =  ( n178 ) ? ( n322 ) : ( SREG_14 ) ;
assign n324 =  ( n159 ) ? ( n318 ) : ( n323 ) ;
assign n325 =  ( n192 ) ? ( SREG_14 ) : ( SREG_14 ) ;
assign n326 =  ( n157 ) ? ( n324 ) : ( n325 ) ;
assign n327 =  ( n6 ) ? ( n313 ) : ( n326 ) ;
assign n328 =  ( n307 ) ? ( n327 ) : ( SREG_14 ) ;
assign n329 =  ( n3 ) == ( 5'd15 )  ;
assign n330 =  ( n148 ) ? ( n149 ) : ( SREG_15 ) ;
assign n331 =  ( n146 ) ? ( n147 ) : ( n330 ) ;
assign n332 =  ( n144 ) ? ( n145 ) : ( n331 ) ;
assign n333 =  ( n142 ) ? ( n143 ) : ( n332 ) ;
assign n334 =  ( n10 ) ? ( n141 ) : ( n333 ) ;
assign n335 =  ( n8 ) ? ( n334 ) : ( SREG_15 ) ;
assign n336 =  ( n172 ) ? ( n149 ) : ( SREG_15 ) ;
assign n337 =  ( n170 ) ? ( n171 ) : ( n336 ) ;
assign n338 =  ( n168 ) ? ( n169 ) : ( n337 ) ;
assign n339 =  ( n166 ) ? ( n167 ) : ( n338 ) ;
assign n340 =  ( n162 ) ? ( n165 ) : ( n339 ) ;
assign n341 =  ( n170 ) ? ( n184 ) : ( n336 ) ;
assign n342 =  ( n168 ) ? ( n183 ) : ( n341 ) ;
assign n343 =  ( n166 ) ? ( n182 ) : ( n342 ) ;
assign n344 =  ( n162 ) ? ( n181 ) : ( n343 ) ;
assign n345 =  ( n178 ) ? ( n344 ) : ( SREG_15 ) ;
assign n346 =  ( n159 ) ? ( n340 ) : ( n345 ) ;
assign n347 =  ( n192 ) ? ( SREG_15 ) : ( SREG_15 ) ;
assign n348 =  ( n157 ) ? ( n346 ) : ( n347 ) ;
assign n349 =  ( n6 ) ? ( n335 ) : ( n348 ) ;
assign n350 =  ( n329 ) ? ( n349 ) : ( SREG_15 ) ;
assign n351 =  ( n3 ) == ( 5'd16 )  ;
assign n352 =  ( n148 ) ? ( n149 ) : ( SREG_16 ) ;
assign n353 =  ( n146 ) ? ( n147 ) : ( n352 ) ;
assign n354 =  ( n144 ) ? ( n145 ) : ( n353 ) ;
assign n355 =  ( n142 ) ? ( n143 ) : ( n354 ) ;
assign n356 =  ( n10 ) ? ( n141 ) : ( n355 ) ;
assign n357 =  ( n8 ) ? ( n356 ) : ( SREG_16 ) ;
assign n358 =  ( n172 ) ? ( n149 ) : ( SREG_16 ) ;
assign n359 =  ( n170 ) ? ( n171 ) : ( n358 ) ;
assign n360 =  ( n168 ) ? ( n169 ) : ( n359 ) ;
assign n361 =  ( n166 ) ? ( n167 ) : ( n360 ) ;
assign n362 =  ( n162 ) ? ( n165 ) : ( n361 ) ;
assign n363 =  ( n170 ) ? ( n184 ) : ( n358 ) ;
assign n364 =  ( n168 ) ? ( n183 ) : ( n363 ) ;
assign n365 =  ( n166 ) ? ( n182 ) : ( n364 ) ;
assign n366 =  ( n162 ) ? ( n181 ) : ( n365 ) ;
assign n367 =  ( n178 ) ? ( n366 ) : ( SREG_16 ) ;
assign n368 =  ( n159 ) ? ( n362 ) : ( n367 ) ;
assign n369 =  ( n192 ) ? ( SREG_16 ) : ( SREG_16 ) ;
assign n370 =  ( n157 ) ? ( n368 ) : ( n369 ) ;
assign n371 =  ( n6 ) ? ( n357 ) : ( n370 ) ;
assign n372 =  ( n351 ) ? ( n371 ) : ( SREG_16 ) ;
assign n373 =  ( n3 ) == ( 5'd17 )  ;
assign n374 =  ( n148 ) ? ( n149 ) : ( SREG_17 ) ;
assign n375 =  ( n146 ) ? ( n147 ) : ( n374 ) ;
assign n376 =  ( n144 ) ? ( n145 ) : ( n375 ) ;
assign n377 =  ( n142 ) ? ( n143 ) : ( n376 ) ;
assign n378 =  ( n10 ) ? ( n141 ) : ( n377 ) ;
assign n379 =  ( n8 ) ? ( n378 ) : ( SREG_17 ) ;
assign n380 =  ( n172 ) ? ( n149 ) : ( SREG_17 ) ;
assign n381 =  ( n170 ) ? ( n171 ) : ( n380 ) ;
assign n382 =  ( n168 ) ? ( n169 ) : ( n381 ) ;
assign n383 =  ( n166 ) ? ( n167 ) : ( n382 ) ;
assign n384 =  ( n162 ) ? ( n165 ) : ( n383 ) ;
assign n385 =  ( n170 ) ? ( n184 ) : ( n380 ) ;
assign n386 =  ( n168 ) ? ( n183 ) : ( n385 ) ;
assign n387 =  ( n166 ) ? ( n182 ) : ( n386 ) ;
assign n388 =  ( n162 ) ? ( n181 ) : ( n387 ) ;
assign n389 =  ( n178 ) ? ( n388 ) : ( SREG_17 ) ;
assign n390 =  ( n159 ) ? ( n384 ) : ( n389 ) ;
assign n391 =  ( n192 ) ? ( SREG_17 ) : ( SREG_17 ) ;
assign n392 =  ( n157 ) ? ( n390 ) : ( n391 ) ;
assign n393 =  ( n6 ) ? ( n379 ) : ( n392 ) ;
assign n394 =  ( n373 ) ? ( n393 ) : ( SREG_17 ) ;
assign n395 =  ( n3 ) == ( 5'd18 )  ;
assign n396 =  ( n148 ) ? ( n149 ) : ( SREG_18 ) ;
assign n397 =  ( n146 ) ? ( n147 ) : ( n396 ) ;
assign n398 =  ( n144 ) ? ( n145 ) : ( n397 ) ;
assign n399 =  ( n142 ) ? ( n143 ) : ( n398 ) ;
assign n400 =  ( n10 ) ? ( n141 ) : ( n399 ) ;
assign n401 =  ( n8 ) ? ( n400 ) : ( SREG_18 ) ;
assign n402 =  ( n172 ) ? ( n149 ) : ( SREG_18 ) ;
assign n403 =  ( n170 ) ? ( n171 ) : ( n402 ) ;
assign n404 =  ( n168 ) ? ( n169 ) : ( n403 ) ;
assign n405 =  ( n166 ) ? ( n167 ) : ( n404 ) ;
assign n406 =  ( n162 ) ? ( n165 ) : ( n405 ) ;
assign n407 =  ( n170 ) ? ( n184 ) : ( n402 ) ;
assign n408 =  ( n168 ) ? ( n183 ) : ( n407 ) ;
assign n409 =  ( n166 ) ? ( n182 ) : ( n408 ) ;
assign n410 =  ( n162 ) ? ( n181 ) : ( n409 ) ;
assign n411 =  ( n178 ) ? ( n410 ) : ( SREG_18 ) ;
assign n412 =  ( n159 ) ? ( n406 ) : ( n411 ) ;
assign n413 =  ( n192 ) ? ( SREG_18 ) : ( SREG_18 ) ;
assign n414 =  ( n157 ) ? ( n412 ) : ( n413 ) ;
assign n415 =  ( n6 ) ? ( n401 ) : ( n414 ) ;
assign n416 =  ( n395 ) ? ( n415 ) : ( SREG_18 ) ;
assign n417 =  ( n3 ) == ( 5'd19 )  ;
assign n418 =  ( n148 ) ? ( n149 ) : ( SREG_19 ) ;
assign n419 =  ( n146 ) ? ( n147 ) : ( n418 ) ;
assign n420 =  ( n144 ) ? ( n145 ) : ( n419 ) ;
assign n421 =  ( n142 ) ? ( n143 ) : ( n420 ) ;
assign n422 =  ( n10 ) ? ( n141 ) : ( n421 ) ;
assign n423 =  ( n8 ) ? ( n422 ) : ( SREG_19 ) ;
assign n424 =  ( n172 ) ? ( n149 ) : ( SREG_19 ) ;
assign n425 =  ( n170 ) ? ( n171 ) : ( n424 ) ;
assign n426 =  ( n168 ) ? ( n169 ) : ( n425 ) ;
assign n427 =  ( n166 ) ? ( n167 ) : ( n426 ) ;
assign n428 =  ( n162 ) ? ( n165 ) : ( n427 ) ;
assign n429 =  ( n170 ) ? ( n184 ) : ( n424 ) ;
assign n430 =  ( n168 ) ? ( n183 ) : ( n429 ) ;
assign n431 =  ( n166 ) ? ( n182 ) : ( n430 ) ;
assign n432 =  ( n162 ) ? ( n181 ) : ( n431 ) ;
assign n433 =  ( n178 ) ? ( n432 ) : ( SREG_19 ) ;
assign n434 =  ( n159 ) ? ( n428 ) : ( n433 ) ;
assign n435 =  ( n192 ) ? ( SREG_19 ) : ( SREG_19 ) ;
assign n436 =  ( n157 ) ? ( n434 ) : ( n435 ) ;
assign n437 =  ( n6 ) ? ( n423 ) : ( n436 ) ;
assign n438 =  ( n417 ) ? ( n437 ) : ( SREG_19 ) ;
assign n439 =  ( n3 ) == ( 5'd2 )  ;
assign n440 =  ( n148 ) ? ( n149 ) : ( SREG_2 ) ;
assign n441 =  ( n146 ) ? ( n147 ) : ( n440 ) ;
assign n442 =  ( n144 ) ? ( n145 ) : ( n441 ) ;
assign n443 =  ( n142 ) ? ( n143 ) : ( n442 ) ;
assign n444 =  ( n10 ) ? ( n141 ) : ( n443 ) ;
assign n445 =  ( n8 ) ? ( n444 ) : ( SREG_2 ) ;
assign n446 =  ( n172 ) ? ( n149 ) : ( SREG_2 ) ;
assign n447 =  ( n170 ) ? ( n171 ) : ( n446 ) ;
assign n448 =  ( n168 ) ? ( n169 ) : ( n447 ) ;
assign n449 =  ( n166 ) ? ( n167 ) : ( n448 ) ;
assign n450 =  ( n162 ) ? ( n165 ) : ( n449 ) ;
assign n451 =  ( n170 ) ? ( n184 ) : ( n446 ) ;
assign n452 =  ( n168 ) ? ( n183 ) : ( n451 ) ;
assign n453 =  ( n166 ) ? ( n182 ) : ( n452 ) ;
assign n454 =  ( n162 ) ? ( n181 ) : ( n453 ) ;
assign n455 =  ( n178 ) ? ( n454 ) : ( SREG_2 ) ;
assign n456 =  ( n159 ) ? ( n450 ) : ( n455 ) ;
assign n457 =  ( n192 ) ? ( SREG_2 ) : ( SREG_2 ) ;
assign n458 =  ( n157 ) ? ( n456 ) : ( n457 ) ;
assign n459 =  ( n6 ) ? ( n445 ) : ( n458 ) ;
assign n460 =  ( n439 ) ? ( n459 ) : ( SREG_2 ) ;
assign n461 =  ( n3 ) == ( 5'd20 )  ;
assign n462 =  ( n148 ) ? ( n149 ) : ( SREG_20 ) ;
assign n463 =  ( n146 ) ? ( n147 ) : ( n462 ) ;
assign n464 =  ( n144 ) ? ( n145 ) : ( n463 ) ;
assign n465 =  ( n142 ) ? ( n143 ) : ( n464 ) ;
assign n466 =  ( n10 ) ? ( n141 ) : ( n465 ) ;
assign n467 =  ( n8 ) ? ( n466 ) : ( SREG_20 ) ;
assign n468 =  ( n172 ) ? ( n149 ) : ( SREG_20 ) ;
assign n469 =  ( n170 ) ? ( n171 ) : ( n468 ) ;
assign n470 =  ( n168 ) ? ( n169 ) : ( n469 ) ;
assign n471 =  ( n166 ) ? ( n167 ) : ( n470 ) ;
assign n472 =  ( n162 ) ? ( n165 ) : ( n471 ) ;
assign n473 =  ( n170 ) ? ( n184 ) : ( n468 ) ;
assign n474 =  ( n168 ) ? ( n183 ) : ( n473 ) ;
assign n475 =  ( n166 ) ? ( n182 ) : ( n474 ) ;
assign n476 =  ( n162 ) ? ( n181 ) : ( n475 ) ;
assign n477 =  ( n178 ) ? ( n476 ) : ( SREG_20 ) ;
assign n478 =  ( n159 ) ? ( n472 ) : ( n477 ) ;
assign n479 =  ( n192 ) ? ( SREG_20 ) : ( SREG_20 ) ;
assign n480 =  ( n157 ) ? ( n478 ) : ( n479 ) ;
assign n481 =  ( n6 ) ? ( n467 ) : ( n480 ) ;
assign n482 =  ( n461 ) ? ( n481 ) : ( SREG_20 ) ;
assign n483 =  ( n3 ) == ( 5'd21 )  ;
assign n484 =  ( n148 ) ? ( n149 ) : ( SREG_21 ) ;
assign n485 =  ( n146 ) ? ( n147 ) : ( n484 ) ;
assign n486 =  ( n144 ) ? ( n145 ) : ( n485 ) ;
assign n487 =  ( n142 ) ? ( n143 ) : ( n486 ) ;
assign n488 =  ( n10 ) ? ( n141 ) : ( n487 ) ;
assign n489 =  ( n8 ) ? ( n488 ) : ( SREG_21 ) ;
assign n490 =  ( n172 ) ? ( n149 ) : ( SREG_21 ) ;
assign n491 =  ( n170 ) ? ( n171 ) : ( n490 ) ;
assign n492 =  ( n168 ) ? ( n169 ) : ( n491 ) ;
assign n493 =  ( n166 ) ? ( n167 ) : ( n492 ) ;
assign n494 =  ( n162 ) ? ( n165 ) : ( n493 ) ;
assign n495 =  ( n170 ) ? ( n184 ) : ( n490 ) ;
assign n496 =  ( n168 ) ? ( n183 ) : ( n495 ) ;
assign n497 =  ( n166 ) ? ( n182 ) : ( n496 ) ;
assign n498 =  ( n162 ) ? ( n181 ) : ( n497 ) ;
assign n499 =  ( n178 ) ? ( n498 ) : ( SREG_21 ) ;
assign n500 =  ( n159 ) ? ( n494 ) : ( n499 ) ;
assign n501 =  ( n192 ) ? ( SREG_21 ) : ( SREG_21 ) ;
assign n502 =  ( n157 ) ? ( n500 ) : ( n501 ) ;
assign n503 =  ( n6 ) ? ( n489 ) : ( n502 ) ;
assign n504 =  ( n483 ) ? ( n503 ) : ( SREG_21 ) ;
assign n505 =  ( n3 ) == ( 5'd22 )  ;
assign n506 =  ( n148 ) ? ( n149 ) : ( SREG_22 ) ;
assign n507 =  ( n146 ) ? ( n147 ) : ( n506 ) ;
assign n508 =  ( n144 ) ? ( n145 ) : ( n507 ) ;
assign n509 =  ( n142 ) ? ( n143 ) : ( n508 ) ;
assign n510 =  ( n10 ) ? ( n141 ) : ( n509 ) ;
assign n511 =  ( n8 ) ? ( n510 ) : ( SREG_22 ) ;
assign n512 =  ( n172 ) ? ( n149 ) : ( SREG_22 ) ;
assign n513 =  ( n170 ) ? ( n171 ) : ( n512 ) ;
assign n514 =  ( n168 ) ? ( n169 ) : ( n513 ) ;
assign n515 =  ( n166 ) ? ( n167 ) : ( n514 ) ;
assign n516 =  ( n162 ) ? ( n165 ) : ( n515 ) ;
assign n517 =  ( n170 ) ? ( n184 ) : ( n512 ) ;
assign n518 =  ( n168 ) ? ( n183 ) : ( n517 ) ;
assign n519 =  ( n166 ) ? ( n182 ) : ( n518 ) ;
assign n520 =  ( n162 ) ? ( n181 ) : ( n519 ) ;
assign n521 =  ( n178 ) ? ( n520 ) : ( SREG_22 ) ;
assign n522 =  ( n159 ) ? ( n516 ) : ( n521 ) ;
assign n523 =  ( n192 ) ? ( SREG_22 ) : ( SREG_22 ) ;
assign n524 =  ( n157 ) ? ( n522 ) : ( n523 ) ;
assign n525 =  ( n6 ) ? ( n511 ) : ( n524 ) ;
assign n526 =  ( n505 ) ? ( n525 ) : ( SREG_22 ) ;
assign n527 =  ( n3 ) == ( 5'd23 )  ;
assign n528 =  ( n148 ) ? ( n149 ) : ( SREG_23 ) ;
assign n529 =  ( n146 ) ? ( n147 ) : ( n528 ) ;
assign n530 =  ( n144 ) ? ( n145 ) : ( n529 ) ;
assign n531 =  ( n142 ) ? ( n143 ) : ( n530 ) ;
assign n532 =  ( n10 ) ? ( n141 ) : ( n531 ) ;
assign n533 =  ( n8 ) ? ( n532 ) : ( SREG_23 ) ;
assign n534 =  ( n172 ) ? ( n149 ) : ( SREG_23 ) ;
assign n535 =  ( n170 ) ? ( n171 ) : ( n534 ) ;
assign n536 =  ( n168 ) ? ( n169 ) : ( n535 ) ;
assign n537 =  ( n166 ) ? ( n167 ) : ( n536 ) ;
assign n538 =  ( n162 ) ? ( n165 ) : ( n537 ) ;
assign n539 =  ( n170 ) ? ( n184 ) : ( n534 ) ;
assign n540 =  ( n168 ) ? ( n183 ) : ( n539 ) ;
assign n541 =  ( n166 ) ? ( n182 ) : ( n540 ) ;
assign n542 =  ( n162 ) ? ( n181 ) : ( n541 ) ;
assign n543 =  ( n178 ) ? ( n542 ) : ( SREG_23 ) ;
assign n544 =  ( n159 ) ? ( n538 ) : ( n543 ) ;
assign n545 =  ( n192 ) ? ( SREG_23 ) : ( SREG_23 ) ;
assign n546 =  ( n157 ) ? ( n544 ) : ( n545 ) ;
assign n547 =  ( n6 ) ? ( n533 ) : ( n546 ) ;
assign n548 =  ( n527 ) ? ( n547 ) : ( SREG_23 ) ;
assign n549 =  ( n3 ) == ( 5'd24 )  ;
assign n550 =  ( n148 ) ? ( n149 ) : ( SREG_24 ) ;
assign n551 =  ( n146 ) ? ( n147 ) : ( n550 ) ;
assign n552 =  ( n144 ) ? ( n145 ) : ( n551 ) ;
assign n553 =  ( n142 ) ? ( n143 ) : ( n552 ) ;
assign n554 =  ( n10 ) ? ( n141 ) : ( n553 ) ;
assign n555 =  ( n8 ) ? ( n554 ) : ( SREG_24 ) ;
assign n556 =  ( n172 ) ? ( n149 ) : ( SREG_24 ) ;
assign n557 =  ( n170 ) ? ( n171 ) : ( n556 ) ;
assign n558 =  ( n168 ) ? ( n169 ) : ( n557 ) ;
assign n559 =  ( n166 ) ? ( n167 ) : ( n558 ) ;
assign n560 =  ( n162 ) ? ( n165 ) : ( n559 ) ;
assign n561 =  ( n170 ) ? ( n184 ) : ( n556 ) ;
assign n562 =  ( n168 ) ? ( n183 ) : ( n561 ) ;
assign n563 =  ( n166 ) ? ( n182 ) : ( n562 ) ;
assign n564 =  ( n162 ) ? ( n181 ) : ( n563 ) ;
assign n565 =  ( n178 ) ? ( n564 ) : ( SREG_24 ) ;
assign n566 =  ( n159 ) ? ( n560 ) : ( n565 ) ;
assign n567 =  ( n192 ) ? ( SREG_24 ) : ( SREG_24 ) ;
assign n568 =  ( n157 ) ? ( n566 ) : ( n567 ) ;
assign n569 =  ( n6 ) ? ( n555 ) : ( n568 ) ;
assign n570 =  ( n549 ) ? ( n569 ) : ( SREG_24 ) ;
assign n571 =  ( n3 ) == ( 5'd25 )  ;
assign n572 =  ( n148 ) ? ( n149 ) : ( SREG_25 ) ;
assign n573 =  ( n146 ) ? ( n147 ) : ( n572 ) ;
assign n574 =  ( n144 ) ? ( n145 ) : ( n573 ) ;
assign n575 =  ( n142 ) ? ( n143 ) : ( n574 ) ;
assign n576 =  ( n10 ) ? ( n141 ) : ( n575 ) ;
assign n577 =  ( n8 ) ? ( n576 ) : ( SREG_25 ) ;
assign n578 =  ( n172 ) ? ( n149 ) : ( SREG_25 ) ;
assign n579 =  ( n170 ) ? ( n171 ) : ( n578 ) ;
assign n580 =  ( n168 ) ? ( n169 ) : ( n579 ) ;
assign n581 =  ( n166 ) ? ( n167 ) : ( n580 ) ;
assign n582 =  ( n162 ) ? ( n165 ) : ( n581 ) ;
assign n583 =  ( n170 ) ? ( n184 ) : ( n578 ) ;
assign n584 =  ( n168 ) ? ( n183 ) : ( n583 ) ;
assign n585 =  ( n166 ) ? ( n182 ) : ( n584 ) ;
assign n586 =  ( n162 ) ? ( n181 ) : ( n585 ) ;
assign n587 =  ( n178 ) ? ( n586 ) : ( SREG_25 ) ;
assign n588 =  ( n159 ) ? ( n582 ) : ( n587 ) ;
assign n589 =  ( n192 ) ? ( SREG_25 ) : ( SREG_25 ) ;
assign n590 =  ( n157 ) ? ( n588 ) : ( n589 ) ;
assign n591 =  ( n6 ) ? ( n577 ) : ( n590 ) ;
assign n592 =  ( n571 ) ? ( n591 ) : ( SREG_25 ) ;
assign n593 =  ( n3 ) == ( 5'd26 )  ;
assign n594 =  ( n148 ) ? ( n149 ) : ( SREG_26 ) ;
assign n595 =  ( n146 ) ? ( n147 ) : ( n594 ) ;
assign n596 =  ( n144 ) ? ( n145 ) : ( n595 ) ;
assign n597 =  ( n142 ) ? ( n143 ) : ( n596 ) ;
assign n598 =  ( n10 ) ? ( n141 ) : ( n597 ) ;
assign n599 =  ( n8 ) ? ( n598 ) : ( SREG_26 ) ;
assign n600 =  ( n172 ) ? ( n149 ) : ( SREG_26 ) ;
assign n601 =  ( n170 ) ? ( n171 ) : ( n600 ) ;
assign n602 =  ( n168 ) ? ( n169 ) : ( n601 ) ;
assign n603 =  ( n166 ) ? ( n167 ) : ( n602 ) ;
assign n604 =  ( n162 ) ? ( n165 ) : ( n603 ) ;
assign n605 =  ( n170 ) ? ( n184 ) : ( n600 ) ;
assign n606 =  ( n168 ) ? ( n183 ) : ( n605 ) ;
assign n607 =  ( n166 ) ? ( n182 ) : ( n606 ) ;
assign n608 =  ( n162 ) ? ( n181 ) : ( n607 ) ;
assign n609 =  ( n178 ) ? ( n608 ) : ( SREG_26 ) ;
assign n610 =  ( n159 ) ? ( n604 ) : ( n609 ) ;
assign n611 =  ( n192 ) ? ( SREG_26 ) : ( SREG_26 ) ;
assign n612 =  ( n157 ) ? ( n610 ) : ( n611 ) ;
assign n613 =  ( n6 ) ? ( n599 ) : ( n612 ) ;
assign n614 =  ( n593 ) ? ( n613 ) : ( SREG_26 ) ;
assign n615 =  ( n3 ) == ( 5'd27 )  ;
assign n616 =  ( n148 ) ? ( n149 ) : ( SREG_27 ) ;
assign n617 =  ( n146 ) ? ( n147 ) : ( n616 ) ;
assign n618 =  ( n144 ) ? ( n145 ) : ( n617 ) ;
assign n619 =  ( n142 ) ? ( n143 ) : ( n618 ) ;
assign n620 =  ( n10 ) ? ( n141 ) : ( n619 ) ;
assign n621 =  ( n8 ) ? ( n620 ) : ( SREG_27 ) ;
assign n622 =  ( n172 ) ? ( n149 ) : ( SREG_27 ) ;
assign n623 =  ( n170 ) ? ( n171 ) : ( n622 ) ;
assign n624 =  ( n168 ) ? ( n169 ) : ( n623 ) ;
assign n625 =  ( n166 ) ? ( n167 ) : ( n624 ) ;
assign n626 =  ( n162 ) ? ( n165 ) : ( n625 ) ;
assign n627 =  ( n170 ) ? ( n184 ) : ( n622 ) ;
assign n628 =  ( n168 ) ? ( n183 ) : ( n627 ) ;
assign n629 =  ( n166 ) ? ( n182 ) : ( n628 ) ;
assign n630 =  ( n162 ) ? ( n181 ) : ( n629 ) ;
assign n631 =  ( n178 ) ? ( n630 ) : ( SREG_27 ) ;
assign n632 =  ( n159 ) ? ( n626 ) : ( n631 ) ;
assign n633 =  ( n192 ) ? ( SREG_27 ) : ( SREG_27 ) ;
assign n634 =  ( n157 ) ? ( n632 ) : ( n633 ) ;
assign n635 =  ( n6 ) ? ( n621 ) : ( n634 ) ;
assign n636 =  ( n615 ) ? ( n635 ) : ( SREG_27 ) ;
assign n637 =  ( n3 ) == ( 5'd28 )  ;
assign n638 =  ( n148 ) ? ( n149 ) : ( SREG_28 ) ;
assign n639 =  ( n146 ) ? ( n147 ) : ( n638 ) ;
assign n640 =  ( n144 ) ? ( n145 ) : ( n639 ) ;
assign n641 =  ( n142 ) ? ( n143 ) : ( n640 ) ;
assign n642 =  ( n10 ) ? ( n141 ) : ( n641 ) ;
assign n643 =  ( n8 ) ? ( n642 ) : ( SREG_28 ) ;
assign n644 =  ( n172 ) ? ( n149 ) : ( SREG_28 ) ;
assign n645 =  ( n170 ) ? ( n171 ) : ( n644 ) ;
assign n646 =  ( n168 ) ? ( n169 ) : ( n645 ) ;
assign n647 =  ( n166 ) ? ( n167 ) : ( n646 ) ;
assign n648 =  ( n162 ) ? ( n165 ) : ( n647 ) ;
assign n649 =  ( n170 ) ? ( n184 ) : ( n644 ) ;
assign n650 =  ( n168 ) ? ( n183 ) : ( n649 ) ;
assign n651 =  ( n166 ) ? ( n182 ) : ( n650 ) ;
assign n652 =  ( n162 ) ? ( n181 ) : ( n651 ) ;
assign n653 =  ( n178 ) ? ( n652 ) : ( SREG_28 ) ;
assign n654 =  ( n159 ) ? ( n648 ) : ( n653 ) ;
assign n655 =  ( n192 ) ? ( SREG_28 ) : ( SREG_28 ) ;
assign n656 =  ( n157 ) ? ( n654 ) : ( n655 ) ;
assign n657 =  ( n6 ) ? ( n643 ) : ( n656 ) ;
assign n658 =  ( n637 ) ? ( n657 ) : ( SREG_28 ) ;
assign n659 =  ( n3 ) == ( 5'd29 )  ;
assign n660 =  ( n148 ) ? ( n149 ) : ( SREG_29 ) ;
assign n661 =  ( n146 ) ? ( n147 ) : ( n660 ) ;
assign n662 =  ( n144 ) ? ( n145 ) : ( n661 ) ;
assign n663 =  ( n142 ) ? ( n143 ) : ( n662 ) ;
assign n664 =  ( n10 ) ? ( n141 ) : ( n663 ) ;
assign n665 =  ( n8 ) ? ( n664 ) : ( SREG_29 ) ;
assign n666 =  ( n172 ) ? ( n149 ) : ( SREG_29 ) ;
assign n667 =  ( n170 ) ? ( n171 ) : ( n666 ) ;
assign n668 =  ( n168 ) ? ( n169 ) : ( n667 ) ;
assign n669 =  ( n166 ) ? ( n167 ) : ( n668 ) ;
assign n670 =  ( n162 ) ? ( n165 ) : ( n669 ) ;
assign n671 =  ( n170 ) ? ( n184 ) : ( n666 ) ;
assign n672 =  ( n168 ) ? ( n183 ) : ( n671 ) ;
assign n673 =  ( n166 ) ? ( n182 ) : ( n672 ) ;
assign n674 =  ( n162 ) ? ( n181 ) : ( n673 ) ;
assign n675 =  ( n178 ) ? ( n674 ) : ( SREG_29 ) ;
assign n676 =  ( n159 ) ? ( n670 ) : ( n675 ) ;
assign n677 =  ( n192 ) ? ( SREG_29 ) : ( SREG_29 ) ;
assign n678 =  ( n157 ) ? ( n676 ) : ( n677 ) ;
assign n679 =  ( n6 ) ? ( n665 ) : ( n678 ) ;
assign n680 =  ( n659 ) ? ( n679 ) : ( SREG_29 ) ;
assign n681 =  ( n3 ) == ( 5'd3 )  ;
assign n682 =  ( n148 ) ? ( n149 ) : ( SREG_3 ) ;
assign n683 =  ( n146 ) ? ( n147 ) : ( n682 ) ;
assign n684 =  ( n144 ) ? ( n145 ) : ( n683 ) ;
assign n685 =  ( n142 ) ? ( n143 ) : ( n684 ) ;
assign n686 =  ( n10 ) ? ( n141 ) : ( n685 ) ;
assign n687 =  ( n8 ) ? ( n686 ) : ( SREG_3 ) ;
assign n688 =  ( n172 ) ? ( n149 ) : ( SREG_3 ) ;
assign n689 =  ( n170 ) ? ( n171 ) : ( n688 ) ;
assign n690 =  ( n168 ) ? ( n169 ) : ( n689 ) ;
assign n691 =  ( n166 ) ? ( n167 ) : ( n690 ) ;
assign n692 =  ( n162 ) ? ( n165 ) : ( n691 ) ;
assign n693 =  ( n170 ) ? ( n184 ) : ( n688 ) ;
assign n694 =  ( n168 ) ? ( n183 ) : ( n693 ) ;
assign n695 =  ( n166 ) ? ( n182 ) : ( n694 ) ;
assign n696 =  ( n162 ) ? ( n181 ) : ( n695 ) ;
assign n697 =  ( n178 ) ? ( n696 ) : ( SREG_3 ) ;
assign n698 =  ( n159 ) ? ( n692 ) : ( n697 ) ;
assign n699 =  ( n192 ) ? ( SREG_3 ) : ( SREG_3 ) ;
assign n700 =  ( n157 ) ? ( n698 ) : ( n699 ) ;
assign n701 =  ( n6 ) ? ( n687 ) : ( n700 ) ;
assign n702 =  ( n681 ) ? ( n701 ) : ( SREG_3 ) ;
assign n703 =  ( n3 ) == ( 5'd30 )  ;
assign n704 =  ( n148 ) ? ( n149 ) : ( SREG_30 ) ;
assign n705 =  ( n146 ) ? ( n147 ) : ( n704 ) ;
assign n706 =  ( n144 ) ? ( n145 ) : ( n705 ) ;
assign n707 =  ( n142 ) ? ( n143 ) : ( n706 ) ;
assign n708 =  ( n10 ) ? ( n141 ) : ( n707 ) ;
assign n709 =  ( n8 ) ? ( n708 ) : ( SREG_30 ) ;
assign n710 =  ( n172 ) ? ( n149 ) : ( SREG_30 ) ;
assign n711 =  ( n170 ) ? ( n171 ) : ( n710 ) ;
assign n712 =  ( n168 ) ? ( n169 ) : ( n711 ) ;
assign n713 =  ( n166 ) ? ( n167 ) : ( n712 ) ;
assign n714 =  ( n162 ) ? ( n165 ) : ( n713 ) ;
assign n715 =  ( n170 ) ? ( n184 ) : ( n710 ) ;
assign n716 =  ( n168 ) ? ( n183 ) : ( n715 ) ;
assign n717 =  ( n166 ) ? ( n182 ) : ( n716 ) ;
assign n718 =  ( n162 ) ? ( n181 ) : ( n717 ) ;
assign n719 =  ( n178 ) ? ( n718 ) : ( SREG_30 ) ;
assign n720 =  ( n159 ) ? ( n714 ) : ( n719 ) ;
assign n721 =  ( n192 ) ? ( SREG_30 ) : ( SREG_30 ) ;
assign n722 =  ( n157 ) ? ( n720 ) : ( n721 ) ;
assign n723 =  ( n6 ) ? ( n709 ) : ( n722 ) ;
assign n724 =  ( n703 ) ? ( n723 ) : ( SREG_30 ) ;
assign n725 =  ( n3 ) == ( 5'd31 )  ;
assign n726 =  ( n148 ) ? ( n149 ) : ( SREG_31 ) ;
assign n727 =  ( n146 ) ? ( n147 ) : ( n726 ) ;
assign n728 =  ( n144 ) ? ( n145 ) : ( n727 ) ;
assign n729 =  ( n142 ) ? ( n143 ) : ( n728 ) ;
assign n730 =  ( n10 ) ? ( n141 ) : ( n729 ) ;
assign n731 =  ( n8 ) ? ( n730 ) : ( SREG_31 ) ;
assign n732 =  ( n172 ) ? ( n149 ) : ( SREG_31 ) ;
assign n733 =  ( n170 ) ? ( n171 ) : ( n732 ) ;
assign n734 =  ( n168 ) ? ( n169 ) : ( n733 ) ;
assign n735 =  ( n166 ) ? ( n167 ) : ( n734 ) ;
assign n736 =  ( n162 ) ? ( n165 ) : ( n735 ) ;
assign n737 =  ( n170 ) ? ( n184 ) : ( n732 ) ;
assign n738 =  ( n168 ) ? ( n183 ) : ( n737 ) ;
assign n739 =  ( n166 ) ? ( n182 ) : ( n738 ) ;
assign n740 =  ( n162 ) ? ( n181 ) : ( n739 ) ;
assign n741 =  ( n178 ) ? ( n740 ) : ( SREG_31 ) ;
assign n742 =  ( n159 ) ? ( n736 ) : ( n741 ) ;
assign n743 =  ( n192 ) ? ( SREG_31 ) : ( SREG_31 ) ;
assign n744 =  ( n157 ) ? ( n742 ) : ( n743 ) ;
assign n745 =  ( n6 ) ? ( n731 ) : ( n744 ) ;
assign n746 =  ( n725 ) ? ( n745 ) : ( SREG_31 ) ;
assign n747 =  ( n3 ) == ( 5'd4 )  ;
assign n748 =  ( n148 ) ? ( n149 ) : ( SREG_4 ) ;
assign n749 =  ( n146 ) ? ( n147 ) : ( n748 ) ;
assign n750 =  ( n144 ) ? ( n145 ) : ( n749 ) ;
assign n751 =  ( n142 ) ? ( n143 ) : ( n750 ) ;
assign n752 =  ( n10 ) ? ( n141 ) : ( n751 ) ;
assign n753 =  ( n8 ) ? ( n752 ) : ( SREG_4 ) ;
assign n754 =  ( n172 ) ? ( n149 ) : ( SREG_4 ) ;
assign n755 =  ( n170 ) ? ( n171 ) : ( n754 ) ;
assign n756 =  ( n168 ) ? ( n169 ) : ( n755 ) ;
assign n757 =  ( n166 ) ? ( n167 ) : ( n756 ) ;
assign n758 =  ( n162 ) ? ( n165 ) : ( n757 ) ;
assign n759 =  ( n170 ) ? ( n184 ) : ( n754 ) ;
assign n760 =  ( n168 ) ? ( n183 ) : ( n759 ) ;
assign n761 =  ( n166 ) ? ( n182 ) : ( n760 ) ;
assign n762 =  ( n162 ) ? ( n181 ) : ( n761 ) ;
assign n763 =  ( n178 ) ? ( n762 ) : ( SREG_4 ) ;
assign n764 =  ( n159 ) ? ( n758 ) : ( n763 ) ;
assign n765 =  ( n192 ) ? ( SREG_4 ) : ( SREG_4 ) ;
assign n766 =  ( n157 ) ? ( n764 ) : ( n765 ) ;
assign n767 =  ( n6 ) ? ( n753 ) : ( n766 ) ;
assign n768 =  ( n747 ) ? ( n767 ) : ( SREG_4 ) ;
assign n769 =  ( n3 ) == ( 5'd5 )  ;
assign n770 =  ( n148 ) ? ( n149 ) : ( SREG_5 ) ;
assign n771 =  ( n146 ) ? ( n147 ) : ( n770 ) ;
assign n772 =  ( n144 ) ? ( n145 ) : ( n771 ) ;
assign n773 =  ( n142 ) ? ( n143 ) : ( n772 ) ;
assign n774 =  ( n10 ) ? ( n141 ) : ( n773 ) ;
assign n775 =  ( n8 ) ? ( n774 ) : ( SREG_5 ) ;
assign n776 =  ( n172 ) ? ( n149 ) : ( SREG_5 ) ;
assign n777 =  ( n170 ) ? ( n171 ) : ( n776 ) ;
assign n778 =  ( n168 ) ? ( n169 ) : ( n777 ) ;
assign n779 =  ( n166 ) ? ( n167 ) : ( n778 ) ;
assign n780 =  ( n162 ) ? ( n165 ) : ( n779 ) ;
assign n781 =  ( n170 ) ? ( n184 ) : ( n776 ) ;
assign n782 =  ( n168 ) ? ( n183 ) : ( n781 ) ;
assign n783 =  ( n166 ) ? ( n182 ) : ( n782 ) ;
assign n784 =  ( n162 ) ? ( n181 ) : ( n783 ) ;
assign n785 =  ( n178 ) ? ( n784 ) : ( SREG_5 ) ;
assign n786 =  ( n159 ) ? ( n780 ) : ( n785 ) ;
assign n787 =  ( n192 ) ? ( SREG_5 ) : ( SREG_5 ) ;
assign n788 =  ( n157 ) ? ( n786 ) : ( n787 ) ;
assign n789 =  ( n6 ) ? ( n775 ) : ( n788 ) ;
assign n790 =  ( n769 ) ? ( n789 ) : ( SREG_5 ) ;
assign n791 =  ( n3 ) == ( 5'd6 )  ;
assign n792 =  ( n148 ) ? ( n149 ) : ( SREG_6 ) ;
assign n793 =  ( n146 ) ? ( n147 ) : ( n792 ) ;
assign n794 =  ( n144 ) ? ( n145 ) : ( n793 ) ;
assign n795 =  ( n142 ) ? ( n143 ) : ( n794 ) ;
assign n796 =  ( n10 ) ? ( n141 ) : ( n795 ) ;
assign n797 =  ( n8 ) ? ( n796 ) : ( SREG_6 ) ;
assign n798 =  ( n172 ) ? ( n149 ) : ( SREG_6 ) ;
assign n799 =  ( n170 ) ? ( n171 ) : ( n798 ) ;
assign n800 =  ( n168 ) ? ( n169 ) : ( n799 ) ;
assign n801 =  ( n166 ) ? ( n167 ) : ( n800 ) ;
assign n802 =  ( n162 ) ? ( n165 ) : ( n801 ) ;
assign n803 =  ( n170 ) ? ( n184 ) : ( n798 ) ;
assign n804 =  ( n168 ) ? ( n183 ) : ( n803 ) ;
assign n805 =  ( n166 ) ? ( n182 ) : ( n804 ) ;
assign n806 =  ( n162 ) ? ( n181 ) : ( n805 ) ;
assign n807 =  ( n178 ) ? ( n806 ) : ( SREG_6 ) ;
assign n808 =  ( n159 ) ? ( n802 ) : ( n807 ) ;
assign n809 =  ( n192 ) ? ( SREG_6 ) : ( SREG_6 ) ;
assign n810 =  ( n157 ) ? ( n808 ) : ( n809 ) ;
assign n811 =  ( n6 ) ? ( n797 ) : ( n810 ) ;
assign n812 =  ( n791 ) ? ( n811 ) : ( SREG_6 ) ;
assign n813 =  ( n3 ) == ( 5'd7 )  ;
assign n814 =  ( n148 ) ? ( n149 ) : ( SREG_7 ) ;
assign n815 =  ( n146 ) ? ( n147 ) : ( n814 ) ;
assign n816 =  ( n144 ) ? ( n145 ) : ( n815 ) ;
assign n817 =  ( n142 ) ? ( n143 ) : ( n816 ) ;
assign n818 =  ( n10 ) ? ( n141 ) : ( n817 ) ;
assign n819 =  ( n8 ) ? ( n818 ) : ( SREG_7 ) ;
assign n820 =  ( n172 ) ? ( n149 ) : ( SREG_7 ) ;
assign n821 =  ( n170 ) ? ( n171 ) : ( n820 ) ;
assign n822 =  ( n168 ) ? ( n169 ) : ( n821 ) ;
assign n823 =  ( n166 ) ? ( n167 ) : ( n822 ) ;
assign n824 =  ( n162 ) ? ( n165 ) : ( n823 ) ;
assign n825 =  ( n170 ) ? ( n184 ) : ( n820 ) ;
assign n826 =  ( n168 ) ? ( n183 ) : ( n825 ) ;
assign n827 =  ( n166 ) ? ( n182 ) : ( n826 ) ;
assign n828 =  ( n162 ) ? ( n181 ) : ( n827 ) ;
assign n829 =  ( n178 ) ? ( n828 ) : ( SREG_7 ) ;
assign n830 =  ( n159 ) ? ( n824 ) : ( n829 ) ;
assign n831 =  ( n192 ) ? ( SREG_7 ) : ( SREG_7 ) ;
assign n832 =  ( n157 ) ? ( n830 ) : ( n831 ) ;
assign n833 =  ( n6 ) ? ( n819 ) : ( n832 ) ;
assign n834 =  ( n813 ) ? ( n833 ) : ( SREG_7 ) ;
assign n835 =  ( n3 ) == ( 5'd8 )  ;
assign n836 =  ( n148 ) ? ( n149 ) : ( SREG_8 ) ;
assign n837 =  ( n146 ) ? ( n147 ) : ( n836 ) ;
assign n838 =  ( n144 ) ? ( n145 ) : ( n837 ) ;
assign n839 =  ( n142 ) ? ( n143 ) : ( n838 ) ;
assign n840 =  ( n10 ) ? ( n141 ) : ( n839 ) ;
assign n841 =  ( n8 ) ? ( n840 ) : ( SREG_8 ) ;
assign n842 =  ( n172 ) ? ( n149 ) : ( SREG_8 ) ;
assign n843 =  ( n170 ) ? ( n171 ) : ( n842 ) ;
assign n844 =  ( n168 ) ? ( n169 ) : ( n843 ) ;
assign n845 =  ( n166 ) ? ( n167 ) : ( n844 ) ;
assign n846 =  ( n162 ) ? ( n165 ) : ( n845 ) ;
assign n847 =  ( n170 ) ? ( n184 ) : ( n842 ) ;
assign n848 =  ( n168 ) ? ( n183 ) : ( n847 ) ;
assign n849 =  ( n166 ) ? ( n182 ) : ( n848 ) ;
assign n850 =  ( n162 ) ? ( n181 ) : ( n849 ) ;
assign n851 =  ( n178 ) ? ( n850 ) : ( SREG_8 ) ;
assign n852 =  ( n159 ) ? ( n846 ) : ( n851 ) ;
assign n853 =  ( n192 ) ? ( SREG_8 ) : ( SREG_8 ) ;
assign n854 =  ( n157 ) ? ( n852 ) : ( n853 ) ;
assign n855 =  ( n6 ) ? ( n841 ) : ( n854 ) ;
assign n856 =  ( n835 ) ? ( n855 ) : ( SREG_8 ) ;
assign n857 =  ( n3 ) == ( 5'd9 )  ;
assign n858 =  ( n148 ) ? ( n149 ) : ( SREG_9 ) ;
assign n859 =  ( n146 ) ? ( n147 ) : ( n858 ) ;
assign n860 =  ( n144 ) ? ( n145 ) : ( n859 ) ;
assign n861 =  ( n142 ) ? ( n143 ) : ( n860 ) ;
assign n862 =  ( n10 ) ? ( n141 ) : ( n861 ) ;
assign n863 =  ( n8 ) ? ( n862 ) : ( SREG_9 ) ;
assign n864 =  ( n172 ) ? ( n149 ) : ( SREG_9 ) ;
assign n865 =  ( n170 ) ? ( n171 ) : ( n864 ) ;
assign n866 =  ( n168 ) ? ( n169 ) : ( n865 ) ;
assign n867 =  ( n166 ) ? ( n167 ) : ( n866 ) ;
assign n868 =  ( n162 ) ? ( n165 ) : ( n867 ) ;
assign n869 =  ( n170 ) ? ( n184 ) : ( n864 ) ;
assign n870 =  ( n168 ) ? ( n183 ) : ( n869 ) ;
assign n871 =  ( n166 ) ? ( n182 ) : ( n870 ) ;
assign n872 =  ( n162 ) ? ( n181 ) : ( n871 ) ;
assign n873 =  ( n178 ) ? ( n872 ) : ( SREG_9 ) ;
assign n874 =  ( n159 ) ? ( n868 ) : ( n873 ) ;
assign n875 =  ( n192 ) ? ( SREG_9 ) : ( SREG_9 ) ;
assign n876 =  ( n157 ) ? ( n874 ) : ( n875 ) ;
assign n877 =  ( n6 ) ? ( n863 ) : ( n876 ) ;
assign n878 =  ( n857 ) ? ( n877 ) : ( SREG_9 ) ;
assign n879 =  ( n7 ) == ( 3'd1 )  ;
assign n880 =  ( 32'd0 ) == ( 32'd15 )  ;
assign n881 =  ( n12 ) & ( n880 )  ;
assign n882 =  ( 32'd0 ) == ( 32'd14 )  ;
assign n883 =  ( n12 ) & ( n882 )  ;
assign n884 =  ( 32'd0 ) == ( 32'd13 )  ;
assign n885 =  ( n12 ) & ( n884 )  ;
assign n886 =  ( 32'd0 ) == ( 32'd12 )  ;
assign n887 =  ( n12 ) & ( n886 )  ;
assign n888 =  ( 32'd0 ) == ( 32'd11 )  ;
assign n889 =  ( n12 ) & ( n888 )  ;
assign n890 =  ( 32'd0 ) == ( 32'd10 )  ;
assign n891 =  ( n12 ) & ( n890 )  ;
assign n892 =  ( 32'd0 ) == ( 32'd9 )  ;
assign n893 =  ( n12 ) & ( n892 )  ;
assign n894 =  ( 32'd0 ) == ( 32'd8 )  ;
assign n895 =  ( n12 ) & ( n894 )  ;
assign n896 =  ( 32'd0 ) == ( 32'd7 )  ;
assign n897 =  ( n12 ) & ( n896 )  ;
assign n898 =  ( 32'd0 ) == ( 32'd6 )  ;
assign n899 =  ( n12 ) & ( n898 )  ;
assign n900 =  ( 32'd0 ) == ( 32'd5 )  ;
assign n901 =  ( n12 ) & ( n900 )  ;
assign n902 =  ( 32'd0 ) == ( 32'd4 )  ;
assign n903 =  ( n12 ) & ( n902 )  ;
assign n904 =  ( 32'd0 ) == ( 32'd3 )  ;
assign n905 =  ( n12 ) & ( n904 )  ;
assign n906 =  ( 32'd0 ) == ( 32'd2 )  ;
assign n907 =  ( n12 ) & ( n906 )  ;
assign n908 =  ( 32'd0 ) == ( 32'd1 )  ;
assign n909 =  ( n12 ) & ( n908 )  ;
assign n910 =  ( 32'd0 ) == ( 32'd0 )  ;
assign n911 =  ( n12 ) & ( n910 )  ;
assign n912 =  ( n13 ) & ( n880 )  ;
assign n913 =  ( n13 ) & ( n882 )  ;
assign n914 =  ( n13 ) & ( n884 )  ;
assign n915 =  ( n13 ) & ( n886 )  ;
assign n916 =  ( n13 ) & ( n888 )  ;
assign n917 =  ( n13 ) & ( n890 )  ;
assign n918 =  ( n13 ) & ( n892 )  ;
assign n919 =  ( n13 ) & ( n894 )  ;
assign n920 =  ( n13 ) & ( n896 )  ;
assign n921 =  ( n13 ) & ( n898 )  ;
assign n922 =  ( n13 ) & ( n900 )  ;
assign n923 =  ( n13 ) & ( n902 )  ;
assign n924 =  ( n13 ) & ( n904 )  ;
assign n925 =  ( n13 ) & ( n906 )  ;
assign n926 =  ( n13 ) & ( n908 )  ;
assign n927 =  ( n13 ) & ( n910 )  ;
assign n928 =  ( n14 ) & ( n880 )  ;
assign n929 =  ( n14 ) & ( n882 )  ;
assign n930 =  ( n14 ) & ( n884 )  ;
assign n931 =  ( n14 ) & ( n886 )  ;
assign n932 =  ( n14 ) & ( n888 )  ;
assign n933 =  ( n14 ) & ( n890 )  ;
assign n934 =  ( n14 ) & ( n892 )  ;
assign n935 =  ( n14 ) & ( n894 )  ;
assign n936 =  ( n14 ) & ( n896 )  ;
assign n937 =  ( n14 ) & ( n898 )  ;
assign n938 =  ( n14 ) & ( n900 )  ;
assign n939 =  ( n14 ) & ( n902 )  ;
assign n940 =  ( n14 ) & ( n904 )  ;
assign n941 =  ( n14 ) & ( n906 )  ;
assign n942 =  ( n14 ) & ( n908 )  ;
assign n943 =  ( n14 ) & ( n910 )  ;
assign n944 =  ( n15 ) & ( n880 )  ;
assign n945 =  ( n15 ) & ( n882 )  ;
assign n946 =  ( n15 ) & ( n884 )  ;
assign n947 =  ( n15 ) & ( n886 )  ;
assign n948 =  ( n15 ) & ( n888 )  ;
assign n949 =  ( n15 ) & ( n890 )  ;
assign n950 =  ( n15 ) & ( n892 )  ;
assign n951 =  ( n15 ) & ( n894 )  ;
assign n952 =  ( n15 ) & ( n896 )  ;
assign n953 =  ( n15 ) & ( n898 )  ;
assign n954 =  ( n15 ) & ( n900 )  ;
assign n955 =  ( n15 ) & ( n902 )  ;
assign n956 =  ( n15 ) & ( n904 )  ;
assign n957 =  ( n15 ) & ( n906 )  ;
assign n958 =  ( n15 ) & ( n908 )  ;
assign n959 =  ( n15 ) & ( n910 )  ;
assign n960 =  ( n16 ) & ( n880 )  ;
assign n961 =  ( n16 ) & ( n882 )  ;
assign n962 =  ( n16 ) & ( n884 )  ;
assign n963 =  ( n16 ) & ( n886 )  ;
assign n964 =  ( n16 ) & ( n888 )  ;
assign n965 =  ( n16 ) & ( n890 )  ;
assign n966 =  ( n16 ) & ( n892 )  ;
assign n967 =  ( n16 ) & ( n894 )  ;
assign n968 =  ( n16 ) & ( n896 )  ;
assign n969 =  ( n16 ) & ( n898 )  ;
assign n970 =  ( n16 ) & ( n900 )  ;
assign n971 =  ( n16 ) & ( n902 )  ;
assign n972 =  ( n16 ) & ( n904 )  ;
assign n973 =  ( n16 ) & ( n906 )  ;
assign n974 =  ( n16 ) & ( n908 )  ;
assign n975 =  ( n16 ) & ( n910 )  ;
assign n976 =  ( n17 ) & ( n880 )  ;
assign n977 =  ( n17 ) & ( n882 )  ;
assign n978 =  ( n17 ) & ( n884 )  ;
assign n979 =  ( n17 ) & ( n886 )  ;
assign n980 =  ( n17 ) & ( n888 )  ;
assign n981 =  ( n17 ) & ( n890 )  ;
assign n982 =  ( n17 ) & ( n892 )  ;
assign n983 =  ( n17 ) & ( n894 )  ;
assign n984 =  ( n17 ) & ( n896 )  ;
assign n985 =  ( n17 ) & ( n898 )  ;
assign n986 =  ( n17 ) & ( n900 )  ;
assign n987 =  ( n17 ) & ( n902 )  ;
assign n988 =  ( n17 ) & ( n904 )  ;
assign n989 =  ( n17 ) & ( n906 )  ;
assign n990 =  ( n17 ) & ( n908 )  ;
assign n991 =  ( n17 ) & ( n910 )  ;
assign n992 =  ( n18 ) & ( n880 )  ;
assign n993 =  ( n18 ) & ( n882 )  ;
assign n994 =  ( n18 ) & ( n884 )  ;
assign n995 =  ( n18 ) & ( n886 )  ;
assign n996 =  ( n18 ) & ( n888 )  ;
assign n997 =  ( n18 ) & ( n890 )  ;
assign n998 =  ( n18 ) & ( n892 )  ;
assign n999 =  ( n18 ) & ( n894 )  ;
assign n1000 =  ( n18 ) & ( n896 )  ;
assign n1001 =  ( n18 ) & ( n898 )  ;
assign n1002 =  ( n18 ) & ( n900 )  ;
assign n1003 =  ( n18 ) & ( n902 )  ;
assign n1004 =  ( n18 ) & ( n904 )  ;
assign n1005 =  ( n18 ) & ( n906 )  ;
assign n1006 =  ( n18 ) & ( n908 )  ;
assign n1007 =  ( n18 ) & ( n910 )  ;
assign n1008 =  ( n19 ) & ( n880 )  ;
assign n1009 =  ( n19 ) & ( n882 )  ;
assign n1010 =  ( n19 ) & ( n884 )  ;
assign n1011 =  ( n19 ) & ( n886 )  ;
assign n1012 =  ( n19 ) & ( n888 )  ;
assign n1013 =  ( n19 ) & ( n890 )  ;
assign n1014 =  ( n19 ) & ( n892 )  ;
assign n1015 =  ( n19 ) & ( n894 )  ;
assign n1016 =  ( n19 ) & ( n896 )  ;
assign n1017 =  ( n19 ) & ( n898 )  ;
assign n1018 =  ( n19 ) & ( n900 )  ;
assign n1019 =  ( n19 ) & ( n902 )  ;
assign n1020 =  ( n19 ) & ( n904 )  ;
assign n1021 =  ( n19 ) & ( n906 )  ;
assign n1022 =  ( n19 ) & ( n908 )  ;
assign n1023 =  ( n19 ) & ( n910 )  ;
assign n1024 =  ( n20 ) & ( n880 )  ;
assign n1025 =  ( n20 ) & ( n882 )  ;
assign n1026 =  ( n20 ) & ( n884 )  ;
assign n1027 =  ( n20 ) & ( n886 )  ;
assign n1028 =  ( n20 ) & ( n888 )  ;
assign n1029 =  ( n20 ) & ( n890 )  ;
assign n1030 =  ( n20 ) & ( n892 )  ;
assign n1031 =  ( n20 ) & ( n894 )  ;
assign n1032 =  ( n20 ) & ( n896 )  ;
assign n1033 =  ( n20 ) & ( n898 )  ;
assign n1034 =  ( n20 ) & ( n900 )  ;
assign n1035 =  ( n20 ) & ( n902 )  ;
assign n1036 =  ( n20 ) & ( n904 )  ;
assign n1037 =  ( n20 ) & ( n906 )  ;
assign n1038 =  ( n20 ) & ( n908 )  ;
assign n1039 =  ( n20 ) & ( n910 )  ;
assign n1040 =  ( n21 ) & ( n880 )  ;
assign n1041 =  ( n21 ) & ( n882 )  ;
assign n1042 =  ( n21 ) & ( n884 )  ;
assign n1043 =  ( n21 ) & ( n886 )  ;
assign n1044 =  ( n21 ) & ( n888 )  ;
assign n1045 =  ( n21 ) & ( n890 )  ;
assign n1046 =  ( n21 ) & ( n892 )  ;
assign n1047 =  ( n21 ) & ( n894 )  ;
assign n1048 =  ( n21 ) & ( n896 )  ;
assign n1049 =  ( n21 ) & ( n898 )  ;
assign n1050 =  ( n21 ) & ( n900 )  ;
assign n1051 =  ( n21 ) & ( n902 )  ;
assign n1052 =  ( n21 ) & ( n904 )  ;
assign n1053 =  ( n21 ) & ( n906 )  ;
assign n1054 =  ( n21 ) & ( n908 )  ;
assign n1055 =  ( n21 ) & ( n910 )  ;
assign n1056 =  ( n22 ) & ( n880 )  ;
assign n1057 =  ( n22 ) & ( n882 )  ;
assign n1058 =  ( n22 ) & ( n884 )  ;
assign n1059 =  ( n22 ) & ( n886 )  ;
assign n1060 =  ( n22 ) & ( n888 )  ;
assign n1061 =  ( n22 ) & ( n890 )  ;
assign n1062 =  ( n22 ) & ( n892 )  ;
assign n1063 =  ( n22 ) & ( n894 )  ;
assign n1064 =  ( n22 ) & ( n896 )  ;
assign n1065 =  ( n22 ) & ( n898 )  ;
assign n1066 =  ( n22 ) & ( n900 )  ;
assign n1067 =  ( n22 ) & ( n902 )  ;
assign n1068 =  ( n22 ) & ( n904 )  ;
assign n1069 =  ( n22 ) & ( n906 )  ;
assign n1070 =  ( n22 ) & ( n908 )  ;
assign n1071 =  ( n22 ) & ( n910 )  ;
assign n1072 =  ( n23 ) & ( n880 )  ;
assign n1073 =  ( n23 ) & ( n882 )  ;
assign n1074 =  ( n23 ) & ( n884 )  ;
assign n1075 =  ( n23 ) & ( n886 )  ;
assign n1076 =  ( n23 ) & ( n888 )  ;
assign n1077 =  ( n23 ) & ( n890 )  ;
assign n1078 =  ( n23 ) & ( n892 )  ;
assign n1079 =  ( n23 ) & ( n894 )  ;
assign n1080 =  ( n23 ) & ( n896 )  ;
assign n1081 =  ( n23 ) & ( n898 )  ;
assign n1082 =  ( n23 ) & ( n900 )  ;
assign n1083 =  ( n23 ) & ( n902 )  ;
assign n1084 =  ( n23 ) & ( n904 )  ;
assign n1085 =  ( n23 ) & ( n906 )  ;
assign n1086 =  ( n23 ) & ( n908 )  ;
assign n1087 =  ( n23 ) & ( n910 )  ;
assign n1088 =  ( n24 ) & ( n880 )  ;
assign n1089 =  ( n24 ) & ( n882 )  ;
assign n1090 =  ( n24 ) & ( n884 )  ;
assign n1091 =  ( n24 ) & ( n886 )  ;
assign n1092 =  ( n24 ) & ( n888 )  ;
assign n1093 =  ( n24 ) & ( n890 )  ;
assign n1094 =  ( n24 ) & ( n892 )  ;
assign n1095 =  ( n24 ) & ( n894 )  ;
assign n1096 =  ( n24 ) & ( n896 )  ;
assign n1097 =  ( n24 ) & ( n898 )  ;
assign n1098 =  ( n24 ) & ( n900 )  ;
assign n1099 =  ( n24 ) & ( n902 )  ;
assign n1100 =  ( n24 ) & ( n904 )  ;
assign n1101 =  ( n24 ) & ( n906 )  ;
assign n1102 =  ( n24 ) & ( n908 )  ;
assign n1103 =  ( n24 ) & ( n910 )  ;
assign n1104 =  ( n25 ) & ( n880 )  ;
assign n1105 =  ( n25 ) & ( n882 )  ;
assign n1106 =  ( n25 ) & ( n884 )  ;
assign n1107 =  ( n25 ) & ( n886 )  ;
assign n1108 =  ( n25 ) & ( n888 )  ;
assign n1109 =  ( n25 ) & ( n890 )  ;
assign n1110 =  ( n25 ) & ( n892 )  ;
assign n1111 =  ( n25 ) & ( n894 )  ;
assign n1112 =  ( n25 ) & ( n896 )  ;
assign n1113 =  ( n25 ) & ( n898 )  ;
assign n1114 =  ( n25 ) & ( n900 )  ;
assign n1115 =  ( n25 ) & ( n902 )  ;
assign n1116 =  ( n25 ) & ( n904 )  ;
assign n1117 =  ( n25 ) & ( n906 )  ;
assign n1118 =  ( n25 ) & ( n908 )  ;
assign n1119 =  ( n25 ) & ( n910 )  ;
assign n1120 =  ( n26 ) & ( n880 )  ;
assign n1121 =  ( n26 ) & ( n882 )  ;
assign n1122 =  ( n26 ) & ( n884 )  ;
assign n1123 =  ( n26 ) & ( n886 )  ;
assign n1124 =  ( n26 ) & ( n888 )  ;
assign n1125 =  ( n26 ) & ( n890 )  ;
assign n1126 =  ( n26 ) & ( n892 )  ;
assign n1127 =  ( n26 ) & ( n894 )  ;
assign n1128 =  ( n26 ) & ( n896 )  ;
assign n1129 =  ( n26 ) & ( n898 )  ;
assign n1130 =  ( n26 ) & ( n900 )  ;
assign n1131 =  ( n26 ) & ( n902 )  ;
assign n1132 =  ( n26 ) & ( n904 )  ;
assign n1133 =  ( n26 ) & ( n906 )  ;
assign n1134 =  ( n26 ) & ( n908 )  ;
assign n1135 =  ( n26 ) & ( n910 )  ;
assign n1136 =  ( n27 ) & ( n880 )  ;
assign n1137 =  ( n27 ) & ( n882 )  ;
assign n1138 =  ( n27 ) & ( n884 )  ;
assign n1139 =  ( n27 ) & ( n886 )  ;
assign n1140 =  ( n27 ) & ( n888 )  ;
assign n1141 =  ( n27 ) & ( n890 )  ;
assign n1142 =  ( n27 ) & ( n892 )  ;
assign n1143 =  ( n27 ) & ( n894 )  ;
assign n1144 =  ( n27 ) & ( n896 )  ;
assign n1145 =  ( n27 ) & ( n898 )  ;
assign n1146 =  ( n27 ) & ( n900 )  ;
assign n1147 =  ( n27 ) & ( n902 )  ;
assign n1148 =  ( n27 ) & ( n904 )  ;
assign n1149 =  ( n27 ) & ( n906 )  ;
assign n1150 =  ( n27 ) & ( n908 )  ;
assign n1151 =  ( n27 ) & ( n910 )  ;
assign n1152 =  ( n28 ) & ( n880 )  ;
assign n1153 =  ( n28 ) & ( n882 )  ;
assign n1154 =  ( n28 ) & ( n884 )  ;
assign n1155 =  ( n28 ) & ( n886 )  ;
assign n1156 =  ( n28 ) & ( n888 )  ;
assign n1157 =  ( n28 ) & ( n890 )  ;
assign n1158 =  ( n28 ) & ( n892 )  ;
assign n1159 =  ( n28 ) & ( n894 )  ;
assign n1160 =  ( n28 ) & ( n896 )  ;
assign n1161 =  ( n28 ) & ( n898 )  ;
assign n1162 =  ( n28 ) & ( n900 )  ;
assign n1163 =  ( n28 ) & ( n902 )  ;
assign n1164 =  ( n28 ) & ( n904 )  ;
assign n1165 =  ( n28 ) & ( n906 )  ;
assign n1166 =  ( n28 ) & ( n908 )  ;
assign n1167 =  ( n28 ) & ( n910 )  ;
assign n1168 =  ( n29 ) & ( n880 )  ;
assign n1169 =  ( n29 ) & ( n882 )  ;
assign n1170 =  ( n29 ) & ( n884 )  ;
assign n1171 =  ( n29 ) & ( n886 )  ;
assign n1172 =  ( n29 ) & ( n888 )  ;
assign n1173 =  ( n29 ) & ( n890 )  ;
assign n1174 =  ( n29 ) & ( n892 )  ;
assign n1175 =  ( n29 ) & ( n894 )  ;
assign n1176 =  ( n29 ) & ( n896 )  ;
assign n1177 =  ( n29 ) & ( n898 )  ;
assign n1178 =  ( n29 ) & ( n900 )  ;
assign n1179 =  ( n29 ) & ( n902 )  ;
assign n1180 =  ( n29 ) & ( n904 )  ;
assign n1181 =  ( n29 ) & ( n906 )  ;
assign n1182 =  ( n29 ) & ( n908 )  ;
assign n1183 =  ( n29 ) & ( n910 )  ;
assign n1184 =  ( n30 ) & ( n880 )  ;
assign n1185 =  ( n30 ) & ( n882 )  ;
assign n1186 =  ( n30 ) & ( n884 )  ;
assign n1187 =  ( n30 ) & ( n886 )  ;
assign n1188 =  ( n30 ) & ( n888 )  ;
assign n1189 =  ( n30 ) & ( n890 )  ;
assign n1190 =  ( n30 ) & ( n892 )  ;
assign n1191 =  ( n30 ) & ( n894 )  ;
assign n1192 =  ( n30 ) & ( n896 )  ;
assign n1193 =  ( n30 ) & ( n898 )  ;
assign n1194 =  ( n30 ) & ( n900 )  ;
assign n1195 =  ( n30 ) & ( n902 )  ;
assign n1196 =  ( n30 ) & ( n904 )  ;
assign n1197 =  ( n30 ) & ( n906 )  ;
assign n1198 =  ( n30 ) & ( n908 )  ;
assign n1199 =  ( n30 ) & ( n910 )  ;
assign n1200 =  ( n31 ) & ( n880 )  ;
assign n1201 =  ( n31 ) & ( n882 )  ;
assign n1202 =  ( n31 ) & ( n884 )  ;
assign n1203 =  ( n31 ) & ( n886 )  ;
assign n1204 =  ( n31 ) & ( n888 )  ;
assign n1205 =  ( n31 ) & ( n890 )  ;
assign n1206 =  ( n31 ) & ( n892 )  ;
assign n1207 =  ( n31 ) & ( n894 )  ;
assign n1208 =  ( n31 ) & ( n896 )  ;
assign n1209 =  ( n31 ) & ( n898 )  ;
assign n1210 =  ( n31 ) & ( n900 )  ;
assign n1211 =  ( n31 ) & ( n902 )  ;
assign n1212 =  ( n31 ) & ( n904 )  ;
assign n1213 =  ( n31 ) & ( n906 )  ;
assign n1214 =  ( n31 ) & ( n908 )  ;
assign n1215 =  ( n31 ) & ( n910 )  ;
assign n1216 =  ( n32 ) & ( n880 )  ;
assign n1217 =  ( n32 ) & ( n882 )  ;
assign n1218 =  ( n32 ) & ( n884 )  ;
assign n1219 =  ( n32 ) & ( n886 )  ;
assign n1220 =  ( n32 ) & ( n888 )  ;
assign n1221 =  ( n32 ) & ( n890 )  ;
assign n1222 =  ( n32 ) & ( n892 )  ;
assign n1223 =  ( n32 ) & ( n894 )  ;
assign n1224 =  ( n32 ) & ( n896 )  ;
assign n1225 =  ( n32 ) & ( n898 )  ;
assign n1226 =  ( n32 ) & ( n900 )  ;
assign n1227 =  ( n32 ) & ( n902 )  ;
assign n1228 =  ( n32 ) & ( n904 )  ;
assign n1229 =  ( n32 ) & ( n906 )  ;
assign n1230 =  ( n32 ) & ( n908 )  ;
assign n1231 =  ( n32 ) & ( n910 )  ;
assign n1232 =  ( n33 ) & ( n880 )  ;
assign n1233 =  ( n33 ) & ( n882 )  ;
assign n1234 =  ( n33 ) & ( n884 )  ;
assign n1235 =  ( n33 ) & ( n886 )  ;
assign n1236 =  ( n33 ) & ( n888 )  ;
assign n1237 =  ( n33 ) & ( n890 )  ;
assign n1238 =  ( n33 ) & ( n892 )  ;
assign n1239 =  ( n33 ) & ( n894 )  ;
assign n1240 =  ( n33 ) & ( n896 )  ;
assign n1241 =  ( n33 ) & ( n898 )  ;
assign n1242 =  ( n33 ) & ( n900 )  ;
assign n1243 =  ( n33 ) & ( n902 )  ;
assign n1244 =  ( n33 ) & ( n904 )  ;
assign n1245 =  ( n33 ) & ( n906 )  ;
assign n1246 =  ( n33 ) & ( n908 )  ;
assign n1247 =  ( n33 ) & ( n910 )  ;
assign n1248 =  ( n34 ) & ( n880 )  ;
assign n1249 =  ( n34 ) & ( n882 )  ;
assign n1250 =  ( n34 ) & ( n884 )  ;
assign n1251 =  ( n34 ) & ( n886 )  ;
assign n1252 =  ( n34 ) & ( n888 )  ;
assign n1253 =  ( n34 ) & ( n890 )  ;
assign n1254 =  ( n34 ) & ( n892 )  ;
assign n1255 =  ( n34 ) & ( n894 )  ;
assign n1256 =  ( n34 ) & ( n896 )  ;
assign n1257 =  ( n34 ) & ( n898 )  ;
assign n1258 =  ( n34 ) & ( n900 )  ;
assign n1259 =  ( n34 ) & ( n902 )  ;
assign n1260 =  ( n34 ) & ( n904 )  ;
assign n1261 =  ( n34 ) & ( n906 )  ;
assign n1262 =  ( n34 ) & ( n908 )  ;
assign n1263 =  ( n34 ) & ( n910 )  ;
assign n1264 =  ( n35 ) & ( n880 )  ;
assign n1265 =  ( n35 ) & ( n882 )  ;
assign n1266 =  ( n35 ) & ( n884 )  ;
assign n1267 =  ( n35 ) & ( n886 )  ;
assign n1268 =  ( n35 ) & ( n888 )  ;
assign n1269 =  ( n35 ) & ( n890 )  ;
assign n1270 =  ( n35 ) & ( n892 )  ;
assign n1271 =  ( n35 ) & ( n894 )  ;
assign n1272 =  ( n35 ) & ( n896 )  ;
assign n1273 =  ( n35 ) & ( n898 )  ;
assign n1274 =  ( n35 ) & ( n900 )  ;
assign n1275 =  ( n35 ) & ( n902 )  ;
assign n1276 =  ( n35 ) & ( n904 )  ;
assign n1277 =  ( n35 ) & ( n906 )  ;
assign n1278 =  ( n35 ) & ( n908 )  ;
assign n1279 =  ( n35 ) & ( n910 )  ;
assign n1280 =  ( n36 ) & ( n880 )  ;
assign n1281 =  ( n36 ) & ( n882 )  ;
assign n1282 =  ( n36 ) & ( n884 )  ;
assign n1283 =  ( n36 ) & ( n886 )  ;
assign n1284 =  ( n36 ) & ( n888 )  ;
assign n1285 =  ( n36 ) & ( n890 )  ;
assign n1286 =  ( n36 ) & ( n892 )  ;
assign n1287 =  ( n36 ) & ( n894 )  ;
assign n1288 =  ( n36 ) & ( n896 )  ;
assign n1289 =  ( n36 ) & ( n898 )  ;
assign n1290 =  ( n36 ) & ( n900 )  ;
assign n1291 =  ( n36 ) & ( n902 )  ;
assign n1292 =  ( n36 ) & ( n904 )  ;
assign n1293 =  ( n36 ) & ( n906 )  ;
assign n1294 =  ( n36 ) & ( n908 )  ;
assign n1295 =  ( n36 ) & ( n910 )  ;
assign n1296 =  ( n37 ) & ( n880 )  ;
assign n1297 =  ( n37 ) & ( n882 )  ;
assign n1298 =  ( n37 ) & ( n884 )  ;
assign n1299 =  ( n37 ) & ( n886 )  ;
assign n1300 =  ( n37 ) & ( n888 )  ;
assign n1301 =  ( n37 ) & ( n890 )  ;
assign n1302 =  ( n37 ) & ( n892 )  ;
assign n1303 =  ( n37 ) & ( n894 )  ;
assign n1304 =  ( n37 ) & ( n896 )  ;
assign n1305 =  ( n37 ) & ( n898 )  ;
assign n1306 =  ( n37 ) & ( n900 )  ;
assign n1307 =  ( n37 ) & ( n902 )  ;
assign n1308 =  ( n37 ) & ( n904 )  ;
assign n1309 =  ( n37 ) & ( n906 )  ;
assign n1310 =  ( n37 ) & ( n908 )  ;
assign n1311 =  ( n37 ) & ( n910 )  ;
assign n1312 =  ( n38 ) & ( n880 )  ;
assign n1313 =  ( n38 ) & ( n882 )  ;
assign n1314 =  ( n38 ) & ( n884 )  ;
assign n1315 =  ( n38 ) & ( n886 )  ;
assign n1316 =  ( n38 ) & ( n888 )  ;
assign n1317 =  ( n38 ) & ( n890 )  ;
assign n1318 =  ( n38 ) & ( n892 )  ;
assign n1319 =  ( n38 ) & ( n894 )  ;
assign n1320 =  ( n38 ) & ( n896 )  ;
assign n1321 =  ( n38 ) & ( n898 )  ;
assign n1322 =  ( n38 ) & ( n900 )  ;
assign n1323 =  ( n38 ) & ( n902 )  ;
assign n1324 =  ( n38 ) & ( n904 )  ;
assign n1325 =  ( n38 ) & ( n906 )  ;
assign n1326 =  ( n38 ) & ( n908 )  ;
assign n1327 =  ( n38 ) & ( n910 )  ;
assign n1328 =  ( n39 ) & ( n880 )  ;
assign n1329 =  ( n39 ) & ( n882 )  ;
assign n1330 =  ( n39 ) & ( n884 )  ;
assign n1331 =  ( n39 ) & ( n886 )  ;
assign n1332 =  ( n39 ) & ( n888 )  ;
assign n1333 =  ( n39 ) & ( n890 )  ;
assign n1334 =  ( n39 ) & ( n892 )  ;
assign n1335 =  ( n39 ) & ( n894 )  ;
assign n1336 =  ( n39 ) & ( n896 )  ;
assign n1337 =  ( n39 ) & ( n898 )  ;
assign n1338 =  ( n39 ) & ( n900 )  ;
assign n1339 =  ( n39 ) & ( n902 )  ;
assign n1340 =  ( n39 ) & ( n904 )  ;
assign n1341 =  ( n39 ) & ( n906 )  ;
assign n1342 =  ( n39 ) & ( n908 )  ;
assign n1343 =  ( n39 ) & ( n910 )  ;
assign n1344 =  ( n40 ) & ( n880 )  ;
assign n1345 =  ( n40 ) & ( n882 )  ;
assign n1346 =  ( n40 ) & ( n884 )  ;
assign n1347 =  ( n40 ) & ( n886 )  ;
assign n1348 =  ( n40 ) & ( n888 )  ;
assign n1349 =  ( n40 ) & ( n890 )  ;
assign n1350 =  ( n40 ) & ( n892 )  ;
assign n1351 =  ( n40 ) & ( n894 )  ;
assign n1352 =  ( n40 ) & ( n896 )  ;
assign n1353 =  ( n40 ) & ( n898 )  ;
assign n1354 =  ( n40 ) & ( n900 )  ;
assign n1355 =  ( n40 ) & ( n902 )  ;
assign n1356 =  ( n40 ) & ( n904 )  ;
assign n1357 =  ( n40 ) & ( n906 )  ;
assign n1358 =  ( n40 ) & ( n908 )  ;
assign n1359 =  ( n40 ) & ( n910 )  ;
assign n1360 =  ( n41 ) & ( n880 )  ;
assign n1361 =  ( n41 ) & ( n882 )  ;
assign n1362 =  ( n41 ) & ( n884 )  ;
assign n1363 =  ( n41 ) & ( n886 )  ;
assign n1364 =  ( n41 ) & ( n888 )  ;
assign n1365 =  ( n41 ) & ( n890 )  ;
assign n1366 =  ( n41 ) & ( n892 )  ;
assign n1367 =  ( n41 ) & ( n894 )  ;
assign n1368 =  ( n41 ) & ( n896 )  ;
assign n1369 =  ( n41 ) & ( n898 )  ;
assign n1370 =  ( n41 ) & ( n900 )  ;
assign n1371 =  ( n41 ) & ( n902 )  ;
assign n1372 =  ( n41 ) & ( n904 )  ;
assign n1373 =  ( n41 ) & ( n906 )  ;
assign n1374 =  ( n41 ) & ( n908 )  ;
assign n1375 =  ( n41 ) & ( n910 )  ;
assign n1376 =  ( n42 ) & ( n880 )  ;
assign n1377 =  ( n42 ) & ( n882 )  ;
assign n1378 =  ( n42 ) & ( n884 )  ;
assign n1379 =  ( n42 ) & ( n886 )  ;
assign n1380 =  ( n42 ) & ( n888 )  ;
assign n1381 =  ( n42 ) & ( n890 )  ;
assign n1382 =  ( n42 ) & ( n892 )  ;
assign n1383 =  ( n42 ) & ( n894 )  ;
assign n1384 =  ( n42 ) & ( n896 )  ;
assign n1385 =  ( n42 ) & ( n898 )  ;
assign n1386 =  ( n42 ) & ( n900 )  ;
assign n1387 =  ( n42 ) & ( n902 )  ;
assign n1388 =  ( n42 ) & ( n904 )  ;
assign n1389 =  ( n42 ) & ( n906 )  ;
assign n1390 =  ( n42 ) & ( n908 )  ;
assign n1391 =  ( n42 ) & ( n910 )  ;
assign n1392 =  ( n43 ) & ( n880 )  ;
assign n1393 =  ( n43 ) & ( n882 )  ;
assign n1394 =  ( n43 ) & ( n884 )  ;
assign n1395 =  ( n43 ) & ( n886 )  ;
assign n1396 =  ( n43 ) & ( n888 )  ;
assign n1397 =  ( n43 ) & ( n890 )  ;
assign n1398 =  ( n43 ) & ( n892 )  ;
assign n1399 =  ( n43 ) & ( n894 )  ;
assign n1400 =  ( n43 ) & ( n896 )  ;
assign n1401 =  ( n43 ) & ( n898 )  ;
assign n1402 =  ( n43 ) & ( n900 )  ;
assign n1403 =  ( n43 ) & ( n902 )  ;
assign n1404 =  ( n43 ) & ( n904 )  ;
assign n1405 =  ( n43 ) & ( n906 )  ;
assign n1406 =  ( n43 ) & ( n908 )  ;
assign n1407 =  ( n43 ) & ( n910 )  ;
assign n1408 =  ( n1407 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n1409 =  ( n1406 ) ? ( VREG_0_1 ) : ( n1408 ) ;
assign n1410 =  ( n1405 ) ? ( VREG_0_2 ) : ( n1409 ) ;
assign n1411 =  ( n1404 ) ? ( VREG_0_3 ) : ( n1410 ) ;
assign n1412 =  ( n1403 ) ? ( VREG_0_4 ) : ( n1411 ) ;
assign n1413 =  ( n1402 ) ? ( VREG_0_5 ) : ( n1412 ) ;
assign n1414 =  ( n1401 ) ? ( VREG_0_6 ) : ( n1413 ) ;
assign n1415 =  ( n1400 ) ? ( VREG_0_7 ) : ( n1414 ) ;
assign n1416 =  ( n1399 ) ? ( VREG_0_8 ) : ( n1415 ) ;
assign n1417 =  ( n1398 ) ? ( VREG_0_9 ) : ( n1416 ) ;
assign n1418 =  ( n1397 ) ? ( VREG_0_10 ) : ( n1417 ) ;
assign n1419 =  ( n1396 ) ? ( VREG_0_11 ) : ( n1418 ) ;
assign n1420 =  ( n1395 ) ? ( VREG_0_12 ) : ( n1419 ) ;
assign n1421 =  ( n1394 ) ? ( VREG_0_13 ) : ( n1420 ) ;
assign n1422 =  ( n1393 ) ? ( VREG_0_14 ) : ( n1421 ) ;
assign n1423 =  ( n1392 ) ? ( VREG_0_15 ) : ( n1422 ) ;
assign n1424 =  ( n1391 ) ? ( VREG_1_0 ) : ( n1423 ) ;
assign n1425 =  ( n1390 ) ? ( VREG_1_1 ) : ( n1424 ) ;
assign n1426 =  ( n1389 ) ? ( VREG_1_2 ) : ( n1425 ) ;
assign n1427 =  ( n1388 ) ? ( VREG_1_3 ) : ( n1426 ) ;
assign n1428 =  ( n1387 ) ? ( VREG_1_4 ) : ( n1427 ) ;
assign n1429 =  ( n1386 ) ? ( VREG_1_5 ) : ( n1428 ) ;
assign n1430 =  ( n1385 ) ? ( VREG_1_6 ) : ( n1429 ) ;
assign n1431 =  ( n1384 ) ? ( VREG_1_7 ) : ( n1430 ) ;
assign n1432 =  ( n1383 ) ? ( VREG_1_8 ) : ( n1431 ) ;
assign n1433 =  ( n1382 ) ? ( VREG_1_9 ) : ( n1432 ) ;
assign n1434 =  ( n1381 ) ? ( VREG_1_10 ) : ( n1433 ) ;
assign n1435 =  ( n1380 ) ? ( VREG_1_11 ) : ( n1434 ) ;
assign n1436 =  ( n1379 ) ? ( VREG_1_12 ) : ( n1435 ) ;
assign n1437 =  ( n1378 ) ? ( VREG_1_13 ) : ( n1436 ) ;
assign n1438 =  ( n1377 ) ? ( VREG_1_14 ) : ( n1437 ) ;
assign n1439 =  ( n1376 ) ? ( VREG_1_15 ) : ( n1438 ) ;
assign n1440 =  ( n1375 ) ? ( VREG_2_0 ) : ( n1439 ) ;
assign n1441 =  ( n1374 ) ? ( VREG_2_1 ) : ( n1440 ) ;
assign n1442 =  ( n1373 ) ? ( VREG_2_2 ) : ( n1441 ) ;
assign n1443 =  ( n1372 ) ? ( VREG_2_3 ) : ( n1442 ) ;
assign n1444 =  ( n1371 ) ? ( VREG_2_4 ) : ( n1443 ) ;
assign n1445 =  ( n1370 ) ? ( VREG_2_5 ) : ( n1444 ) ;
assign n1446 =  ( n1369 ) ? ( VREG_2_6 ) : ( n1445 ) ;
assign n1447 =  ( n1368 ) ? ( VREG_2_7 ) : ( n1446 ) ;
assign n1448 =  ( n1367 ) ? ( VREG_2_8 ) : ( n1447 ) ;
assign n1449 =  ( n1366 ) ? ( VREG_2_9 ) : ( n1448 ) ;
assign n1450 =  ( n1365 ) ? ( VREG_2_10 ) : ( n1449 ) ;
assign n1451 =  ( n1364 ) ? ( VREG_2_11 ) : ( n1450 ) ;
assign n1452 =  ( n1363 ) ? ( VREG_2_12 ) : ( n1451 ) ;
assign n1453 =  ( n1362 ) ? ( VREG_2_13 ) : ( n1452 ) ;
assign n1454 =  ( n1361 ) ? ( VREG_2_14 ) : ( n1453 ) ;
assign n1455 =  ( n1360 ) ? ( VREG_2_15 ) : ( n1454 ) ;
assign n1456 =  ( n1359 ) ? ( VREG_3_0 ) : ( n1455 ) ;
assign n1457 =  ( n1358 ) ? ( VREG_3_1 ) : ( n1456 ) ;
assign n1458 =  ( n1357 ) ? ( VREG_3_2 ) : ( n1457 ) ;
assign n1459 =  ( n1356 ) ? ( VREG_3_3 ) : ( n1458 ) ;
assign n1460 =  ( n1355 ) ? ( VREG_3_4 ) : ( n1459 ) ;
assign n1461 =  ( n1354 ) ? ( VREG_3_5 ) : ( n1460 ) ;
assign n1462 =  ( n1353 ) ? ( VREG_3_6 ) : ( n1461 ) ;
assign n1463 =  ( n1352 ) ? ( VREG_3_7 ) : ( n1462 ) ;
assign n1464 =  ( n1351 ) ? ( VREG_3_8 ) : ( n1463 ) ;
assign n1465 =  ( n1350 ) ? ( VREG_3_9 ) : ( n1464 ) ;
assign n1466 =  ( n1349 ) ? ( VREG_3_10 ) : ( n1465 ) ;
assign n1467 =  ( n1348 ) ? ( VREG_3_11 ) : ( n1466 ) ;
assign n1468 =  ( n1347 ) ? ( VREG_3_12 ) : ( n1467 ) ;
assign n1469 =  ( n1346 ) ? ( VREG_3_13 ) : ( n1468 ) ;
assign n1470 =  ( n1345 ) ? ( VREG_3_14 ) : ( n1469 ) ;
assign n1471 =  ( n1344 ) ? ( VREG_3_15 ) : ( n1470 ) ;
assign n1472 =  ( n1343 ) ? ( VREG_4_0 ) : ( n1471 ) ;
assign n1473 =  ( n1342 ) ? ( VREG_4_1 ) : ( n1472 ) ;
assign n1474 =  ( n1341 ) ? ( VREG_4_2 ) : ( n1473 ) ;
assign n1475 =  ( n1340 ) ? ( VREG_4_3 ) : ( n1474 ) ;
assign n1476 =  ( n1339 ) ? ( VREG_4_4 ) : ( n1475 ) ;
assign n1477 =  ( n1338 ) ? ( VREG_4_5 ) : ( n1476 ) ;
assign n1478 =  ( n1337 ) ? ( VREG_4_6 ) : ( n1477 ) ;
assign n1479 =  ( n1336 ) ? ( VREG_4_7 ) : ( n1478 ) ;
assign n1480 =  ( n1335 ) ? ( VREG_4_8 ) : ( n1479 ) ;
assign n1481 =  ( n1334 ) ? ( VREG_4_9 ) : ( n1480 ) ;
assign n1482 =  ( n1333 ) ? ( VREG_4_10 ) : ( n1481 ) ;
assign n1483 =  ( n1332 ) ? ( VREG_4_11 ) : ( n1482 ) ;
assign n1484 =  ( n1331 ) ? ( VREG_4_12 ) : ( n1483 ) ;
assign n1485 =  ( n1330 ) ? ( VREG_4_13 ) : ( n1484 ) ;
assign n1486 =  ( n1329 ) ? ( VREG_4_14 ) : ( n1485 ) ;
assign n1487 =  ( n1328 ) ? ( VREG_4_15 ) : ( n1486 ) ;
assign n1488 =  ( n1327 ) ? ( VREG_5_0 ) : ( n1487 ) ;
assign n1489 =  ( n1326 ) ? ( VREG_5_1 ) : ( n1488 ) ;
assign n1490 =  ( n1325 ) ? ( VREG_5_2 ) : ( n1489 ) ;
assign n1491 =  ( n1324 ) ? ( VREG_5_3 ) : ( n1490 ) ;
assign n1492 =  ( n1323 ) ? ( VREG_5_4 ) : ( n1491 ) ;
assign n1493 =  ( n1322 ) ? ( VREG_5_5 ) : ( n1492 ) ;
assign n1494 =  ( n1321 ) ? ( VREG_5_6 ) : ( n1493 ) ;
assign n1495 =  ( n1320 ) ? ( VREG_5_7 ) : ( n1494 ) ;
assign n1496 =  ( n1319 ) ? ( VREG_5_8 ) : ( n1495 ) ;
assign n1497 =  ( n1318 ) ? ( VREG_5_9 ) : ( n1496 ) ;
assign n1498 =  ( n1317 ) ? ( VREG_5_10 ) : ( n1497 ) ;
assign n1499 =  ( n1316 ) ? ( VREG_5_11 ) : ( n1498 ) ;
assign n1500 =  ( n1315 ) ? ( VREG_5_12 ) : ( n1499 ) ;
assign n1501 =  ( n1314 ) ? ( VREG_5_13 ) : ( n1500 ) ;
assign n1502 =  ( n1313 ) ? ( VREG_5_14 ) : ( n1501 ) ;
assign n1503 =  ( n1312 ) ? ( VREG_5_15 ) : ( n1502 ) ;
assign n1504 =  ( n1311 ) ? ( VREG_6_0 ) : ( n1503 ) ;
assign n1505 =  ( n1310 ) ? ( VREG_6_1 ) : ( n1504 ) ;
assign n1506 =  ( n1309 ) ? ( VREG_6_2 ) : ( n1505 ) ;
assign n1507 =  ( n1308 ) ? ( VREG_6_3 ) : ( n1506 ) ;
assign n1508 =  ( n1307 ) ? ( VREG_6_4 ) : ( n1507 ) ;
assign n1509 =  ( n1306 ) ? ( VREG_6_5 ) : ( n1508 ) ;
assign n1510 =  ( n1305 ) ? ( VREG_6_6 ) : ( n1509 ) ;
assign n1511 =  ( n1304 ) ? ( VREG_6_7 ) : ( n1510 ) ;
assign n1512 =  ( n1303 ) ? ( VREG_6_8 ) : ( n1511 ) ;
assign n1513 =  ( n1302 ) ? ( VREG_6_9 ) : ( n1512 ) ;
assign n1514 =  ( n1301 ) ? ( VREG_6_10 ) : ( n1513 ) ;
assign n1515 =  ( n1300 ) ? ( VREG_6_11 ) : ( n1514 ) ;
assign n1516 =  ( n1299 ) ? ( VREG_6_12 ) : ( n1515 ) ;
assign n1517 =  ( n1298 ) ? ( VREG_6_13 ) : ( n1516 ) ;
assign n1518 =  ( n1297 ) ? ( VREG_6_14 ) : ( n1517 ) ;
assign n1519 =  ( n1296 ) ? ( VREG_6_15 ) : ( n1518 ) ;
assign n1520 =  ( n1295 ) ? ( VREG_7_0 ) : ( n1519 ) ;
assign n1521 =  ( n1294 ) ? ( VREG_7_1 ) : ( n1520 ) ;
assign n1522 =  ( n1293 ) ? ( VREG_7_2 ) : ( n1521 ) ;
assign n1523 =  ( n1292 ) ? ( VREG_7_3 ) : ( n1522 ) ;
assign n1524 =  ( n1291 ) ? ( VREG_7_4 ) : ( n1523 ) ;
assign n1525 =  ( n1290 ) ? ( VREG_7_5 ) : ( n1524 ) ;
assign n1526 =  ( n1289 ) ? ( VREG_7_6 ) : ( n1525 ) ;
assign n1527 =  ( n1288 ) ? ( VREG_7_7 ) : ( n1526 ) ;
assign n1528 =  ( n1287 ) ? ( VREG_7_8 ) : ( n1527 ) ;
assign n1529 =  ( n1286 ) ? ( VREG_7_9 ) : ( n1528 ) ;
assign n1530 =  ( n1285 ) ? ( VREG_7_10 ) : ( n1529 ) ;
assign n1531 =  ( n1284 ) ? ( VREG_7_11 ) : ( n1530 ) ;
assign n1532 =  ( n1283 ) ? ( VREG_7_12 ) : ( n1531 ) ;
assign n1533 =  ( n1282 ) ? ( VREG_7_13 ) : ( n1532 ) ;
assign n1534 =  ( n1281 ) ? ( VREG_7_14 ) : ( n1533 ) ;
assign n1535 =  ( n1280 ) ? ( VREG_7_15 ) : ( n1534 ) ;
assign n1536 =  ( n1279 ) ? ( VREG_8_0 ) : ( n1535 ) ;
assign n1537 =  ( n1278 ) ? ( VREG_8_1 ) : ( n1536 ) ;
assign n1538 =  ( n1277 ) ? ( VREG_8_2 ) : ( n1537 ) ;
assign n1539 =  ( n1276 ) ? ( VREG_8_3 ) : ( n1538 ) ;
assign n1540 =  ( n1275 ) ? ( VREG_8_4 ) : ( n1539 ) ;
assign n1541 =  ( n1274 ) ? ( VREG_8_5 ) : ( n1540 ) ;
assign n1542 =  ( n1273 ) ? ( VREG_8_6 ) : ( n1541 ) ;
assign n1543 =  ( n1272 ) ? ( VREG_8_7 ) : ( n1542 ) ;
assign n1544 =  ( n1271 ) ? ( VREG_8_8 ) : ( n1543 ) ;
assign n1545 =  ( n1270 ) ? ( VREG_8_9 ) : ( n1544 ) ;
assign n1546 =  ( n1269 ) ? ( VREG_8_10 ) : ( n1545 ) ;
assign n1547 =  ( n1268 ) ? ( VREG_8_11 ) : ( n1546 ) ;
assign n1548 =  ( n1267 ) ? ( VREG_8_12 ) : ( n1547 ) ;
assign n1549 =  ( n1266 ) ? ( VREG_8_13 ) : ( n1548 ) ;
assign n1550 =  ( n1265 ) ? ( VREG_8_14 ) : ( n1549 ) ;
assign n1551 =  ( n1264 ) ? ( VREG_8_15 ) : ( n1550 ) ;
assign n1552 =  ( n1263 ) ? ( VREG_9_0 ) : ( n1551 ) ;
assign n1553 =  ( n1262 ) ? ( VREG_9_1 ) : ( n1552 ) ;
assign n1554 =  ( n1261 ) ? ( VREG_9_2 ) : ( n1553 ) ;
assign n1555 =  ( n1260 ) ? ( VREG_9_3 ) : ( n1554 ) ;
assign n1556 =  ( n1259 ) ? ( VREG_9_4 ) : ( n1555 ) ;
assign n1557 =  ( n1258 ) ? ( VREG_9_5 ) : ( n1556 ) ;
assign n1558 =  ( n1257 ) ? ( VREG_9_6 ) : ( n1557 ) ;
assign n1559 =  ( n1256 ) ? ( VREG_9_7 ) : ( n1558 ) ;
assign n1560 =  ( n1255 ) ? ( VREG_9_8 ) : ( n1559 ) ;
assign n1561 =  ( n1254 ) ? ( VREG_9_9 ) : ( n1560 ) ;
assign n1562 =  ( n1253 ) ? ( VREG_9_10 ) : ( n1561 ) ;
assign n1563 =  ( n1252 ) ? ( VREG_9_11 ) : ( n1562 ) ;
assign n1564 =  ( n1251 ) ? ( VREG_9_12 ) : ( n1563 ) ;
assign n1565 =  ( n1250 ) ? ( VREG_9_13 ) : ( n1564 ) ;
assign n1566 =  ( n1249 ) ? ( VREG_9_14 ) : ( n1565 ) ;
assign n1567 =  ( n1248 ) ? ( VREG_9_15 ) : ( n1566 ) ;
assign n1568 =  ( n1247 ) ? ( VREG_10_0 ) : ( n1567 ) ;
assign n1569 =  ( n1246 ) ? ( VREG_10_1 ) : ( n1568 ) ;
assign n1570 =  ( n1245 ) ? ( VREG_10_2 ) : ( n1569 ) ;
assign n1571 =  ( n1244 ) ? ( VREG_10_3 ) : ( n1570 ) ;
assign n1572 =  ( n1243 ) ? ( VREG_10_4 ) : ( n1571 ) ;
assign n1573 =  ( n1242 ) ? ( VREG_10_5 ) : ( n1572 ) ;
assign n1574 =  ( n1241 ) ? ( VREG_10_6 ) : ( n1573 ) ;
assign n1575 =  ( n1240 ) ? ( VREG_10_7 ) : ( n1574 ) ;
assign n1576 =  ( n1239 ) ? ( VREG_10_8 ) : ( n1575 ) ;
assign n1577 =  ( n1238 ) ? ( VREG_10_9 ) : ( n1576 ) ;
assign n1578 =  ( n1237 ) ? ( VREG_10_10 ) : ( n1577 ) ;
assign n1579 =  ( n1236 ) ? ( VREG_10_11 ) : ( n1578 ) ;
assign n1580 =  ( n1235 ) ? ( VREG_10_12 ) : ( n1579 ) ;
assign n1581 =  ( n1234 ) ? ( VREG_10_13 ) : ( n1580 ) ;
assign n1582 =  ( n1233 ) ? ( VREG_10_14 ) : ( n1581 ) ;
assign n1583 =  ( n1232 ) ? ( VREG_10_15 ) : ( n1582 ) ;
assign n1584 =  ( n1231 ) ? ( VREG_11_0 ) : ( n1583 ) ;
assign n1585 =  ( n1230 ) ? ( VREG_11_1 ) : ( n1584 ) ;
assign n1586 =  ( n1229 ) ? ( VREG_11_2 ) : ( n1585 ) ;
assign n1587 =  ( n1228 ) ? ( VREG_11_3 ) : ( n1586 ) ;
assign n1588 =  ( n1227 ) ? ( VREG_11_4 ) : ( n1587 ) ;
assign n1589 =  ( n1226 ) ? ( VREG_11_5 ) : ( n1588 ) ;
assign n1590 =  ( n1225 ) ? ( VREG_11_6 ) : ( n1589 ) ;
assign n1591 =  ( n1224 ) ? ( VREG_11_7 ) : ( n1590 ) ;
assign n1592 =  ( n1223 ) ? ( VREG_11_8 ) : ( n1591 ) ;
assign n1593 =  ( n1222 ) ? ( VREG_11_9 ) : ( n1592 ) ;
assign n1594 =  ( n1221 ) ? ( VREG_11_10 ) : ( n1593 ) ;
assign n1595 =  ( n1220 ) ? ( VREG_11_11 ) : ( n1594 ) ;
assign n1596 =  ( n1219 ) ? ( VREG_11_12 ) : ( n1595 ) ;
assign n1597 =  ( n1218 ) ? ( VREG_11_13 ) : ( n1596 ) ;
assign n1598 =  ( n1217 ) ? ( VREG_11_14 ) : ( n1597 ) ;
assign n1599 =  ( n1216 ) ? ( VREG_11_15 ) : ( n1598 ) ;
assign n1600 =  ( n1215 ) ? ( VREG_12_0 ) : ( n1599 ) ;
assign n1601 =  ( n1214 ) ? ( VREG_12_1 ) : ( n1600 ) ;
assign n1602 =  ( n1213 ) ? ( VREG_12_2 ) : ( n1601 ) ;
assign n1603 =  ( n1212 ) ? ( VREG_12_3 ) : ( n1602 ) ;
assign n1604 =  ( n1211 ) ? ( VREG_12_4 ) : ( n1603 ) ;
assign n1605 =  ( n1210 ) ? ( VREG_12_5 ) : ( n1604 ) ;
assign n1606 =  ( n1209 ) ? ( VREG_12_6 ) : ( n1605 ) ;
assign n1607 =  ( n1208 ) ? ( VREG_12_7 ) : ( n1606 ) ;
assign n1608 =  ( n1207 ) ? ( VREG_12_8 ) : ( n1607 ) ;
assign n1609 =  ( n1206 ) ? ( VREG_12_9 ) : ( n1608 ) ;
assign n1610 =  ( n1205 ) ? ( VREG_12_10 ) : ( n1609 ) ;
assign n1611 =  ( n1204 ) ? ( VREG_12_11 ) : ( n1610 ) ;
assign n1612 =  ( n1203 ) ? ( VREG_12_12 ) : ( n1611 ) ;
assign n1613 =  ( n1202 ) ? ( VREG_12_13 ) : ( n1612 ) ;
assign n1614 =  ( n1201 ) ? ( VREG_12_14 ) : ( n1613 ) ;
assign n1615 =  ( n1200 ) ? ( VREG_12_15 ) : ( n1614 ) ;
assign n1616 =  ( n1199 ) ? ( VREG_13_0 ) : ( n1615 ) ;
assign n1617 =  ( n1198 ) ? ( VREG_13_1 ) : ( n1616 ) ;
assign n1618 =  ( n1197 ) ? ( VREG_13_2 ) : ( n1617 ) ;
assign n1619 =  ( n1196 ) ? ( VREG_13_3 ) : ( n1618 ) ;
assign n1620 =  ( n1195 ) ? ( VREG_13_4 ) : ( n1619 ) ;
assign n1621 =  ( n1194 ) ? ( VREG_13_5 ) : ( n1620 ) ;
assign n1622 =  ( n1193 ) ? ( VREG_13_6 ) : ( n1621 ) ;
assign n1623 =  ( n1192 ) ? ( VREG_13_7 ) : ( n1622 ) ;
assign n1624 =  ( n1191 ) ? ( VREG_13_8 ) : ( n1623 ) ;
assign n1625 =  ( n1190 ) ? ( VREG_13_9 ) : ( n1624 ) ;
assign n1626 =  ( n1189 ) ? ( VREG_13_10 ) : ( n1625 ) ;
assign n1627 =  ( n1188 ) ? ( VREG_13_11 ) : ( n1626 ) ;
assign n1628 =  ( n1187 ) ? ( VREG_13_12 ) : ( n1627 ) ;
assign n1629 =  ( n1186 ) ? ( VREG_13_13 ) : ( n1628 ) ;
assign n1630 =  ( n1185 ) ? ( VREG_13_14 ) : ( n1629 ) ;
assign n1631 =  ( n1184 ) ? ( VREG_13_15 ) : ( n1630 ) ;
assign n1632 =  ( n1183 ) ? ( VREG_14_0 ) : ( n1631 ) ;
assign n1633 =  ( n1182 ) ? ( VREG_14_1 ) : ( n1632 ) ;
assign n1634 =  ( n1181 ) ? ( VREG_14_2 ) : ( n1633 ) ;
assign n1635 =  ( n1180 ) ? ( VREG_14_3 ) : ( n1634 ) ;
assign n1636 =  ( n1179 ) ? ( VREG_14_4 ) : ( n1635 ) ;
assign n1637 =  ( n1178 ) ? ( VREG_14_5 ) : ( n1636 ) ;
assign n1638 =  ( n1177 ) ? ( VREG_14_6 ) : ( n1637 ) ;
assign n1639 =  ( n1176 ) ? ( VREG_14_7 ) : ( n1638 ) ;
assign n1640 =  ( n1175 ) ? ( VREG_14_8 ) : ( n1639 ) ;
assign n1641 =  ( n1174 ) ? ( VREG_14_9 ) : ( n1640 ) ;
assign n1642 =  ( n1173 ) ? ( VREG_14_10 ) : ( n1641 ) ;
assign n1643 =  ( n1172 ) ? ( VREG_14_11 ) : ( n1642 ) ;
assign n1644 =  ( n1171 ) ? ( VREG_14_12 ) : ( n1643 ) ;
assign n1645 =  ( n1170 ) ? ( VREG_14_13 ) : ( n1644 ) ;
assign n1646 =  ( n1169 ) ? ( VREG_14_14 ) : ( n1645 ) ;
assign n1647 =  ( n1168 ) ? ( VREG_14_15 ) : ( n1646 ) ;
assign n1648 =  ( n1167 ) ? ( VREG_15_0 ) : ( n1647 ) ;
assign n1649 =  ( n1166 ) ? ( VREG_15_1 ) : ( n1648 ) ;
assign n1650 =  ( n1165 ) ? ( VREG_15_2 ) : ( n1649 ) ;
assign n1651 =  ( n1164 ) ? ( VREG_15_3 ) : ( n1650 ) ;
assign n1652 =  ( n1163 ) ? ( VREG_15_4 ) : ( n1651 ) ;
assign n1653 =  ( n1162 ) ? ( VREG_15_5 ) : ( n1652 ) ;
assign n1654 =  ( n1161 ) ? ( VREG_15_6 ) : ( n1653 ) ;
assign n1655 =  ( n1160 ) ? ( VREG_15_7 ) : ( n1654 ) ;
assign n1656 =  ( n1159 ) ? ( VREG_15_8 ) : ( n1655 ) ;
assign n1657 =  ( n1158 ) ? ( VREG_15_9 ) : ( n1656 ) ;
assign n1658 =  ( n1157 ) ? ( VREG_15_10 ) : ( n1657 ) ;
assign n1659 =  ( n1156 ) ? ( VREG_15_11 ) : ( n1658 ) ;
assign n1660 =  ( n1155 ) ? ( VREG_15_12 ) : ( n1659 ) ;
assign n1661 =  ( n1154 ) ? ( VREG_15_13 ) : ( n1660 ) ;
assign n1662 =  ( n1153 ) ? ( VREG_15_14 ) : ( n1661 ) ;
assign n1663 =  ( n1152 ) ? ( VREG_15_15 ) : ( n1662 ) ;
assign n1664 =  ( n1151 ) ? ( VREG_16_0 ) : ( n1663 ) ;
assign n1665 =  ( n1150 ) ? ( VREG_16_1 ) : ( n1664 ) ;
assign n1666 =  ( n1149 ) ? ( VREG_16_2 ) : ( n1665 ) ;
assign n1667 =  ( n1148 ) ? ( VREG_16_3 ) : ( n1666 ) ;
assign n1668 =  ( n1147 ) ? ( VREG_16_4 ) : ( n1667 ) ;
assign n1669 =  ( n1146 ) ? ( VREG_16_5 ) : ( n1668 ) ;
assign n1670 =  ( n1145 ) ? ( VREG_16_6 ) : ( n1669 ) ;
assign n1671 =  ( n1144 ) ? ( VREG_16_7 ) : ( n1670 ) ;
assign n1672 =  ( n1143 ) ? ( VREG_16_8 ) : ( n1671 ) ;
assign n1673 =  ( n1142 ) ? ( VREG_16_9 ) : ( n1672 ) ;
assign n1674 =  ( n1141 ) ? ( VREG_16_10 ) : ( n1673 ) ;
assign n1675 =  ( n1140 ) ? ( VREG_16_11 ) : ( n1674 ) ;
assign n1676 =  ( n1139 ) ? ( VREG_16_12 ) : ( n1675 ) ;
assign n1677 =  ( n1138 ) ? ( VREG_16_13 ) : ( n1676 ) ;
assign n1678 =  ( n1137 ) ? ( VREG_16_14 ) : ( n1677 ) ;
assign n1679 =  ( n1136 ) ? ( VREG_16_15 ) : ( n1678 ) ;
assign n1680 =  ( n1135 ) ? ( VREG_17_0 ) : ( n1679 ) ;
assign n1681 =  ( n1134 ) ? ( VREG_17_1 ) : ( n1680 ) ;
assign n1682 =  ( n1133 ) ? ( VREG_17_2 ) : ( n1681 ) ;
assign n1683 =  ( n1132 ) ? ( VREG_17_3 ) : ( n1682 ) ;
assign n1684 =  ( n1131 ) ? ( VREG_17_4 ) : ( n1683 ) ;
assign n1685 =  ( n1130 ) ? ( VREG_17_5 ) : ( n1684 ) ;
assign n1686 =  ( n1129 ) ? ( VREG_17_6 ) : ( n1685 ) ;
assign n1687 =  ( n1128 ) ? ( VREG_17_7 ) : ( n1686 ) ;
assign n1688 =  ( n1127 ) ? ( VREG_17_8 ) : ( n1687 ) ;
assign n1689 =  ( n1126 ) ? ( VREG_17_9 ) : ( n1688 ) ;
assign n1690 =  ( n1125 ) ? ( VREG_17_10 ) : ( n1689 ) ;
assign n1691 =  ( n1124 ) ? ( VREG_17_11 ) : ( n1690 ) ;
assign n1692 =  ( n1123 ) ? ( VREG_17_12 ) : ( n1691 ) ;
assign n1693 =  ( n1122 ) ? ( VREG_17_13 ) : ( n1692 ) ;
assign n1694 =  ( n1121 ) ? ( VREG_17_14 ) : ( n1693 ) ;
assign n1695 =  ( n1120 ) ? ( VREG_17_15 ) : ( n1694 ) ;
assign n1696 =  ( n1119 ) ? ( VREG_18_0 ) : ( n1695 ) ;
assign n1697 =  ( n1118 ) ? ( VREG_18_1 ) : ( n1696 ) ;
assign n1698 =  ( n1117 ) ? ( VREG_18_2 ) : ( n1697 ) ;
assign n1699 =  ( n1116 ) ? ( VREG_18_3 ) : ( n1698 ) ;
assign n1700 =  ( n1115 ) ? ( VREG_18_4 ) : ( n1699 ) ;
assign n1701 =  ( n1114 ) ? ( VREG_18_5 ) : ( n1700 ) ;
assign n1702 =  ( n1113 ) ? ( VREG_18_6 ) : ( n1701 ) ;
assign n1703 =  ( n1112 ) ? ( VREG_18_7 ) : ( n1702 ) ;
assign n1704 =  ( n1111 ) ? ( VREG_18_8 ) : ( n1703 ) ;
assign n1705 =  ( n1110 ) ? ( VREG_18_9 ) : ( n1704 ) ;
assign n1706 =  ( n1109 ) ? ( VREG_18_10 ) : ( n1705 ) ;
assign n1707 =  ( n1108 ) ? ( VREG_18_11 ) : ( n1706 ) ;
assign n1708 =  ( n1107 ) ? ( VREG_18_12 ) : ( n1707 ) ;
assign n1709 =  ( n1106 ) ? ( VREG_18_13 ) : ( n1708 ) ;
assign n1710 =  ( n1105 ) ? ( VREG_18_14 ) : ( n1709 ) ;
assign n1711 =  ( n1104 ) ? ( VREG_18_15 ) : ( n1710 ) ;
assign n1712 =  ( n1103 ) ? ( VREG_19_0 ) : ( n1711 ) ;
assign n1713 =  ( n1102 ) ? ( VREG_19_1 ) : ( n1712 ) ;
assign n1714 =  ( n1101 ) ? ( VREG_19_2 ) : ( n1713 ) ;
assign n1715 =  ( n1100 ) ? ( VREG_19_3 ) : ( n1714 ) ;
assign n1716 =  ( n1099 ) ? ( VREG_19_4 ) : ( n1715 ) ;
assign n1717 =  ( n1098 ) ? ( VREG_19_5 ) : ( n1716 ) ;
assign n1718 =  ( n1097 ) ? ( VREG_19_6 ) : ( n1717 ) ;
assign n1719 =  ( n1096 ) ? ( VREG_19_7 ) : ( n1718 ) ;
assign n1720 =  ( n1095 ) ? ( VREG_19_8 ) : ( n1719 ) ;
assign n1721 =  ( n1094 ) ? ( VREG_19_9 ) : ( n1720 ) ;
assign n1722 =  ( n1093 ) ? ( VREG_19_10 ) : ( n1721 ) ;
assign n1723 =  ( n1092 ) ? ( VREG_19_11 ) : ( n1722 ) ;
assign n1724 =  ( n1091 ) ? ( VREG_19_12 ) : ( n1723 ) ;
assign n1725 =  ( n1090 ) ? ( VREG_19_13 ) : ( n1724 ) ;
assign n1726 =  ( n1089 ) ? ( VREG_19_14 ) : ( n1725 ) ;
assign n1727 =  ( n1088 ) ? ( VREG_19_15 ) : ( n1726 ) ;
assign n1728 =  ( n1087 ) ? ( VREG_20_0 ) : ( n1727 ) ;
assign n1729 =  ( n1086 ) ? ( VREG_20_1 ) : ( n1728 ) ;
assign n1730 =  ( n1085 ) ? ( VREG_20_2 ) : ( n1729 ) ;
assign n1731 =  ( n1084 ) ? ( VREG_20_3 ) : ( n1730 ) ;
assign n1732 =  ( n1083 ) ? ( VREG_20_4 ) : ( n1731 ) ;
assign n1733 =  ( n1082 ) ? ( VREG_20_5 ) : ( n1732 ) ;
assign n1734 =  ( n1081 ) ? ( VREG_20_6 ) : ( n1733 ) ;
assign n1735 =  ( n1080 ) ? ( VREG_20_7 ) : ( n1734 ) ;
assign n1736 =  ( n1079 ) ? ( VREG_20_8 ) : ( n1735 ) ;
assign n1737 =  ( n1078 ) ? ( VREG_20_9 ) : ( n1736 ) ;
assign n1738 =  ( n1077 ) ? ( VREG_20_10 ) : ( n1737 ) ;
assign n1739 =  ( n1076 ) ? ( VREG_20_11 ) : ( n1738 ) ;
assign n1740 =  ( n1075 ) ? ( VREG_20_12 ) : ( n1739 ) ;
assign n1741 =  ( n1074 ) ? ( VREG_20_13 ) : ( n1740 ) ;
assign n1742 =  ( n1073 ) ? ( VREG_20_14 ) : ( n1741 ) ;
assign n1743 =  ( n1072 ) ? ( VREG_20_15 ) : ( n1742 ) ;
assign n1744 =  ( n1071 ) ? ( VREG_21_0 ) : ( n1743 ) ;
assign n1745 =  ( n1070 ) ? ( VREG_21_1 ) : ( n1744 ) ;
assign n1746 =  ( n1069 ) ? ( VREG_21_2 ) : ( n1745 ) ;
assign n1747 =  ( n1068 ) ? ( VREG_21_3 ) : ( n1746 ) ;
assign n1748 =  ( n1067 ) ? ( VREG_21_4 ) : ( n1747 ) ;
assign n1749 =  ( n1066 ) ? ( VREG_21_5 ) : ( n1748 ) ;
assign n1750 =  ( n1065 ) ? ( VREG_21_6 ) : ( n1749 ) ;
assign n1751 =  ( n1064 ) ? ( VREG_21_7 ) : ( n1750 ) ;
assign n1752 =  ( n1063 ) ? ( VREG_21_8 ) : ( n1751 ) ;
assign n1753 =  ( n1062 ) ? ( VREG_21_9 ) : ( n1752 ) ;
assign n1754 =  ( n1061 ) ? ( VREG_21_10 ) : ( n1753 ) ;
assign n1755 =  ( n1060 ) ? ( VREG_21_11 ) : ( n1754 ) ;
assign n1756 =  ( n1059 ) ? ( VREG_21_12 ) : ( n1755 ) ;
assign n1757 =  ( n1058 ) ? ( VREG_21_13 ) : ( n1756 ) ;
assign n1758 =  ( n1057 ) ? ( VREG_21_14 ) : ( n1757 ) ;
assign n1759 =  ( n1056 ) ? ( VREG_21_15 ) : ( n1758 ) ;
assign n1760 =  ( n1055 ) ? ( VREG_22_0 ) : ( n1759 ) ;
assign n1761 =  ( n1054 ) ? ( VREG_22_1 ) : ( n1760 ) ;
assign n1762 =  ( n1053 ) ? ( VREG_22_2 ) : ( n1761 ) ;
assign n1763 =  ( n1052 ) ? ( VREG_22_3 ) : ( n1762 ) ;
assign n1764 =  ( n1051 ) ? ( VREG_22_4 ) : ( n1763 ) ;
assign n1765 =  ( n1050 ) ? ( VREG_22_5 ) : ( n1764 ) ;
assign n1766 =  ( n1049 ) ? ( VREG_22_6 ) : ( n1765 ) ;
assign n1767 =  ( n1048 ) ? ( VREG_22_7 ) : ( n1766 ) ;
assign n1768 =  ( n1047 ) ? ( VREG_22_8 ) : ( n1767 ) ;
assign n1769 =  ( n1046 ) ? ( VREG_22_9 ) : ( n1768 ) ;
assign n1770 =  ( n1045 ) ? ( VREG_22_10 ) : ( n1769 ) ;
assign n1771 =  ( n1044 ) ? ( VREG_22_11 ) : ( n1770 ) ;
assign n1772 =  ( n1043 ) ? ( VREG_22_12 ) : ( n1771 ) ;
assign n1773 =  ( n1042 ) ? ( VREG_22_13 ) : ( n1772 ) ;
assign n1774 =  ( n1041 ) ? ( VREG_22_14 ) : ( n1773 ) ;
assign n1775 =  ( n1040 ) ? ( VREG_22_15 ) : ( n1774 ) ;
assign n1776 =  ( n1039 ) ? ( VREG_23_0 ) : ( n1775 ) ;
assign n1777 =  ( n1038 ) ? ( VREG_23_1 ) : ( n1776 ) ;
assign n1778 =  ( n1037 ) ? ( VREG_23_2 ) : ( n1777 ) ;
assign n1779 =  ( n1036 ) ? ( VREG_23_3 ) : ( n1778 ) ;
assign n1780 =  ( n1035 ) ? ( VREG_23_4 ) : ( n1779 ) ;
assign n1781 =  ( n1034 ) ? ( VREG_23_5 ) : ( n1780 ) ;
assign n1782 =  ( n1033 ) ? ( VREG_23_6 ) : ( n1781 ) ;
assign n1783 =  ( n1032 ) ? ( VREG_23_7 ) : ( n1782 ) ;
assign n1784 =  ( n1031 ) ? ( VREG_23_8 ) : ( n1783 ) ;
assign n1785 =  ( n1030 ) ? ( VREG_23_9 ) : ( n1784 ) ;
assign n1786 =  ( n1029 ) ? ( VREG_23_10 ) : ( n1785 ) ;
assign n1787 =  ( n1028 ) ? ( VREG_23_11 ) : ( n1786 ) ;
assign n1788 =  ( n1027 ) ? ( VREG_23_12 ) : ( n1787 ) ;
assign n1789 =  ( n1026 ) ? ( VREG_23_13 ) : ( n1788 ) ;
assign n1790 =  ( n1025 ) ? ( VREG_23_14 ) : ( n1789 ) ;
assign n1791 =  ( n1024 ) ? ( VREG_23_15 ) : ( n1790 ) ;
assign n1792 =  ( n1023 ) ? ( VREG_24_0 ) : ( n1791 ) ;
assign n1793 =  ( n1022 ) ? ( VREG_24_1 ) : ( n1792 ) ;
assign n1794 =  ( n1021 ) ? ( VREG_24_2 ) : ( n1793 ) ;
assign n1795 =  ( n1020 ) ? ( VREG_24_3 ) : ( n1794 ) ;
assign n1796 =  ( n1019 ) ? ( VREG_24_4 ) : ( n1795 ) ;
assign n1797 =  ( n1018 ) ? ( VREG_24_5 ) : ( n1796 ) ;
assign n1798 =  ( n1017 ) ? ( VREG_24_6 ) : ( n1797 ) ;
assign n1799 =  ( n1016 ) ? ( VREG_24_7 ) : ( n1798 ) ;
assign n1800 =  ( n1015 ) ? ( VREG_24_8 ) : ( n1799 ) ;
assign n1801 =  ( n1014 ) ? ( VREG_24_9 ) : ( n1800 ) ;
assign n1802 =  ( n1013 ) ? ( VREG_24_10 ) : ( n1801 ) ;
assign n1803 =  ( n1012 ) ? ( VREG_24_11 ) : ( n1802 ) ;
assign n1804 =  ( n1011 ) ? ( VREG_24_12 ) : ( n1803 ) ;
assign n1805 =  ( n1010 ) ? ( VREG_24_13 ) : ( n1804 ) ;
assign n1806 =  ( n1009 ) ? ( VREG_24_14 ) : ( n1805 ) ;
assign n1807 =  ( n1008 ) ? ( VREG_24_15 ) : ( n1806 ) ;
assign n1808 =  ( n1007 ) ? ( VREG_25_0 ) : ( n1807 ) ;
assign n1809 =  ( n1006 ) ? ( VREG_25_1 ) : ( n1808 ) ;
assign n1810 =  ( n1005 ) ? ( VREG_25_2 ) : ( n1809 ) ;
assign n1811 =  ( n1004 ) ? ( VREG_25_3 ) : ( n1810 ) ;
assign n1812 =  ( n1003 ) ? ( VREG_25_4 ) : ( n1811 ) ;
assign n1813 =  ( n1002 ) ? ( VREG_25_5 ) : ( n1812 ) ;
assign n1814 =  ( n1001 ) ? ( VREG_25_6 ) : ( n1813 ) ;
assign n1815 =  ( n1000 ) ? ( VREG_25_7 ) : ( n1814 ) ;
assign n1816 =  ( n999 ) ? ( VREG_25_8 ) : ( n1815 ) ;
assign n1817 =  ( n998 ) ? ( VREG_25_9 ) : ( n1816 ) ;
assign n1818 =  ( n997 ) ? ( VREG_25_10 ) : ( n1817 ) ;
assign n1819 =  ( n996 ) ? ( VREG_25_11 ) : ( n1818 ) ;
assign n1820 =  ( n995 ) ? ( VREG_25_12 ) : ( n1819 ) ;
assign n1821 =  ( n994 ) ? ( VREG_25_13 ) : ( n1820 ) ;
assign n1822 =  ( n993 ) ? ( VREG_25_14 ) : ( n1821 ) ;
assign n1823 =  ( n992 ) ? ( VREG_25_15 ) : ( n1822 ) ;
assign n1824 =  ( n991 ) ? ( VREG_26_0 ) : ( n1823 ) ;
assign n1825 =  ( n990 ) ? ( VREG_26_1 ) : ( n1824 ) ;
assign n1826 =  ( n989 ) ? ( VREG_26_2 ) : ( n1825 ) ;
assign n1827 =  ( n988 ) ? ( VREG_26_3 ) : ( n1826 ) ;
assign n1828 =  ( n987 ) ? ( VREG_26_4 ) : ( n1827 ) ;
assign n1829 =  ( n986 ) ? ( VREG_26_5 ) : ( n1828 ) ;
assign n1830 =  ( n985 ) ? ( VREG_26_6 ) : ( n1829 ) ;
assign n1831 =  ( n984 ) ? ( VREG_26_7 ) : ( n1830 ) ;
assign n1832 =  ( n983 ) ? ( VREG_26_8 ) : ( n1831 ) ;
assign n1833 =  ( n982 ) ? ( VREG_26_9 ) : ( n1832 ) ;
assign n1834 =  ( n981 ) ? ( VREG_26_10 ) : ( n1833 ) ;
assign n1835 =  ( n980 ) ? ( VREG_26_11 ) : ( n1834 ) ;
assign n1836 =  ( n979 ) ? ( VREG_26_12 ) : ( n1835 ) ;
assign n1837 =  ( n978 ) ? ( VREG_26_13 ) : ( n1836 ) ;
assign n1838 =  ( n977 ) ? ( VREG_26_14 ) : ( n1837 ) ;
assign n1839 =  ( n976 ) ? ( VREG_26_15 ) : ( n1838 ) ;
assign n1840 =  ( n975 ) ? ( VREG_27_0 ) : ( n1839 ) ;
assign n1841 =  ( n974 ) ? ( VREG_27_1 ) : ( n1840 ) ;
assign n1842 =  ( n973 ) ? ( VREG_27_2 ) : ( n1841 ) ;
assign n1843 =  ( n972 ) ? ( VREG_27_3 ) : ( n1842 ) ;
assign n1844 =  ( n971 ) ? ( VREG_27_4 ) : ( n1843 ) ;
assign n1845 =  ( n970 ) ? ( VREG_27_5 ) : ( n1844 ) ;
assign n1846 =  ( n969 ) ? ( VREG_27_6 ) : ( n1845 ) ;
assign n1847 =  ( n968 ) ? ( VREG_27_7 ) : ( n1846 ) ;
assign n1848 =  ( n967 ) ? ( VREG_27_8 ) : ( n1847 ) ;
assign n1849 =  ( n966 ) ? ( VREG_27_9 ) : ( n1848 ) ;
assign n1850 =  ( n965 ) ? ( VREG_27_10 ) : ( n1849 ) ;
assign n1851 =  ( n964 ) ? ( VREG_27_11 ) : ( n1850 ) ;
assign n1852 =  ( n963 ) ? ( VREG_27_12 ) : ( n1851 ) ;
assign n1853 =  ( n962 ) ? ( VREG_27_13 ) : ( n1852 ) ;
assign n1854 =  ( n961 ) ? ( VREG_27_14 ) : ( n1853 ) ;
assign n1855 =  ( n960 ) ? ( VREG_27_15 ) : ( n1854 ) ;
assign n1856 =  ( n959 ) ? ( VREG_28_0 ) : ( n1855 ) ;
assign n1857 =  ( n958 ) ? ( VREG_28_1 ) : ( n1856 ) ;
assign n1858 =  ( n957 ) ? ( VREG_28_2 ) : ( n1857 ) ;
assign n1859 =  ( n956 ) ? ( VREG_28_3 ) : ( n1858 ) ;
assign n1860 =  ( n955 ) ? ( VREG_28_4 ) : ( n1859 ) ;
assign n1861 =  ( n954 ) ? ( VREG_28_5 ) : ( n1860 ) ;
assign n1862 =  ( n953 ) ? ( VREG_28_6 ) : ( n1861 ) ;
assign n1863 =  ( n952 ) ? ( VREG_28_7 ) : ( n1862 ) ;
assign n1864 =  ( n951 ) ? ( VREG_28_8 ) : ( n1863 ) ;
assign n1865 =  ( n950 ) ? ( VREG_28_9 ) : ( n1864 ) ;
assign n1866 =  ( n949 ) ? ( VREG_28_10 ) : ( n1865 ) ;
assign n1867 =  ( n948 ) ? ( VREG_28_11 ) : ( n1866 ) ;
assign n1868 =  ( n947 ) ? ( VREG_28_12 ) : ( n1867 ) ;
assign n1869 =  ( n946 ) ? ( VREG_28_13 ) : ( n1868 ) ;
assign n1870 =  ( n945 ) ? ( VREG_28_14 ) : ( n1869 ) ;
assign n1871 =  ( n944 ) ? ( VREG_28_15 ) : ( n1870 ) ;
assign n1872 =  ( n943 ) ? ( VREG_29_0 ) : ( n1871 ) ;
assign n1873 =  ( n942 ) ? ( VREG_29_1 ) : ( n1872 ) ;
assign n1874 =  ( n941 ) ? ( VREG_29_2 ) : ( n1873 ) ;
assign n1875 =  ( n940 ) ? ( VREG_29_3 ) : ( n1874 ) ;
assign n1876 =  ( n939 ) ? ( VREG_29_4 ) : ( n1875 ) ;
assign n1877 =  ( n938 ) ? ( VREG_29_5 ) : ( n1876 ) ;
assign n1878 =  ( n937 ) ? ( VREG_29_6 ) : ( n1877 ) ;
assign n1879 =  ( n936 ) ? ( VREG_29_7 ) : ( n1878 ) ;
assign n1880 =  ( n935 ) ? ( VREG_29_8 ) : ( n1879 ) ;
assign n1881 =  ( n934 ) ? ( VREG_29_9 ) : ( n1880 ) ;
assign n1882 =  ( n933 ) ? ( VREG_29_10 ) : ( n1881 ) ;
assign n1883 =  ( n932 ) ? ( VREG_29_11 ) : ( n1882 ) ;
assign n1884 =  ( n931 ) ? ( VREG_29_12 ) : ( n1883 ) ;
assign n1885 =  ( n930 ) ? ( VREG_29_13 ) : ( n1884 ) ;
assign n1886 =  ( n929 ) ? ( VREG_29_14 ) : ( n1885 ) ;
assign n1887 =  ( n928 ) ? ( VREG_29_15 ) : ( n1886 ) ;
assign n1888 =  ( n927 ) ? ( VREG_30_0 ) : ( n1887 ) ;
assign n1889 =  ( n926 ) ? ( VREG_30_1 ) : ( n1888 ) ;
assign n1890 =  ( n925 ) ? ( VREG_30_2 ) : ( n1889 ) ;
assign n1891 =  ( n924 ) ? ( VREG_30_3 ) : ( n1890 ) ;
assign n1892 =  ( n923 ) ? ( VREG_30_4 ) : ( n1891 ) ;
assign n1893 =  ( n922 ) ? ( VREG_30_5 ) : ( n1892 ) ;
assign n1894 =  ( n921 ) ? ( VREG_30_6 ) : ( n1893 ) ;
assign n1895 =  ( n920 ) ? ( VREG_30_7 ) : ( n1894 ) ;
assign n1896 =  ( n919 ) ? ( VREG_30_8 ) : ( n1895 ) ;
assign n1897 =  ( n918 ) ? ( VREG_30_9 ) : ( n1896 ) ;
assign n1898 =  ( n917 ) ? ( VREG_30_10 ) : ( n1897 ) ;
assign n1899 =  ( n916 ) ? ( VREG_30_11 ) : ( n1898 ) ;
assign n1900 =  ( n915 ) ? ( VREG_30_12 ) : ( n1899 ) ;
assign n1901 =  ( n914 ) ? ( VREG_30_13 ) : ( n1900 ) ;
assign n1902 =  ( n913 ) ? ( VREG_30_14 ) : ( n1901 ) ;
assign n1903 =  ( n912 ) ? ( VREG_30_15 ) : ( n1902 ) ;
assign n1904 =  ( n911 ) ? ( VREG_31_0 ) : ( n1903 ) ;
assign n1905 =  ( n909 ) ? ( VREG_31_1 ) : ( n1904 ) ;
assign n1906 =  ( n907 ) ? ( VREG_31_2 ) : ( n1905 ) ;
assign n1907 =  ( n905 ) ? ( VREG_31_3 ) : ( n1906 ) ;
assign n1908 =  ( n903 ) ? ( VREG_31_4 ) : ( n1907 ) ;
assign n1909 =  ( n901 ) ? ( VREG_31_5 ) : ( n1908 ) ;
assign n1910 =  ( n899 ) ? ( VREG_31_6 ) : ( n1909 ) ;
assign n1911 =  ( n897 ) ? ( VREG_31_7 ) : ( n1910 ) ;
assign n1912 =  ( n895 ) ? ( VREG_31_8 ) : ( n1911 ) ;
assign n1913 =  ( n893 ) ? ( VREG_31_9 ) : ( n1912 ) ;
assign n1914 =  ( n891 ) ? ( VREG_31_10 ) : ( n1913 ) ;
assign n1915 =  ( n889 ) ? ( VREG_31_11 ) : ( n1914 ) ;
assign n1916 =  ( n887 ) ? ( VREG_31_12 ) : ( n1915 ) ;
assign n1917 =  ( n885 ) ? ( VREG_31_13 ) : ( n1916 ) ;
assign n1918 =  ( n883 ) ? ( VREG_31_14 ) : ( n1917 ) ;
assign n1919 =  ( n881 ) ? ( VREG_31_15 ) : ( n1918 ) ;
assign n1920 =  ( n1919 ) + ( n140 )  ;
assign n1921 =  ( n1919 ) - ( n140 )  ;
assign n1922 =  ( n1919 ) & ( n140 )  ;
assign n1923 =  ( n1919 ) | ( n140 )  ;
assign n1924 =  ( ( n1919 ) * ( n140 ))  ;
assign n1925 =  ( n148 ) ? ( n1924 ) : ( VREG_0_0 ) ;
assign n1926 =  ( n146 ) ? ( n1923 ) : ( n1925 ) ;
assign n1927 =  ( n144 ) ? ( n1922 ) : ( n1926 ) ;
assign n1928 =  ( n142 ) ? ( n1921 ) : ( n1927 ) ;
assign n1929 =  ( n10 ) ? ( n1920 ) : ( n1928 ) ;
assign n1930 =  ( n7 ) == ( 3'd4 )  ;
assign n1931 =  ( n77 ) & ( n880 )  ;
assign n1932 =  ( n77 ) & ( n882 )  ;
assign n1933 =  ( n77 ) & ( n884 )  ;
assign n1934 =  ( n77 ) & ( n886 )  ;
assign n1935 =  ( n77 ) & ( n888 )  ;
assign n1936 =  ( n77 ) & ( n890 )  ;
assign n1937 =  ( n77 ) & ( n892 )  ;
assign n1938 =  ( n77 ) & ( n894 )  ;
assign n1939 =  ( n77 ) & ( n896 )  ;
assign n1940 =  ( n77 ) & ( n898 )  ;
assign n1941 =  ( n77 ) & ( n900 )  ;
assign n1942 =  ( n77 ) & ( n902 )  ;
assign n1943 =  ( n77 ) & ( n904 )  ;
assign n1944 =  ( n77 ) & ( n906 )  ;
assign n1945 =  ( n77 ) & ( n908 )  ;
assign n1946 =  ( n77 ) & ( n910 )  ;
assign n1947 =  ( n78 ) & ( n880 )  ;
assign n1948 =  ( n78 ) & ( n882 )  ;
assign n1949 =  ( n78 ) & ( n884 )  ;
assign n1950 =  ( n78 ) & ( n886 )  ;
assign n1951 =  ( n78 ) & ( n888 )  ;
assign n1952 =  ( n78 ) & ( n890 )  ;
assign n1953 =  ( n78 ) & ( n892 )  ;
assign n1954 =  ( n78 ) & ( n894 )  ;
assign n1955 =  ( n78 ) & ( n896 )  ;
assign n1956 =  ( n78 ) & ( n898 )  ;
assign n1957 =  ( n78 ) & ( n900 )  ;
assign n1958 =  ( n78 ) & ( n902 )  ;
assign n1959 =  ( n78 ) & ( n904 )  ;
assign n1960 =  ( n78 ) & ( n906 )  ;
assign n1961 =  ( n78 ) & ( n908 )  ;
assign n1962 =  ( n78 ) & ( n910 )  ;
assign n1963 =  ( n79 ) & ( n880 )  ;
assign n1964 =  ( n79 ) & ( n882 )  ;
assign n1965 =  ( n79 ) & ( n884 )  ;
assign n1966 =  ( n79 ) & ( n886 )  ;
assign n1967 =  ( n79 ) & ( n888 )  ;
assign n1968 =  ( n79 ) & ( n890 )  ;
assign n1969 =  ( n79 ) & ( n892 )  ;
assign n1970 =  ( n79 ) & ( n894 )  ;
assign n1971 =  ( n79 ) & ( n896 )  ;
assign n1972 =  ( n79 ) & ( n898 )  ;
assign n1973 =  ( n79 ) & ( n900 )  ;
assign n1974 =  ( n79 ) & ( n902 )  ;
assign n1975 =  ( n79 ) & ( n904 )  ;
assign n1976 =  ( n79 ) & ( n906 )  ;
assign n1977 =  ( n79 ) & ( n908 )  ;
assign n1978 =  ( n79 ) & ( n910 )  ;
assign n1979 =  ( n80 ) & ( n880 )  ;
assign n1980 =  ( n80 ) & ( n882 )  ;
assign n1981 =  ( n80 ) & ( n884 )  ;
assign n1982 =  ( n80 ) & ( n886 )  ;
assign n1983 =  ( n80 ) & ( n888 )  ;
assign n1984 =  ( n80 ) & ( n890 )  ;
assign n1985 =  ( n80 ) & ( n892 )  ;
assign n1986 =  ( n80 ) & ( n894 )  ;
assign n1987 =  ( n80 ) & ( n896 )  ;
assign n1988 =  ( n80 ) & ( n898 )  ;
assign n1989 =  ( n80 ) & ( n900 )  ;
assign n1990 =  ( n80 ) & ( n902 )  ;
assign n1991 =  ( n80 ) & ( n904 )  ;
assign n1992 =  ( n80 ) & ( n906 )  ;
assign n1993 =  ( n80 ) & ( n908 )  ;
assign n1994 =  ( n80 ) & ( n910 )  ;
assign n1995 =  ( n81 ) & ( n880 )  ;
assign n1996 =  ( n81 ) & ( n882 )  ;
assign n1997 =  ( n81 ) & ( n884 )  ;
assign n1998 =  ( n81 ) & ( n886 )  ;
assign n1999 =  ( n81 ) & ( n888 )  ;
assign n2000 =  ( n81 ) & ( n890 )  ;
assign n2001 =  ( n81 ) & ( n892 )  ;
assign n2002 =  ( n81 ) & ( n894 )  ;
assign n2003 =  ( n81 ) & ( n896 )  ;
assign n2004 =  ( n81 ) & ( n898 )  ;
assign n2005 =  ( n81 ) & ( n900 )  ;
assign n2006 =  ( n81 ) & ( n902 )  ;
assign n2007 =  ( n81 ) & ( n904 )  ;
assign n2008 =  ( n81 ) & ( n906 )  ;
assign n2009 =  ( n81 ) & ( n908 )  ;
assign n2010 =  ( n81 ) & ( n910 )  ;
assign n2011 =  ( n82 ) & ( n880 )  ;
assign n2012 =  ( n82 ) & ( n882 )  ;
assign n2013 =  ( n82 ) & ( n884 )  ;
assign n2014 =  ( n82 ) & ( n886 )  ;
assign n2015 =  ( n82 ) & ( n888 )  ;
assign n2016 =  ( n82 ) & ( n890 )  ;
assign n2017 =  ( n82 ) & ( n892 )  ;
assign n2018 =  ( n82 ) & ( n894 )  ;
assign n2019 =  ( n82 ) & ( n896 )  ;
assign n2020 =  ( n82 ) & ( n898 )  ;
assign n2021 =  ( n82 ) & ( n900 )  ;
assign n2022 =  ( n82 ) & ( n902 )  ;
assign n2023 =  ( n82 ) & ( n904 )  ;
assign n2024 =  ( n82 ) & ( n906 )  ;
assign n2025 =  ( n82 ) & ( n908 )  ;
assign n2026 =  ( n82 ) & ( n910 )  ;
assign n2027 =  ( n83 ) & ( n880 )  ;
assign n2028 =  ( n83 ) & ( n882 )  ;
assign n2029 =  ( n83 ) & ( n884 )  ;
assign n2030 =  ( n83 ) & ( n886 )  ;
assign n2031 =  ( n83 ) & ( n888 )  ;
assign n2032 =  ( n83 ) & ( n890 )  ;
assign n2033 =  ( n83 ) & ( n892 )  ;
assign n2034 =  ( n83 ) & ( n894 )  ;
assign n2035 =  ( n83 ) & ( n896 )  ;
assign n2036 =  ( n83 ) & ( n898 )  ;
assign n2037 =  ( n83 ) & ( n900 )  ;
assign n2038 =  ( n83 ) & ( n902 )  ;
assign n2039 =  ( n83 ) & ( n904 )  ;
assign n2040 =  ( n83 ) & ( n906 )  ;
assign n2041 =  ( n83 ) & ( n908 )  ;
assign n2042 =  ( n83 ) & ( n910 )  ;
assign n2043 =  ( n84 ) & ( n880 )  ;
assign n2044 =  ( n84 ) & ( n882 )  ;
assign n2045 =  ( n84 ) & ( n884 )  ;
assign n2046 =  ( n84 ) & ( n886 )  ;
assign n2047 =  ( n84 ) & ( n888 )  ;
assign n2048 =  ( n84 ) & ( n890 )  ;
assign n2049 =  ( n84 ) & ( n892 )  ;
assign n2050 =  ( n84 ) & ( n894 )  ;
assign n2051 =  ( n84 ) & ( n896 )  ;
assign n2052 =  ( n84 ) & ( n898 )  ;
assign n2053 =  ( n84 ) & ( n900 )  ;
assign n2054 =  ( n84 ) & ( n902 )  ;
assign n2055 =  ( n84 ) & ( n904 )  ;
assign n2056 =  ( n84 ) & ( n906 )  ;
assign n2057 =  ( n84 ) & ( n908 )  ;
assign n2058 =  ( n84 ) & ( n910 )  ;
assign n2059 =  ( n85 ) & ( n880 )  ;
assign n2060 =  ( n85 ) & ( n882 )  ;
assign n2061 =  ( n85 ) & ( n884 )  ;
assign n2062 =  ( n85 ) & ( n886 )  ;
assign n2063 =  ( n85 ) & ( n888 )  ;
assign n2064 =  ( n85 ) & ( n890 )  ;
assign n2065 =  ( n85 ) & ( n892 )  ;
assign n2066 =  ( n85 ) & ( n894 )  ;
assign n2067 =  ( n85 ) & ( n896 )  ;
assign n2068 =  ( n85 ) & ( n898 )  ;
assign n2069 =  ( n85 ) & ( n900 )  ;
assign n2070 =  ( n85 ) & ( n902 )  ;
assign n2071 =  ( n85 ) & ( n904 )  ;
assign n2072 =  ( n85 ) & ( n906 )  ;
assign n2073 =  ( n85 ) & ( n908 )  ;
assign n2074 =  ( n85 ) & ( n910 )  ;
assign n2075 =  ( n86 ) & ( n880 )  ;
assign n2076 =  ( n86 ) & ( n882 )  ;
assign n2077 =  ( n86 ) & ( n884 )  ;
assign n2078 =  ( n86 ) & ( n886 )  ;
assign n2079 =  ( n86 ) & ( n888 )  ;
assign n2080 =  ( n86 ) & ( n890 )  ;
assign n2081 =  ( n86 ) & ( n892 )  ;
assign n2082 =  ( n86 ) & ( n894 )  ;
assign n2083 =  ( n86 ) & ( n896 )  ;
assign n2084 =  ( n86 ) & ( n898 )  ;
assign n2085 =  ( n86 ) & ( n900 )  ;
assign n2086 =  ( n86 ) & ( n902 )  ;
assign n2087 =  ( n86 ) & ( n904 )  ;
assign n2088 =  ( n86 ) & ( n906 )  ;
assign n2089 =  ( n86 ) & ( n908 )  ;
assign n2090 =  ( n86 ) & ( n910 )  ;
assign n2091 =  ( n87 ) & ( n880 )  ;
assign n2092 =  ( n87 ) & ( n882 )  ;
assign n2093 =  ( n87 ) & ( n884 )  ;
assign n2094 =  ( n87 ) & ( n886 )  ;
assign n2095 =  ( n87 ) & ( n888 )  ;
assign n2096 =  ( n87 ) & ( n890 )  ;
assign n2097 =  ( n87 ) & ( n892 )  ;
assign n2098 =  ( n87 ) & ( n894 )  ;
assign n2099 =  ( n87 ) & ( n896 )  ;
assign n2100 =  ( n87 ) & ( n898 )  ;
assign n2101 =  ( n87 ) & ( n900 )  ;
assign n2102 =  ( n87 ) & ( n902 )  ;
assign n2103 =  ( n87 ) & ( n904 )  ;
assign n2104 =  ( n87 ) & ( n906 )  ;
assign n2105 =  ( n87 ) & ( n908 )  ;
assign n2106 =  ( n87 ) & ( n910 )  ;
assign n2107 =  ( n88 ) & ( n880 )  ;
assign n2108 =  ( n88 ) & ( n882 )  ;
assign n2109 =  ( n88 ) & ( n884 )  ;
assign n2110 =  ( n88 ) & ( n886 )  ;
assign n2111 =  ( n88 ) & ( n888 )  ;
assign n2112 =  ( n88 ) & ( n890 )  ;
assign n2113 =  ( n88 ) & ( n892 )  ;
assign n2114 =  ( n88 ) & ( n894 )  ;
assign n2115 =  ( n88 ) & ( n896 )  ;
assign n2116 =  ( n88 ) & ( n898 )  ;
assign n2117 =  ( n88 ) & ( n900 )  ;
assign n2118 =  ( n88 ) & ( n902 )  ;
assign n2119 =  ( n88 ) & ( n904 )  ;
assign n2120 =  ( n88 ) & ( n906 )  ;
assign n2121 =  ( n88 ) & ( n908 )  ;
assign n2122 =  ( n88 ) & ( n910 )  ;
assign n2123 =  ( n89 ) & ( n880 )  ;
assign n2124 =  ( n89 ) & ( n882 )  ;
assign n2125 =  ( n89 ) & ( n884 )  ;
assign n2126 =  ( n89 ) & ( n886 )  ;
assign n2127 =  ( n89 ) & ( n888 )  ;
assign n2128 =  ( n89 ) & ( n890 )  ;
assign n2129 =  ( n89 ) & ( n892 )  ;
assign n2130 =  ( n89 ) & ( n894 )  ;
assign n2131 =  ( n89 ) & ( n896 )  ;
assign n2132 =  ( n89 ) & ( n898 )  ;
assign n2133 =  ( n89 ) & ( n900 )  ;
assign n2134 =  ( n89 ) & ( n902 )  ;
assign n2135 =  ( n89 ) & ( n904 )  ;
assign n2136 =  ( n89 ) & ( n906 )  ;
assign n2137 =  ( n89 ) & ( n908 )  ;
assign n2138 =  ( n89 ) & ( n910 )  ;
assign n2139 =  ( n90 ) & ( n880 )  ;
assign n2140 =  ( n90 ) & ( n882 )  ;
assign n2141 =  ( n90 ) & ( n884 )  ;
assign n2142 =  ( n90 ) & ( n886 )  ;
assign n2143 =  ( n90 ) & ( n888 )  ;
assign n2144 =  ( n90 ) & ( n890 )  ;
assign n2145 =  ( n90 ) & ( n892 )  ;
assign n2146 =  ( n90 ) & ( n894 )  ;
assign n2147 =  ( n90 ) & ( n896 )  ;
assign n2148 =  ( n90 ) & ( n898 )  ;
assign n2149 =  ( n90 ) & ( n900 )  ;
assign n2150 =  ( n90 ) & ( n902 )  ;
assign n2151 =  ( n90 ) & ( n904 )  ;
assign n2152 =  ( n90 ) & ( n906 )  ;
assign n2153 =  ( n90 ) & ( n908 )  ;
assign n2154 =  ( n90 ) & ( n910 )  ;
assign n2155 =  ( n91 ) & ( n880 )  ;
assign n2156 =  ( n91 ) & ( n882 )  ;
assign n2157 =  ( n91 ) & ( n884 )  ;
assign n2158 =  ( n91 ) & ( n886 )  ;
assign n2159 =  ( n91 ) & ( n888 )  ;
assign n2160 =  ( n91 ) & ( n890 )  ;
assign n2161 =  ( n91 ) & ( n892 )  ;
assign n2162 =  ( n91 ) & ( n894 )  ;
assign n2163 =  ( n91 ) & ( n896 )  ;
assign n2164 =  ( n91 ) & ( n898 )  ;
assign n2165 =  ( n91 ) & ( n900 )  ;
assign n2166 =  ( n91 ) & ( n902 )  ;
assign n2167 =  ( n91 ) & ( n904 )  ;
assign n2168 =  ( n91 ) & ( n906 )  ;
assign n2169 =  ( n91 ) & ( n908 )  ;
assign n2170 =  ( n91 ) & ( n910 )  ;
assign n2171 =  ( n92 ) & ( n880 )  ;
assign n2172 =  ( n92 ) & ( n882 )  ;
assign n2173 =  ( n92 ) & ( n884 )  ;
assign n2174 =  ( n92 ) & ( n886 )  ;
assign n2175 =  ( n92 ) & ( n888 )  ;
assign n2176 =  ( n92 ) & ( n890 )  ;
assign n2177 =  ( n92 ) & ( n892 )  ;
assign n2178 =  ( n92 ) & ( n894 )  ;
assign n2179 =  ( n92 ) & ( n896 )  ;
assign n2180 =  ( n92 ) & ( n898 )  ;
assign n2181 =  ( n92 ) & ( n900 )  ;
assign n2182 =  ( n92 ) & ( n902 )  ;
assign n2183 =  ( n92 ) & ( n904 )  ;
assign n2184 =  ( n92 ) & ( n906 )  ;
assign n2185 =  ( n92 ) & ( n908 )  ;
assign n2186 =  ( n92 ) & ( n910 )  ;
assign n2187 =  ( n93 ) & ( n880 )  ;
assign n2188 =  ( n93 ) & ( n882 )  ;
assign n2189 =  ( n93 ) & ( n884 )  ;
assign n2190 =  ( n93 ) & ( n886 )  ;
assign n2191 =  ( n93 ) & ( n888 )  ;
assign n2192 =  ( n93 ) & ( n890 )  ;
assign n2193 =  ( n93 ) & ( n892 )  ;
assign n2194 =  ( n93 ) & ( n894 )  ;
assign n2195 =  ( n93 ) & ( n896 )  ;
assign n2196 =  ( n93 ) & ( n898 )  ;
assign n2197 =  ( n93 ) & ( n900 )  ;
assign n2198 =  ( n93 ) & ( n902 )  ;
assign n2199 =  ( n93 ) & ( n904 )  ;
assign n2200 =  ( n93 ) & ( n906 )  ;
assign n2201 =  ( n93 ) & ( n908 )  ;
assign n2202 =  ( n93 ) & ( n910 )  ;
assign n2203 =  ( n94 ) & ( n880 )  ;
assign n2204 =  ( n94 ) & ( n882 )  ;
assign n2205 =  ( n94 ) & ( n884 )  ;
assign n2206 =  ( n94 ) & ( n886 )  ;
assign n2207 =  ( n94 ) & ( n888 )  ;
assign n2208 =  ( n94 ) & ( n890 )  ;
assign n2209 =  ( n94 ) & ( n892 )  ;
assign n2210 =  ( n94 ) & ( n894 )  ;
assign n2211 =  ( n94 ) & ( n896 )  ;
assign n2212 =  ( n94 ) & ( n898 )  ;
assign n2213 =  ( n94 ) & ( n900 )  ;
assign n2214 =  ( n94 ) & ( n902 )  ;
assign n2215 =  ( n94 ) & ( n904 )  ;
assign n2216 =  ( n94 ) & ( n906 )  ;
assign n2217 =  ( n94 ) & ( n908 )  ;
assign n2218 =  ( n94 ) & ( n910 )  ;
assign n2219 =  ( n95 ) & ( n880 )  ;
assign n2220 =  ( n95 ) & ( n882 )  ;
assign n2221 =  ( n95 ) & ( n884 )  ;
assign n2222 =  ( n95 ) & ( n886 )  ;
assign n2223 =  ( n95 ) & ( n888 )  ;
assign n2224 =  ( n95 ) & ( n890 )  ;
assign n2225 =  ( n95 ) & ( n892 )  ;
assign n2226 =  ( n95 ) & ( n894 )  ;
assign n2227 =  ( n95 ) & ( n896 )  ;
assign n2228 =  ( n95 ) & ( n898 )  ;
assign n2229 =  ( n95 ) & ( n900 )  ;
assign n2230 =  ( n95 ) & ( n902 )  ;
assign n2231 =  ( n95 ) & ( n904 )  ;
assign n2232 =  ( n95 ) & ( n906 )  ;
assign n2233 =  ( n95 ) & ( n908 )  ;
assign n2234 =  ( n95 ) & ( n910 )  ;
assign n2235 =  ( n96 ) & ( n880 )  ;
assign n2236 =  ( n96 ) & ( n882 )  ;
assign n2237 =  ( n96 ) & ( n884 )  ;
assign n2238 =  ( n96 ) & ( n886 )  ;
assign n2239 =  ( n96 ) & ( n888 )  ;
assign n2240 =  ( n96 ) & ( n890 )  ;
assign n2241 =  ( n96 ) & ( n892 )  ;
assign n2242 =  ( n96 ) & ( n894 )  ;
assign n2243 =  ( n96 ) & ( n896 )  ;
assign n2244 =  ( n96 ) & ( n898 )  ;
assign n2245 =  ( n96 ) & ( n900 )  ;
assign n2246 =  ( n96 ) & ( n902 )  ;
assign n2247 =  ( n96 ) & ( n904 )  ;
assign n2248 =  ( n96 ) & ( n906 )  ;
assign n2249 =  ( n96 ) & ( n908 )  ;
assign n2250 =  ( n96 ) & ( n910 )  ;
assign n2251 =  ( n97 ) & ( n880 )  ;
assign n2252 =  ( n97 ) & ( n882 )  ;
assign n2253 =  ( n97 ) & ( n884 )  ;
assign n2254 =  ( n97 ) & ( n886 )  ;
assign n2255 =  ( n97 ) & ( n888 )  ;
assign n2256 =  ( n97 ) & ( n890 )  ;
assign n2257 =  ( n97 ) & ( n892 )  ;
assign n2258 =  ( n97 ) & ( n894 )  ;
assign n2259 =  ( n97 ) & ( n896 )  ;
assign n2260 =  ( n97 ) & ( n898 )  ;
assign n2261 =  ( n97 ) & ( n900 )  ;
assign n2262 =  ( n97 ) & ( n902 )  ;
assign n2263 =  ( n97 ) & ( n904 )  ;
assign n2264 =  ( n97 ) & ( n906 )  ;
assign n2265 =  ( n97 ) & ( n908 )  ;
assign n2266 =  ( n97 ) & ( n910 )  ;
assign n2267 =  ( n98 ) & ( n880 )  ;
assign n2268 =  ( n98 ) & ( n882 )  ;
assign n2269 =  ( n98 ) & ( n884 )  ;
assign n2270 =  ( n98 ) & ( n886 )  ;
assign n2271 =  ( n98 ) & ( n888 )  ;
assign n2272 =  ( n98 ) & ( n890 )  ;
assign n2273 =  ( n98 ) & ( n892 )  ;
assign n2274 =  ( n98 ) & ( n894 )  ;
assign n2275 =  ( n98 ) & ( n896 )  ;
assign n2276 =  ( n98 ) & ( n898 )  ;
assign n2277 =  ( n98 ) & ( n900 )  ;
assign n2278 =  ( n98 ) & ( n902 )  ;
assign n2279 =  ( n98 ) & ( n904 )  ;
assign n2280 =  ( n98 ) & ( n906 )  ;
assign n2281 =  ( n98 ) & ( n908 )  ;
assign n2282 =  ( n98 ) & ( n910 )  ;
assign n2283 =  ( n99 ) & ( n880 )  ;
assign n2284 =  ( n99 ) & ( n882 )  ;
assign n2285 =  ( n99 ) & ( n884 )  ;
assign n2286 =  ( n99 ) & ( n886 )  ;
assign n2287 =  ( n99 ) & ( n888 )  ;
assign n2288 =  ( n99 ) & ( n890 )  ;
assign n2289 =  ( n99 ) & ( n892 )  ;
assign n2290 =  ( n99 ) & ( n894 )  ;
assign n2291 =  ( n99 ) & ( n896 )  ;
assign n2292 =  ( n99 ) & ( n898 )  ;
assign n2293 =  ( n99 ) & ( n900 )  ;
assign n2294 =  ( n99 ) & ( n902 )  ;
assign n2295 =  ( n99 ) & ( n904 )  ;
assign n2296 =  ( n99 ) & ( n906 )  ;
assign n2297 =  ( n99 ) & ( n908 )  ;
assign n2298 =  ( n99 ) & ( n910 )  ;
assign n2299 =  ( n100 ) & ( n880 )  ;
assign n2300 =  ( n100 ) & ( n882 )  ;
assign n2301 =  ( n100 ) & ( n884 )  ;
assign n2302 =  ( n100 ) & ( n886 )  ;
assign n2303 =  ( n100 ) & ( n888 )  ;
assign n2304 =  ( n100 ) & ( n890 )  ;
assign n2305 =  ( n100 ) & ( n892 )  ;
assign n2306 =  ( n100 ) & ( n894 )  ;
assign n2307 =  ( n100 ) & ( n896 )  ;
assign n2308 =  ( n100 ) & ( n898 )  ;
assign n2309 =  ( n100 ) & ( n900 )  ;
assign n2310 =  ( n100 ) & ( n902 )  ;
assign n2311 =  ( n100 ) & ( n904 )  ;
assign n2312 =  ( n100 ) & ( n906 )  ;
assign n2313 =  ( n100 ) & ( n908 )  ;
assign n2314 =  ( n100 ) & ( n910 )  ;
assign n2315 =  ( n101 ) & ( n880 )  ;
assign n2316 =  ( n101 ) & ( n882 )  ;
assign n2317 =  ( n101 ) & ( n884 )  ;
assign n2318 =  ( n101 ) & ( n886 )  ;
assign n2319 =  ( n101 ) & ( n888 )  ;
assign n2320 =  ( n101 ) & ( n890 )  ;
assign n2321 =  ( n101 ) & ( n892 )  ;
assign n2322 =  ( n101 ) & ( n894 )  ;
assign n2323 =  ( n101 ) & ( n896 )  ;
assign n2324 =  ( n101 ) & ( n898 )  ;
assign n2325 =  ( n101 ) & ( n900 )  ;
assign n2326 =  ( n101 ) & ( n902 )  ;
assign n2327 =  ( n101 ) & ( n904 )  ;
assign n2328 =  ( n101 ) & ( n906 )  ;
assign n2329 =  ( n101 ) & ( n908 )  ;
assign n2330 =  ( n101 ) & ( n910 )  ;
assign n2331 =  ( n102 ) & ( n880 )  ;
assign n2332 =  ( n102 ) & ( n882 )  ;
assign n2333 =  ( n102 ) & ( n884 )  ;
assign n2334 =  ( n102 ) & ( n886 )  ;
assign n2335 =  ( n102 ) & ( n888 )  ;
assign n2336 =  ( n102 ) & ( n890 )  ;
assign n2337 =  ( n102 ) & ( n892 )  ;
assign n2338 =  ( n102 ) & ( n894 )  ;
assign n2339 =  ( n102 ) & ( n896 )  ;
assign n2340 =  ( n102 ) & ( n898 )  ;
assign n2341 =  ( n102 ) & ( n900 )  ;
assign n2342 =  ( n102 ) & ( n902 )  ;
assign n2343 =  ( n102 ) & ( n904 )  ;
assign n2344 =  ( n102 ) & ( n906 )  ;
assign n2345 =  ( n102 ) & ( n908 )  ;
assign n2346 =  ( n102 ) & ( n910 )  ;
assign n2347 =  ( n103 ) & ( n880 )  ;
assign n2348 =  ( n103 ) & ( n882 )  ;
assign n2349 =  ( n103 ) & ( n884 )  ;
assign n2350 =  ( n103 ) & ( n886 )  ;
assign n2351 =  ( n103 ) & ( n888 )  ;
assign n2352 =  ( n103 ) & ( n890 )  ;
assign n2353 =  ( n103 ) & ( n892 )  ;
assign n2354 =  ( n103 ) & ( n894 )  ;
assign n2355 =  ( n103 ) & ( n896 )  ;
assign n2356 =  ( n103 ) & ( n898 )  ;
assign n2357 =  ( n103 ) & ( n900 )  ;
assign n2358 =  ( n103 ) & ( n902 )  ;
assign n2359 =  ( n103 ) & ( n904 )  ;
assign n2360 =  ( n103 ) & ( n906 )  ;
assign n2361 =  ( n103 ) & ( n908 )  ;
assign n2362 =  ( n103 ) & ( n910 )  ;
assign n2363 =  ( n104 ) & ( n880 )  ;
assign n2364 =  ( n104 ) & ( n882 )  ;
assign n2365 =  ( n104 ) & ( n884 )  ;
assign n2366 =  ( n104 ) & ( n886 )  ;
assign n2367 =  ( n104 ) & ( n888 )  ;
assign n2368 =  ( n104 ) & ( n890 )  ;
assign n2369 =  ( n104 ) & ( n892 )  ;
assign n2370 =  ( n104 ) & ( n894 )  ;
assign n2371 =  ( n104 ) & ( n896 )  ;
assign n2372 =  ( n104 ) & ( n898 )  ;
assign n2373 =  ( n104 ) & ( n900 )  ;
assign n2374 =  ( n104 ) & ( n902 )  ;
assign n2375 =  ( n104 ) & ( n904 )  ;
assign n2376 =  ( n104 ) & ( n906 )  ;
assign n2377 =  ( n104 ) & ( n908 )  ;
assign n2378 =  ( n104 ) & ( n910 )  ;
assign n2379 =  ( n105 ) & ( n880 )  ;
assign n2380 =  ( n105 ) & ( n882 )  ;
assign n2381 =  ( n105 ) & ( n884 )  ;
assign n2382 =  ( n105 ) & ( n886 )  ;
assign n2383 =  ( n105 ) & ( n888 )  ;
assign n2384 =  ( n105 ) & ( n890 )  ;
assign n2385 =  ( n105 ) & ( n892 )  ;
assign n2386 =  ( n105 ) & ( n894 )  ;
assign n2387 =  ( n105 ) & ( n896 )  ;
assign n2388 =  ( n105 ) & ( n898 )  ;
assign n2389 =  ( n105 ) & ( n900 )  ;
assign n2390 =  ( n105 ) & ( n902 )  ;
assign n2391 =  ( n105 ) & ( n904 )  ;
assign n2392 =  ( n105 ) & ( n906 )  ;
assign n2393 =  ( n105 ) & ( n908 )  ;
assign n2394 =  ( n105 ) & ( n910 )  ;
assign n2395 =  ( n106 ) & ( n880 )  ;
assign n2396 =  ( n106 ) & ( n882 )  ;
assign n2397 =  ( n106 ) & ( n884 )  ;
assign n2398 =  ( n106 ) & ( n886 )  ;
assign n2399 =  ( n106 ) & ( n888 )  ;
assign n2400 =  ( n106 ) & ( n890 )  ;
assign n2401 =  ( n106 ) & ( n892 )  ;
assign n2402 =  ( n106 ) & ( n894 )  ;
assign n2403 =  ( n106 ) & ( n896 )  ;
assign n2404 =  ( n106 ) & ( n898 )  ;
assign n2405 =  ( n106 ) & ( n900 )  ;
assign n2406 =  ( n106 ) & ( n902 )  ;
assign n2407 =  ( n106 ) & ( n904 )  ;
assign n2408 =  ( n106 ) & ( n906 )  ;
assign n2409 =  ( n106 ) & ( n908 )  ;
assign n2410 =  ( n106 ) & ( n910 )  ;
assign n2411 =  ( n107 ) & ( n880 )  ;
assign n2412 =  ( n107 ) & ( n882 )  ;
assign n2413 =  ( n107 ) & ( n884 )  ;
assign n2414 =  ( n107 ) & ( n886 )  ;
assign n2415 =  ( n107 ) & ( n888 )  ;
assign n2416 =  ( n107 ) & ( n890 )  ;
assign n2417 =  ( n107 ) & ( n892 )  ;
assign n2418 =  ( n107 ) & ( n894 )  ;
assign n2419 =  ( n107 ) & ( n896 )  ;
assign n2420 =  ( n107 ) & ( n898 )  ;
assign n2421 =  ( n107 ) & ( n900 )  ;
assign n2422 =  ( n107 ) & ( n902 )  ;
assign n2423 =  ( n107 ) & ( n904 )  ;
assign n2424 =  ( n107 ) & ( n906 )  ;
assign n2425 =  ( n107 ) & ( n908 )  ;
assign n2426 =  ( n107 ) & ( n910 )  ;
assign n2427 =  ( n108 ) & ( n880 )  ;
assign n2428 =  ( n108 ) & ( n882 )  ;
assign n2429 =  ( n108 ) & ( n884 )  ;
assign n2430 =  ( n108 ) & ( n886 )  ;
assign n2431 =  ( n108 ) & ( n888 )  ;
assign n2432 =  ( n108 ) & ( n890 )  ;
assign n2433 =  ( n108 ) & ( n892 )  ;
assign n2434 =  ( n108 ) & ( n894 )  ;
assign n2435 =  ( n108 ) & ( n896 )  ;
assign n2436 =  ( n108 ) & ( n898 )  ;
assign n2437 =  ( n108 ) & ( n900 )  ;
assign n2438 =  ( n108 ) & ( n902 )  ;
assign n2439 =  ( n108 ) & ( n904 )  ;
assign n2440 =  ( n108 ) & ( n906 )  ;
assign n2441 =  ( n108 ) & ( n908 )  ;
assign n2442 =  ( n108 ) & ( n910 )  ;
assign n2443 =  ( n2442 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n2444 =  ( n2441 ) ? ( VREG_0_1 ) : ( n2443 ) ;
assign n2445 =  ( n2440 ) ? ( VREG_0_2 ) : ( n2444 ) ;
assign n2446 =  ( n2439 ) ? ( VREG_0_3 ) : ( n2445 ) ;
assign n2447 =  ( n2438 ) ? ( VREG_0_4 ) : ( n2446 ) ;
assign n2448 =  ( n2437 ) ? ( VREG_0_5 ) : ( n2447 ) ;
assign n2449 =  ( n2436 ) ? ( VREG_0_6 ) : ( n2448 ) ;
assign n2450 =  ( n2435 ) ? ( VREG_0_7 ) : ( n2449 ) ;
assign n2451 =  ( n2434 ) ? ( VREG_0_8 ) : ( n2450 ) ;
assign n2452 =  ( n2433 ) ? ( VREG_0_9 ) : ( n2451 ) ;
assign n2453 =  ( n2432 ) ? ( VREG_0_10 ) : ( n2452 ) ;
assign n2454 =  ( n2431 ) ? ( VREG_0_11 ) : ( n2453 ) ;
assign n2455 =  ( n2430 ) ? ( VREG_0_12 ) : ( n2454 ) ;
assign n2456 =  ( n2429 ) ? ( VREG_0_13 ) : ( n2455 ) ;
assign n2457 =  ( n2428 ) ? ( VREG_0_14 ) : ( n2456 ) ;
assign n2458 =  ( n2427 ) ? ( VREG_0_15 ) : ( n2457 ) ;
assign n2459 =  ( n2426 ) ? ( VREG_1_0 ) : ( n2458 ) ;
assign n2460 =  ( n2425 ) ? ( VREG_1_1 ) : ( n2459 ) ;
assign n2461 =  ( n2424 ) ? ( VREG_1_2 ) : ( n2460 ) ;
assign n2462 =  ( n2423 ) ? ( VREG_1_3 ) : ( n2461 ) ;
assign n2463 =  ( n2422 ) ? ( VREG_1_4 ) : ( n2462 ) ;
assign n2464 =  ( n2421 ) ? ( VREG_1_5 ) : ( n2463 ) ;
assign n2465 =  ( n2420 ) ? ( VREG_1_6 ) : ( n2464 ) ;
assign n2466 =  ( n2419 ) ? ( VREG_1_7 ) : ( n2465 ) ;
assign n2467 =  ( n2418 ) ? ( VREG_1_8 ) : ( n2466 ) ;
assign n2468 =  ( n2417 ) ? ( VREG_1_9 ) : ( n2467 ) ;
assign n2469 =  ( n2416 ) ? ( VREG_1_10 ) : ( n2468 ) ;
assign n2470 =  ( n2415 ) ? ( VREG_1_11 ) : ( n2469 ) ;
assign n2471 =  ( n2414 ) ? ( VREG_1_12 ) : ( n2470 ) ;
assign n2472 =  ( n2413 ) ? ( VREG_1_13 ) : ( n2471 ) ;
assign n2473 =  ( n2412 ) ? ( VREG_1_14 ) : ( n2472 ) ;
assign n2474 =  ( n2411 ) ? ( VREG_1_15 ) : ( n2473 ) ;
assign n2475 =  ( n2410 ) ? ( VREG_2_0 ) : ( n2474 ) ;
assign n2476 =  ( n2409 ) ? ( VREG_2_1 ) : ( n2475 ) ;
assign n2477 =  ( n2408 ) ? ( VREG_2_2 ) : ( n2476 ) ;
assign n2478 =  ( n2407 ) ? ( VREG_2_3 ) : ( n2477 ) ;
assign n2479 =  ( n2406 ) ? ( VREG_2_4 ) : ( n2478 ) ;
assign n2480 =  ( n2405 ) ? ( VREG_2_5 ) : ( n2479 ) ;
assign n2481 =  ( n2404 ) ? ( VREG_2_6 ) : ( n2480 ) ;
assign n2482 =  ( n2403 ) ? ( VREG_2_7 ) : ( n2481 ) ;
assign n2483 =  ( n2402 ) ? ( VREG_2_8 ) : ( n2482 ) ;
assign n2484 =  ( n2401 ) ? ( VREG_2_9 ) : ( n2483 ) ;
assign n2485 =  ( n2400 ) ? ( VREG_2_10 ) : ( n2484 ) ;
assign n2486 =  ( n2399 ) ? ( VREG_2_11 ) : ( n2485 ) ;
assign n2487 =  ( n2398 ) ? ( VREG_2_12 ) : ( n2486 ) ;
assign n2488 =  ( n2397 ) ? ( VREG_2_13 ) : ( n2487 ) ;
assign n2489 =  ( n2396 ) ? ( VREG_2_14 ) : ( n2488 ) ;
assign n2490 =  ( n2395 ) ? ( VREG_2_15 ) : ( n2489 ) ;
assign n2491 =  ( n2394 ) ? ( VREG_3_0 ) : ( n2490 ) ;
assign n2492 =  ( n2393 ) ? ( VREG_3_1 ) : ( n2491 ) ;
assign n2493 =  ( n2392 ) ? ( VREG_3_2 ) : ( n2492 ) ;
assign n2494 =  ( n2391 ) ? ( VREG_3_3 ) : ( n2493 ) ;
assign n2495 =  ( n2390 ) ? ( VREG_3_4 ) : ( n2494 ) ;
assign n2496 =  ( n2389 ) ? ( VREG_3_5 ) : ( n2495 ) ;
assign n2497 =  ( n2388 ) ? ( VREG_3_6 ) : ( n2496 ) ;
assign n2498 =  ( n2387 ) ? ( VREG_3_7 ) : ( n2497 ) ;
assign n2499 =  ( n2386 ) ? ( VREG_3_8 ) : ( n2498 ) ;
assign n2500 =  ( n2385 ) ? ( VREG_3_9 ) : ( n2499 ) ;
assign n2501 =  ( n2384 ) ? ( VREG_3_10 ) : ( n2500 ) ;
assign n2502 =  ( n2383 ) ? ( VREG_3_11 ) : ( n2501 ) ;
assign n2503 =  ( n2382 ) ? ( VREG_3_12 ) : ( n2502 ) ;
assign n2504 =  ( n2381 ) ? ( VREG_3_13 ) : ( n2503 ) ;
assign n2505 =  ( n2380 ) ? ( VREG_3_14 ) : ( n2504 ) ;
assign n2506 =  ( n2379 ) ? ( VREG_3_15 ) : ( n2505 ) ;
assign n2507 =  ( n2378 ) ? ( VREG_4_0 ) : ( n2506 ) ;
assign n2508 =  ( n2377 ) ? ( VREG_4_1 ) : ( n2507 ) ;
assign n2509 =  ( n2376 ) ? ( VREG_4_2 ) : ( n2508 ) ;
assign n2510 =  ( n2375 ) ? ( VREG_4_3 ) : ( n2509 ) ;
assign n2511 =  ( n2374 ) ? ( VREG_4_4 ) : ( n2510 ) ;
assign n2512 =  ( n2373 ) ? ( VREG_4_5 ) : ( n2511 ) ;
assign n2513 =  ( n2372 ) ? ( VREG_4_6 ) : ( n2512 ) ;
assign n2514 =  ( n2371 ) ? ( VREG_4_7 ) : ( n2513 ) ;
assign n2515 =  ( n2370 ) ? ( VREG_4_8 ) : ( n2514 ) ;
assign n2516 =  ( n2369 ) ? ( VREG_4_9 ) : ( n2515 ) ;
assign n2517 =  ( n2368 ) ? ( VREG_4_10 ) : ( n2516 ) ;
assign n2518 =  ( n2367 ) ? ( VREG_4_11 ) : ( n2517 ) ;
assign n2519 =  ( n2366 ) ? ( VREG_4_12 ) : ( n2518 ) ;
assign n2520 =  ( n2365 ) ? ( VREG_4_13 ) : ( n2519 ) ;
assign n2521 =  ( n2364 ) ? ( VREG_4_14 ) : ( n2520 ) ;
assign n2522 =  ( n2363 ) ? ( VREG_4_15 ) : ( n2521 ) ;
assign n2523 =  ( n2362 ) ? ( VREG_5_0 ) : ( n2522 ) ;
assign n2524 =  ( n2361 ) ? ( VREG_5_1 ) : ( n2523 ) ;
assign n2525 =  ( n2360 ) ? ( VREG_5_2 ) : ( n2524 ) ;
assign n2526 =  ( n2359 ) ? ( VREG_5_3 ) : ( n2525 ) ;
assign n2527 =  ( n2358 ) ? ( VREG_5_4 ) : ( n2526 ) ;
assign n2528 =  ( n2357 ) ? ( VREG_5_5 ) : ( n2527 ) ;
assign n2529 =  ( n2356 ) ? ( VREG_5_6 ) : ( n2528 ) ;
assign n2530 =  ( n2355 ) ? ( VREG_5_7 ) : ( n2529 ) ;
assign n2531 =  ( n2354 ) ? ( VREG_5_8 ) : ( n2530 ) ;
assign n2532 =  ( n2353 ) ? ( VREG_5_9 ) : ( n2531 ) ;
assign n2533 =  ( n2352 ) ? ( VREG_5_10 ) : ( n2532 ) ;
assign n2534 =  ( n2351 ) ? ( VREG_5_11 ) : ( n2533 ) ;
assign n2535 =  ( n2350 ) ? ( VREG_5_12 ) : ( n2534 ) ;
assign n2536 =  ( n2349 ) ? ( VREG_5_13 ) : ( n2535 ) ;
assign n2537 =  ( n2348 ) ? ( VREG_5_14 ) : ( n2536 ) ;
assign n2538 =  ( n2347 ) ? ( VREG_5_15 ) : ( n2537 ) ;
assign n2539 =  ( n2346 ) ? ( VREG_6_0 ) : ( n2538 ) ;
assign n2540 =  ( n2345 ) ? ( VREG_6_1 ) : ( n2539 ) ;
assign n2541 =  ( n2344 ) ? ( VREG_6_2 ) : ( n2540 ) ;
assign n2542 =  ( n2343 ) ? ( VREG_6_3 ) : ( n2541 ) ;
assign n2543 =  ( n2342 ) ? ( VREG_6_4 ) : ( n2542 ) ;
assign n2544 =  ( n2341 ) ? ( VREG_6_5 ) : ( n2543 ) ;
assign n2545 =  ( n2340 ) ? ( VREG_6_6 ) : ( n2544 ) ;
assign n2546 =  ( n2339 ) ? ( VREG_6_7 ) : ( n2545 ) ;
assign n2547 =  ( n2338 ) ? ( VREG_6_8 ) : ( n2546 ) ;
assign n2548 =  ( n2337 ) ? ( VREG_6_9 ) : ( n2547 ) ;
assign n2549 =  ( n2336 ) ? ( VREG_6_10 ) : ( n2548 ) ;
assign n2550 =  ( n2335 ) ? ( VREG_6_11 ) : ( n2549 ) ;
assign n2551 =  ( n2334 ) ? ( VREG_6_12 ) : ( n2550 ) ;
assign n2552 =  ( n2333 ) ? ( VREG_6_13 ) : ( n2551 ) ;
assign n2553 =  ( n2332 ) ? ( VREG_6_14 ) : ( n2552 ) ;
assign n2554 =  ( n2331 ) ? ( VREG_6_15 ) : ( n2553 ) ;
assign n2555 =  ( n2330 ) ? ( VREG_7_0 ) : ( n2554 ) ;
assign n2556 =  ( n2329 ) ? ( VREG_7_1 ) : ( n2555 ) ;
assign n2557 =  ( n2328 ) ? ( VREG_7_2 ) : ( n2556 ) ;
assign n2558 =  ( n2327 ) ? ( VREG_7_3 ) : ( n2557 ) ;
assign n2559 =  ( n2326 ) ? ( VREG_7_4 ) : ( n2558 ) ;
assign n2560 =  ( n2325 ) ? ( VREG_7_5 ) : ( n2559 ) ;
assign n2561 =  ( n2324 ) ? ( VREG_7_6 ) : ( n2560 ) ;
assign n2562 =  ( n2323 ) ? ( VREG_7_7 ) : ( n2561 ) ;
assign n2563 =  ( n2322 ) ? ( VREG_7_8 ) : ( n2562 ) ;
assign n2564 =  ( n2321 ) ? ( VREG_7_9 ) : ( n2563 ) ;
assign n2565 =  ( n2320 ) ? ( VREG_7_10 ) : ( n2564 ) ;
assign n2566 =  ( n2319 ) ? ( VREG_7_11 ) : ( n2565 ) ;
assign n2567 =  ( n2318 ) ? ( VREG_7_12 ) : ( n2566 ) ;
assign n2568 =  ( n2317 ) ? ( VREG_7_13 ) : ( n2567 ) ;
assign n2569 =  ( n2316 ) ? ( VREG_7_14 ) : ( n2568 ) ;
assign n2570 =  ( n2315 ) ? ( VREG_7_15 ) : ( n2569 ) ;
assign n2571 =  ( n2314 ) ? ( VREG_8_0 ) : ( n2570 ) ;
assign n2572 =  ( n2313 ) ? ( VREG_8_1 ) : ( n2571 ) ;
assign n2573 =  ( n2312 ) ? ( VREG_8_2 ) : ( n2572 ) ;
assign n2574 =  ( n2311 ) ? ( VREG_8_3 ) : ( n2573 ) ;
assign n2575 =  ( n2310 ) ? ( VREG_8_4 ) : ( n2574 ) ;
assign n2576 =  ( n2309 ) ? ( VREG_8_5 ) : ( n2575 ) ;
assign n2577 =  ( n2308 ) ? ( VREG_8_6 ) : ( n2576 ) ;
assign n2578 =  ( n2307 ) ? ( VREG_8_7 ) : ( n2577 ) ;
assign n2579 =  ( n2306 ) ? ( VREG_8_8 ) : ( n2578 ) ;
assign n2580 =  ( n2305 ) ? ( VREG_8_9 ) : ( n2579 ) ;
assign n2581 =  ( n2304 ) ? ( VREG_8_10 ) : ( n2580 ) ;
assign n2582 =  ( n2303 ) ? ( VREG_8_11 ) : ( n2581 ) ;
assign n2583 =  ( n2302 ) ? ( VREG_8_12 ) : ( n2582 ) ;
assign n2584 =  ( n2301 ) ? ( VREG_8_13 ) : ( n2583 ) ;
assign n2585 =  ( n2300 ) ? ( VREG_8_14 ) : ( n2584 ) ;
assign n2586 =  ( n2299 ) ? ( VREG_8_15 ) : ( n2585 ) ;
assign n2587 =  ( n2298 ) ? ( VREG_9_0 ) : ( n2586 ) ;
assign n2588 =  ( n2297 ) ? ( VREG_9_1 ) : ( n2587 ) ;
assign n2589 =  ( n2296 ) ? ( VREG_9_2 ) : ( n2588 ) ;
assign n2590 =  ( n2295 ) ? ( VREG_9_3 ) : ( n2589 ) ;
assign n2591 =  ( n2294 ) ? ( VREG_9_4 ) : ( n2590 ) ;
assign n2592 =  ( n2293 ) ? ( VREG_9_5 ) : ( n2591 ) ;
assign n2593 =  ( n2292 ) ? ( VREG_9_6 ) : ( n2592 ) ;
assign n2594 =  ( n2291 ) ? ( VREG_9_7 ) : ( n2593 ) ;
assign n2595 =  ( n2290 ) ? ( VREG_9_8 ) : ( n2594 ) ;
assign n2596 =  ( n2289 ) ? ( VREG_9_9 ) : ( n2595 ) ;
assign n2597 =  ( n2288 ) ? ( VREG_9_10 ) : ( n2596 ) ;
assign n2598 =  ( n2287 ) ? ( VREG_9_11 ) : ( n2597 ) ;
assign n2599 =  ( n2286 ) ? ( VREG_9_12 ) : ( n2598 ) ;
assign n2600 =  ( n2285 ) ? ( VREG_9_13 ) : ( n2599 ) ;
assign n2601 =  ( n2284 ) ? ( VREG_9_14 ) : ( n2600 ) ;
assign n2602 =  ( n2283 ) ? ( VREG_9_15 ) : ( n2601 ) ;
assign n2603 =  ( n2282 ) ? ( VREG_10_0 ) : ( n2602 ) ;
assign n2604 =  ( n2281 ) ? ( VREG_10_1 ) : ( n2603 ) ;
assign n2605 =  ( n2280 ) ? ( VREG_10_2 ) : ( n2604 ) ;
assign n2606 =  ( n2279 ) ? ( VREG_10_3 ) : ( n2605 ) ;
assign n2607 =  ( n2278 ) ? ( VREG_10_4 ) : ( n2606 ) ;
assign n2608 =  ( n2277 ) ? ( VREG_10_5 ) : ( n2607 ) ;
assign n2609 =  ( n2276 ) ? ( VREG_10_6 ) : ( n2608 ) ;
assign n2610 =  ( n2275 ) ? ( VREG_10_7 ) : ( n2609 ) ;
assign n2611 =  ( n2274 ) ? ( VREG_10_8 ) : ( n2610 ) ;
assign n2612 =  ( n2273 ) ? ( VREG_10_9 ) : ( n2611 ) ;
assign n2613 =  ( n2272 ) ? ( VREG_10_10 ) : ( n2612 ) ;
assign n2614 =  ( n2271 ) ? ( VREG_10_11 ) : ( n2613 ) ;
assign n2615 =  ( n2270 ) ? ( VREG_10_12 ) : ( n2614 ) ;
assign n2616 =  ( n2269 ) ? ( VREG_10_13 ) : ( n2615 ) ;
assign n2617 =  ( n2268 ) ? ( VREG_10_14 ) : ( n2616 ) ;
assign n2618 =  ( n2267 ) ? ( VREG_10_15 ) : ( n2617 ) ;
assign n2619 =  ( n2266 ) ? ( VREG_11_0 ) : ( n2618 ) ;
assign n2620 =  ( n2265 ) ? ( VREG_11_1 ) : ( n2619 ) ;
assign n2621 =  ( n2264 ) ? ( VREG_11_2 ) : ( n2620 ) ;
assign n2622 =  ( n2263 ) ? ( VREG_11_3 ) : ( n2621 ) ;
assign n2623 =  ( n2262 ) ? ( VREG_11_4 ) : ( n2622 ) ;
assign n2624 =  ( n2261 ) ? ( VREG_11_5 ) : ( n2623 ) ;
assign n2625 =  ( n2260 ) ? ( VREG_11_6 ) : ( n2624 ) ;
assign n2626 =  ( n2259 ) ? ( VREG_11_7 ) : ( n2625 ) ;
assign n2627 =  ( n2258 ) ? ( VREG_11_8 ) : ( n2626 ) ;
assign n2628 =  ( n2257 ) ? ( VREG_11_9 ) : ( n2627 ) ;
assign n2629 =  ( n2256 ) ? ( VREG_11_10 ) : ( n2628 ) ;
assign n2630 =  ( n2255 ) ? ( VREG_11_11 ) : ( n2629 ) ;
assign n2631 =  ( n2254 ) ? ( VREG_11_12 ) : ( n2630 ) ;
assign n2632 =  ( n2253 ) ? ( VREG_11_13 ) : ( n2631 ) ;
assign n2633 =  ( n2252 ) ? ( VREG_11_14 ) : ( n2632 ) ;
assign n2634 =  ( n2251 ) ? ( VREG_11_15 ) : ( n2633 ) ;
assign n2635 =  ( n2250 ) ? ( VREG_12_0 ) : ( n2634 ) ;
assign n2636 =  ( n2249 ) ? ( VREG_12_1 ) : ( n2635 ) ;
assign n2637 =  ( n2248 ) ? ( VREG_12_2 ) : ( n2636 ) ;
assign n2638 =  ( n2247 ) ? ( VREG_12_3 ) : ( n2637 ) ;
assign n2639 =  ( n2246 ) ? ( VREG_12_4 ) : ( n2638 ) ;
assign n2640 =  ( n2245 ) ? ( VREG_12_5 ) : ( n2639 ) ;
assign n2641 =  ( n2244 ) ? ( VREG_12_6 ) : ( n2640 ) ;
assign n2642 =  ( n2243 ) ? ( VREG_12_7 ) : ( n2641 ) ;
assign n2643 =  ( n2242 ) ? ( VREG_12_8 ) : ( n2642 ) ;
assign n2644 =  ( n2241 ) ? ( VREG_12_9 ) : ( n2643 ) ;
assign n2645 =  ( n2240 ) ? ( VREG_12_10 ) : ( n2644 ) ;
assign n2646 =  ( n2239 ) ? ( VREG_12_11 ) : ( n2645 ) ;
assign n2647 =  ( n2238 ) ? ( VREG_12_12 ) : ( n2646 ) ;
assign n2648 =  ( n2237 ) ? ( VREG_12_13 ) : ( n2647 ) ;
assign n2649 =  ( n2236 ) ? ( VREG_12_14 ) : ( n2648 ) ;
assign n2650 =  ( n2235 ) ? ( VREG_12_15 ) : ( n2649 ) ;
assign n2651 =  ( n2234 ) ? ( VREG_13_0 ) : ( n2650 ) ;
assign n2652 =  ( n2233 ) ? ( VREG_13_1 ) : ( n2651 ) ;
assign n2653 =  ( n2232 ) ? ( VREG_13_2 ) : ( n2652 ) ;
assign n2654 =  ( n2231 ) ? ( VREG_13_3 ) : ( n2653 ) ;
assign n2655 =  ( n2230 ) ? ( VREG_13_4 ) : ( n2654 ) ;
assign n2656 =  ( n2229 ) ? ( VREG_13_5 ) : ( n2655 ) ;
assign n2657 =  ( n2228 ) ? ( VREG_13_6 ) : ( n2656 ) ;
assign n2658 =  ( n2227 ) ? ( VREG_13_7 ) : ( n2657 ) ;
assign n2659 =  ( n2226 ) ? ( VREG_13_8 ) : ( n2658 ) ;
assign n2660 =  ( n2225 ) ? ( VREG_13_9 ) : ( n2659 ) ;
assign n2661 =  ( n2224 ) ? ( VREG_13_10 ) : ( n2660 ) ;
assign n2662 =  ( n2223 ) ? ( VREG_13_11 ) : ( n2661 ) ;
assign n2663 =  ( n2222 ) ? ( VREG_13_12 ) : ( n2662 ) ;
assign n2664 =  ( n2221 ) ? ( VREG_13_13 ) : ( n2663 ) ;
assign n2665 =  ( n2220 ) ? ( VREG_13_14 ) : ( n2664 ) ;
assign n2666 =  ( n2219 ) ? ( VREG_13_15 ) : ( n2665 ) ;
assign n2667 =  ( n2218 ) ? ( VREG_14_0 ) : ( n2666 ) ;
assign n2668 =  ( n2217 ) ? ( VREG_14_1 ) : ( n2667 ) ;
assign n2669 =  ( n2216 ) ? ( VREG_14_2 ) : ( n2668 ) ;
assign n2670 =  ( n2215 ) ? ( VREG_14_3 ) : ( n2669 ) ;
assign n2671 =  ( n2214 ) ? ( VREG_14_4 ) : ( n2670 ) ;
assign n2672 =  ( n2213 ) ? ( VREG_14_5 ) : ( n2671 ) ;
assign n2673 =  ( n2212 ) ? ( VREG_14_6 ) : ( n2672 ) ;
assign n2674 =  ( n2211 ) ? ( VREG_14_7 ) : ( n2673 ) ;
assign n2675 =  ( n2210 ) ? ( VREG_14_8 ) : ( n2674 ) ;
assign n2676 =  ( n2209 ) ? ( VREG_14_9 ) : ( n2675 ) ;
assign n2677 =  ( n2208 ) ? ( VREG_14_10 ) : ( n2676 ) ;
assign n2678 =  ( n2207 ) ? ( VREG_14_11 ) : ( n2677 ) ;
assign n2679 =  ( n2206 ) ? ( VREG_14_12 ) : ( n2678 ) ;
assign n2680 =  ( n2205 ) ? ( VREG_14_13 ) : ( n2679 ) ;
assign n2681 =  ( n2204 ) ? ( VREG_14_14 ) : ( n2680 ) ;
assign n2682 =  ( n2203 ) ? ( VREG_14_15 ) : ( n2681 ) ;
assign n2683 =  ( n2202 ) ? ( VREG_15_0 ) : ( n2682 ) ;
assign n2684 =  ( n2201 ) ? ( VREG_15_1 ) : ( n2683 ) ;
assign n2685 =  ( n2200 ) ? ( VREG_15_2 ) : ( n2684 ) ;
assign n2686 =  ( n2199 ) ? ( VREG_15_3 ) : ( n2685 ) ;
assign n2687 =  ( n2198 ) ? ( VREG_15_4 ) : ( n2686 ) ;
assign n2688 =  ( n2197 ) ? ( VREG_15_5 ) : ( n2687 ) ;
assign n2689 =  ( n2196 ) ? ( VREG_15_6 ) : ( n2688 ) ;
assign n2690 =  ( n2195 ) ? ( VREG_15_7 ) : ( n2689 ) ;
assign n2691 =  ( n2194 ) ? ( VREG_15_8 ) : ( n2690 ) ;
assign n2692 =  ( n2193 ) ? ( VREG_15_9 ) : ( n2691 ) ;
assign n2693 =  ( n2192 ) ? ( VREG_15_10 ) : ( n2692 ) ;
assign n2694 =  ( n2191 ) ? ( VREG_15_11 ) : ( n2693 ) ;
assign n2695 =  ( n2190 ) ? ( VREG_15_12 ) : ( n2694 ) ;
assign n2696 =  ( n2189 ) ? ( VREG_15_13 ) : ( n2695 ) ;
assign n2697 =  ( n2188 ) ? ( VREG_15_14 ) : ( n2696 ) ;
assign n2698 =  ( n2187 ) ? ( VREG_15_15 ) : ( n2697 ) ;
assign n2699 =  ( n2186 ) ? ( VREG_16_0 ) : ( n2698 ) ;
assign n2700 =  ( n2185 ) ? ( VREG_16_1 ) : ( n2699 ) ;
assign n2701 =  ( n2184 ) ? ( VREG_16_2 ) : ( n2700 ) ;
assign n2702 =  ( n2183 ) ? ( VREG_16_3 ) : ( n2701 ) ;
assign n2703 =  ( n2182 ) ? ( VREG_16_4 ) : ( n2702 ) ;
assign n2704 =  ( n2181 ) ? ( VREG_16_5 ) : ( n2703 ) ;
assign n2705 =  ( n2180 ) ? ( VREG_16_6 ) : ( n2704 ) ;
assign n2706 =  ( n2179 ) ? ( VREG_16_7 ) : ( n2705 ) ;
assign n2707 =  ( n2178 ) ? ( VREG_16_8 ) : ( n2706 ) ;
assign n2708 =  ( n2177 ) ? ( VREG_16_9 ) : ( n2707 ) ;
assign n2709 =  ( n2176 ) ? ( VREG_16_10 ) : ( n2708 ) ;
assign n2710 =  ( n2175 ) ? ( VREG_16_11 ) : ( n2709 ) ;
assign n2711 =  ( n2174 ) ? ( VREG_16_12 ) : ( n2710 ) ;
assign n2712 =  ( n2173 ) ? ( VREG_16_13 ) : ( n2711 ) ;
assign n2713 =  ( n2172 ) ? ( VREG_16_14 ) : ( n2712 ) ;
assign n2714 =  ( n2171 ) ? ( VREG_16_15 ) : ( n2713 ) ;
assign n2715 =  ( n2170 ) ? ( VREG_17_0 ) : ( n2714 ) ;
assign n2716 =  ( n2169 ) ? ( VREG_17_1 ) : ( n2715 ) ;
assign n2717 =  ( n2168 ) ? ( VREG_17_2 ) : ( n2716 ) ;
assign n2718 =  ( n2167 ) ? ( VREG_17_3 ) : ( n2717 ) ;
assign n2719 =  ( n2166 ) ? ( VREG_17_4 ) : ( n2718 ) ;
assign n2720 =  ( n2165 ) ? ( VREG_17_5 ) : ( n2719 ) ;
assign n2721 =  ( n2164 ) ? ( VREG_17_6 ) : ( n2720 ) ;
assign n2722 =  ( n2163 ) ? ( VREG_17_7 ) : ( n2721 ) ;
assign n2723 =  ( n2162 ) ? ( VREG_17_8 ) : ( n2722 ) ;
assign n2724 =  ( n2161 ) ? ( VREG_17_9 ) : ( n2723 ) ;
assign n2725 =  ( n2160 ) ? ( VREG_17_10 ) : ( n2724 ) ;
assign n2726 =  ( n2159 ) ? ( VREG_17_11 ) : ( n2725 ) ;
assign n2727 =  ( n2158 ) ? ( VREG_17_12 ) : ( n2726 ) ;
assign n2728 =  ( n2157 ) ? ( VREG_17_13 ) : ( n2727 ) ;
assign n2729 =  ( n2156 ) ? ( VREG_17_14 ) : ( n2728 ) ;
assign n2730 =  ( n2155 ) ? ( VREG_17_15 ) : ( n2729 ) ;
assign n2731 =  ( n2154 ) ? ( VREG_18_0 ) : ( n2730 ) ;
assign n2732 =  ( n2153 ) ? ( VREG_18_1 ) : ( n2731 ) ;
assign n2733 =  ( n2152 ) ? ( VREG_18_2 ) : ( n2732 ) ;
assign n2734 =  ( n2151 ) ? ( VREG_18_3 ) : ( n2733 ) ;
assign n2735 =  ( n2150 ) ? ( VREG_18_4 ) : ( n2734 ) ;
assign n2736 =  ( n2149 ) ? ( VREG_18_5 ) : ( n2735 ) ;
assign n2737 =  ( n2148 ) ? ( VREG_18_6 ) : ( n2736 ) ;
assign n2738 =  ( n2147 ) ? ( VREG_18_7 ) : ( n2737 ) ;
assign n2739 =  ( n2146 ) ? ( VREG_18_8 ) : ( n2738 ) ;
assign n2740 =  ( n2145 ) ? ( VREG_18_9 ) : ( n2739 ) ;
assign n2741 =  ( n2144 ) ? ( VREG_18_10 ) : ( n2740 ) ;
assign n2742 =  ( n2143 ) ? ( VREG_18_11 ) : ( n2741 ) ;
assign n2743 =  ( n2142 ) ? ( VREG_18_12 ) : ( n2742 ) ;
assign n2744 =  ( n2141 ) ? ( VREG_18_13 ) : ( n2743 ) ;
assign n2745 =  ( n2140 ) ? ( VREG_18_14 ) : ( n2744 ) ;
assign n2746 =  ( n2139 ) ? ( VREG_18_15 ) : ( n2745 ) ;
assign n2747 =  ( n2138 ) ? ( VREG_19_0 ) : ( n2746 ) ;
assign n2748 =  ( n2137 ) ? ( VREG_19_1 ) : ( n2747 ) ;
assign n2749 =  ( n2136 ) ? ( VREG_19_2 ) : ( n2748 ) ;
assign n2750 =  ( n2135 ) ? ( VREG_19_3 ) : ( n2749 ) ;
assign n2751 =  ( n2134 ) ? ( VREG_19_4 ) : ( n2750 ) ;
assign n2752 =  ( n2133 ) ? ( VREG_19_5 ) : ( n2751 ) ;
assign n2753 =  ( n2132 ) ? ( VREG_19_6 ) : ( n2752 ) ;
assign n2754 =  ( n2131 ) ? ( VREG_19_7 ) : ( n2753 ) ;
assign n2755 =  ( n2130 ) ? ( VREG_19_8 ) : ( n2754 ) ;
assign n2756 =  ( n2129 ) ? ( VREG_19_9 ) : ( n2755 ) ;
assign n2757 =  ( n2128 ) ? ( VREG_19_10 ) : ( n2756 ) ;
assign n2758 =  ( n2127 ) ? ( VREG_19_11 ) : ( n2757 ) ;
assign n2759 =  ( n2126 ) ? ( VREG_19_12 ) : ( n2758 ) ;
assign n2760 =  ( n2125 ) ? ( VREG_19_13 ) : ( n2759 ) ;
assign n2761 =  ( n2124 ) ? ( VREG_19_14 ) : ( n2760 ) ;
assign n2762 =  ( n2123 ) ? ( VREG_19_15 ) : ( n2761 ) ;
assign n2763 =  ( n2122 ) ? ( VREG_20_0 ) : ( n2762 ) ;
assign n2764 =  ( n2121 ) ? ( VREG_20_1 ) : ( n2763 ) ;
assign n2765 =  ( n2120 ) ? ( VREG_20_2 ) : ( n2764 ) ;
assign n2766 =  ( n2119 ) ? ( VREG_20_3 ) : ( n2765 ) ;
assign n2767 =  ( n2118 ) ? ( VREG_20_4 ) : ( n2766 ) ;
assign n2768 =  ( n2117 ) ? ( VREG_20_5 ) : ( n2767 ) ;
assign n2769 =  ( n2116 ) ? ( VREG_20_6 ) : ( n2768 ) ;
assign n2770 =  ( n2115 ) ? ( VREG_20_7 ) : ( n2769 ) ;
assign n2771 =  ( n2114 ) ? ( VREG_20_8 ) : ( n2770 ) ;
assign n2772 =  ( n2113 ) ? ( VREG_20_9 ) : ( n2771 ) ;
assign n2773 =  ( n2112 ) ? ( VREG_20_10 ) : ( n2772 ) ;
assign n2774 =  ( n2111 ) ? ( VREG_20_11 ) : ( n2773 ) ;
assign n2775 =  ( n2110 ) ? ( VREG_20_12 ) : ( n2774 ) ;
assign n2776 =  ( n2109 ) ? ( VREG_20_13 ) : ( n2775 ) ;
assign n2777 =  ( n2108 ) ? ( VREG_20_14 ) : ( n2776 ) ;
assign n2778 =  ( n2107 ) ? ( VREG_20_15 ) : ( n2777 ) ;
assign n2779 =  ( n2106 ) ? ( VREG_21_0 ) : ( n2778 ) ;
assign n2780 =  ( n2105 ) ? ( VREG_21_1 ) : ( n2779 ) ;
assign n2781 =  ( n2104 ) ? ( VREG_21_2 ) : ( n2780 ) ;
assign n2782 =  ( n2103 ) ? ( VREG_21_3 ) : ( n2781 ) ;
assign n2783 =  ( n2102 ) ? ( VREG_21_4 ) : ( n2782 ) ;
assign n2784 =  ( n2101 ) ? ( VREG_21_5 ) : ( n2783 ) ;
assign n2785 =  ( n2100 ) ? ( VREG_21_6 ) : ( n2784 ) ;
assign n2786 =  ( n2099 ) ? ( VREG_21_7 ) : ( n2785 ) ;
assign n2787 =  ( n2098 ) ? ( VREG_21_8 ) : ( n2786 ) ;
assign n2788 =  ( n2097 ) ? ( VREG_21_9 ) : ( n2787 ) ;
assign n2789 =  ( n2096 ) ? ( VREG_21_10 ) : ( n2788 ) ;
assign n2790 =  ( n2095 ) ? ( VREG_21_11 ) : ( n2789 ) ;
assign n2791 =  ( n2094 ) ? ( VREG_21_12 ) : ( n2790 ) ;
assign n2792 =  ( n2093 ) ? ( VREG_21_13 ) : ( n2791 ) ;
assign n2793 =  ( n2092 ) ? ( VREG_21_14 ) : ( n2792 ) ;
assign n2794 =  ( n2091 ) ? ( VREG_21_15 ) : ( n2793 ) ;
assign n2795 =  ( n2090 ) ? ( VREG_22_0 ) : ( n2794 ) ;
assign n2796 =  ( n2089 ) ? ( VREG_22_1 ) : ( n2795 ) ;
assign n2797 =  ( n2088 ) ? ( VREG_22_2 ) : ( n2796 ) ;
assign n2798 =  ( n2087 ) ? ( VREG_22_3 ) : ( n2797 ) ;
assign n2799 =  ( n2086 ) ? ( VREG_22_4 ) : ( n2798 ) ;
assign n2800 =  ( n2085 ) ? ( VREG_22_5 ) : ( n2799 ) ;
assign n2801 =  ( n2084 ) ? ( VREG_22_6 ) : ( n2800 ) ;
assign n2802 =  ( n2083 ) ? ( VREG_22_7 ) : ( n2801 ) ;
assign n2803 =  ( n2082 ) ? ( VREG_22_8 ) : ( n2802 ) ;
assign n2804 =  ( n2081 ) ? ( VREG_22_9 ) : ( n2803 ) ;
assign n2805 =  ( n2080 ) ? ( VREG_22_10 ) : ( n2804 ) ;
assign n2806 =  ( n2079 ) ? ( VREG_22_11 ) : ( n2805 ) ;
assign n2807 =  ( n2078 ) ? ( VREG_22_12 ) : ( n2806 ) ;
assign n2808 =  ( n2077 ) ? ( VREG_22_13 ) : ( n2807 ) ;
assign n2809 =  ( n2076 ) ? ( VREG_22_14 ) : ( n2808 ) ;
assign n2810 =  ( n2075 ) ? ( VREG_22_15 ) : ( n2809 ) ;
assign n2811 =  ( n2074 ) ? ( VREG_23_0 ) : ( n2810 ) ;
assign n2812 =  ( n2073 ) ? ( VREG_23_1 ) : ( n2811 ) ;
assign n2813 =  ( n2072 ) ? ( VREG_23_2 ) : ( n2812 ) ;
assign n2814 =  ( n2071 ) ? ( VREG_23_3 ) : ( n2813 ) ;
assign n2815 =  ( n2070 ) ? ( VREG_23_4 ) : ( n2814 ) ;
assign n2816 =  ( n2069 ) ? ( VREG_23_5 ) : ( n2815 ) ;
assign n2817 =  ( n2068 ) ? ( VREG_23_6 ) : ( n2816 ) ;
assign n2818 =  ( n2067 ) ? ( VREG_23_7 ) : ( n2817 ) ;
assign n2819 =  ( n2066 ) ? ( VREG_23_8 ) : ( n2818 ) ;
assign n2820 =  ( n2065 ) ? ( VREG_23_9 ) : ( n2819 ) ;
assign n2821 =  ( n2064 ) ? ( VREG_23_10 ) : ( n2820 ) ;
assign n2822 =  ( n2063 ) ? ( VREG_23_11 ) : ( n2821 ) ;
assign n2823 =  ( n2062 ) ? ( VREG_23_12 ) : ( n2822 ) ;
assign n2824 =  ( n2061 ) ? ( VREG_23_13 ) : ( n2823 ) ;
assign n2825 =  ( n2060 ) ? ( VREG_23_14 ) : ( n2824 ) ;
assign n2826 =  ( n2059 ) ? ( VREG_23_15 ) : ( n2825 ) ;
assign n2827 =  ( n2058 ) ? ( VREG_24_0 ) : ( n2826 ) ;
assign n2828 =  ( n2057 ) ? ( VREG_24_1 ) : ( n2827 ) ;
assign n2829 =  ( n2056 ) ? ( VREG_24_2 ) : ( n2828 ) ;
assign n2830 =  ( n2055 ) ? ( VREG_24_3 ) : ( n2829 ) ;
assign n2831 =  ( n2054 ) ? ( VREG_24_4 ) : ( n2830 ) ;
assign n2832 =  ( n2053 ) ? ( VREG_24_5 ) : ( n2831 ) ;
assign n2833 =  ( n2052 ) ? ( VREG_24_6 ) : ( n2832 ) ;
assign n2834 =  ( n2051 ) ? ( VREG_24_7 ) : ( n2833 ) ;
assign n2835 =  ( n2050 ) ? ( VREG_24_8 ) : ( n2834 ) ;
assign n2836 =  ( n2049 ) ? ( VREG_24_9 ) : ( n2835 ) ;
assign n2837 =  ( n2048 ) ? ( VREG_24_10 ) : ( n2836 ) ;
assign n2838 =  ( n2047 ) ? ( VREG_24_11 ) : ( n2837 ) ;
assign n2839 =  ( n2046 ) ? ( VREG_24_12 ) : ( n2838 ) ;
assign n2840 =  ( n2045 ) ? ( VREG_24_13 ) : ( n2839 ) ;
assign n2841 =  ( n2044 ) ? ( VREG_24_14 ) : ( n2840 ) ;
assign n2842 =  ( n2043 ) ? ( VREG_24_15 ) : ( n2841 ) ;
assign n2843 =  ( n2042 ) ? ( VREG_25_0 ) : ( n2842 ) ;
assign n2844 =  ( n2041 ) ? ( VREG_25_1 ) : ( n2843 ) ;
assign n2845 =  ( n2040 ) ? ( VREG_25_2 ) : ( n2844 ) ;
assign n2846 =  ( n2039 ) ? ( VREG_25_3 ) : ( n2845 ) ;
assign n2847 =  ( n2038 ) ? ( VREG_25_4 ) : ( n2846 ) ;
assign n2848 =  ( n2037 ) ? ( VREG_25_5 ) : ( n2847 ) ;
assign n2849 =  ( n2036 ) ? ( VREG_25_6 ) : ( n2848 ) ;
assign n2850 =  ( n2035 ) ? ( VREG_25_7 ) : ( n2849 ) ;
assign n2851 =  ( n2034 ) ? ( VREG_25_8 ) : ( n2850 ) ;
assign n2852 =  ( n2033 ) ? ( VREG_25_9 ) : ( n2851 ) ;
assign n2853 =  ( n2032 ) ? ( VREG_25_10 ) : ( n2852 ) ;
assign n2854 =  ( n2031 ) ? ( VREG_25_11 ) : ( n2853 ) ;
assign n2855 =  ( n2030 ) ? ( VREG_25_12 ) : ( n2854 ) ;
assign n2856 =  ( n2029 ) ? ( VREG_25_13 ) : ( n2855 ) ;
assign n2857 =  ( n2028 ) ? ( VREG_25_14 ) : ( n2856 ) ;
assign n2858 =  ( n2027 ) ? ( VREG_25_15 ) : ( n2857 ) ;
assign n2859 =  ( n2026 ) ? ( VREG_26_0 ) : ( n2858 ) ;
assign n2860 =  ( n2025 ) ? ( VREG_26_1 ) : ( n2859 ) ;
assign n2861 =  ( n2024 ) ? ( VREG_26_2 ) : ( n2860 ) ;
assign n2862 =  ( n2023 ) ? ( VREG_26_3 ) : ( n2861 ) ;
assign n2863 =  ( n2022 ) ? ( VREG_26_4 ) : ( n2862 ) ;
assign n2864 =  ( n2021 ) ? ( VREG_26_5 ) : ( n2863 ) ;
assign n2865 =  ( n2020 ) ? ( VREG_26_6 ) : ( n2864 ) ;
assign n2866 =  ( n2019 ) ? ( VREG_26_7 ) : ( n2865 ) ;
assign n2867 =  ( n2018 ) ? ( VREG_26_8 ) : ( n2866 ) ;
assign n2868 =  ( n2017 ) ? ( VREG_26_9 ) : ( n2867 ) ;
assign n2869 =  ( n2016 ) ? ( VREG_26_10 ) : ( n2868 ) ;
assign n2870 =  ( n2015 ) ? ( VREG_26_11 ) : ( n2869 ) ;
assign n2871 =  ( n2014 ) ? ( VREG_26_12 ) : ( n2870 ) ;
assign n2872 =  ( n2013 ) ? ( VREG_26_13 ) : ( n2871 ) ;
assign n2873 =  ( n2012 ) ? ( VREG_26_14 ) : ( n2872 ) ;
assign n2874 =  ( n2011 ) ? ( VREG_26_15 ) : ( n2873 ) ;
assign n2875 =  ( n2010 ) ? ( VREG_27_0 ) : ( n2874 ) ;
assign n2876 =  ( n2009 ) ? ( VREG_27_1 ) : ( n2875 ) ;
assign n2877 =  ( n2008 ) ? ( VREG_27_2 ) : ( n2876 ) ;
assign n2878 =  ( n2007 ) ? ( VREG_27_3 ) : ( n2877 ) ;
assign n2879 =  ( n2006 ) ? ( VREG_27_4 ) : ( n2878 ) ;
assign n2880 =  ( n2005 ) ? ( VREG_27_5 ) : ( n2879 ) ;
assign n2881 =  ( n2004 ) ? ( VREG_27_6 ) : ( n2880 ) ;
assign n2882 =  ( n2003 ) ? ( VREG_27_7 ) : ( n2881 ) ;
assign n2883 =  ( n2002 ) ? ( VREG_27_8 ) : ( n2882 ) ;
assign n2884 =  ( n2001 ) ? ( VREG_27_9 ) : ( n2883 ) ;
assign n2885 =  ( n2000 ) ? ( VREG_27_10 ) : ( n2884 ) ;
assign n2886 =  ( n1999 ) ? ( VREG_27_11 ) : ( n2885 ) ;
assign n2887 =  ( n1998 ) ? ( VREG_27_12 ) : ( n2886 ) ;
assign n2888 =  ( n1997 ) ? ( VREG_27_13 ) : ( n2887 ) ;
assign n2889 =  ( n1996 ) ? ( VREG_27_14 ) : ( n2888 ) ;
assign n2890 =  ( n1995 ) ? ( VREG_27_15 ) : ( n2889 ) ;
assign n2891 =  ( n1994 ) ? ( VREG_28_0 ) : ( n2890 ) ;
assign n2892 =  ( n1993 ) ? ( VREG_28_1 ) : ( n2891 ) ;
assign n2893 =  ( n1992 ) ? ( VREG_28_2 ) : ( n2892 ) ;
assign n2894 =  ( n1991 ) ? ( VREG_28_3 ) : ( n2893 ) ;
assign n2895 =  ( n1990 ) ? ( VREG_28_4 ) : ( n2894 ) ;
assign n2896 =  ( n1989 ) ? ( VREG_28_5 ) : ( n2895 ) ;
assign n2897 =  ( n1988 ) ? ( VREG_28_6 ) : ( n2896 ) ;
assign n2898 =  ( n1987 ) ? ( VREG_28_7 ) : ( n2897 ) ;
assign n2899 =  ( n1986 ) ? ( VREG_28_8 ) : ( n2898 ) ;
assign n2900 =  ( n1985 ) ? ( VREG_28_9 ) : ( n2899 ) ;
assign n2901 =  ( n1984 ) ? ( VREG_28_10 ) : ( n2900 ) ;
assign n2902 =  ( n1983 ) ? ( VREG_28_11 ) : ( n2901 ) ;
assign n2903 =  ( n1982 ) ? ( VREG_28_12 ) : ( n2902 ) ;
assign n2904 =  ( n1981 ) ? ( VREG_28_13 ) : ( n2903 ) ;
assign n2905 =  ( n1980 ) ? ( VREG_28_14 ) : ( n2904 ) ;
assign n2906 =  ( n1979 ) ? ( VREG_28_15 ) : ( n2905 ) ;
assign n2907 =  ( n1978 ) ? ( VREG_29_0 ) : ( n2906 ) ;
assign n2908 =  ( n1977 ) ? ( VREG_29_1 ) : ( n2907 ) ;
assign n2909 =  ( n1976 ) ? ( VREG_29_2 ) : ( n2908 ) ;
assign n2910 =  ( n1975 ) ? ( VREG_29_3 ) : ( n2909 ) ;
assign n2911 =  ( n1974 ) ? ( VREG_29_4 ) : ( n2910 ) ;
assign n2912 =  ( n1973 ) ? ( VREG_29_5 ) : ( n2911 ) ;
assign n2913 =  ( n1972 ) ? ( VREG_29_6 ) : ( n2912 ) ;
assign n2914 =  ( n1971 ) ? ( VREG_29_7 ) : ( n2913 ) ;
assign n2915 =  ( n1970 ) ? ( VREG_29_8 ) : ( n2914 ) ;
assign n2916 =  ( n1969 ) ? ( VREG_29_9 ) : ( n2915 ) ;
assign n2917 =  ( n1968 ) ? ( VREG_29_10 ) : ( n2916 ) ;
assign n2918 =  ( n1967 ) ? ( VREG_29_11 ) : ( n2917 ) ;
assign n2919 =  ( n1966 ) ? ( VREG_29_12 ) : ( n2918 ) ;
assign n2920 =  ( n1965 ) ? ( VREG_29_13 ) : ( n2919 ) ;
assign n2921 =  ( n1964 ) ? ( VREG_29_14 ) : ( n2920 ) ;
assign n2922 =  ( n1963 ) ? ( VREG_29_15 ) : ( n2921 ) ;
assign n2923 =  ( n1962 ) ? ( VREG_30_0 ) : ( n2922 ) ;
assign n2924 =  ( n1961 ) ? ( VREG_30_1 ) : ( n2923 ) ;
assign n2925 =  ( n1960 ) ? ( VREG_30_2 ) : ( n2924 ) ;
assign n2926 =  ( n1959 ) ? ( VREG_30_3 ) : ( n2925 ) ;
assign n2927 =  ( n1958 ) ? ( VREG_30_4 ) : ( n2926 ) ;
assign n2928 =  ( n1957 ) ? ( VREG_30_5 ) : ( n2927 ) ;
assign n2929 =  ( n1956 ) ? ( VREG_30_6 ) : ( n2928 ) ;
assign n2930 =  ( n1955 ) ? ( VREG_30_7 ) : ( n2929 ) ;
assign n2931 =  ( n1954 ) ? ( VREG_30_8 ) : ( n2930 ) ;
assign n2932 =  ( n1953 ) ? ( VREG_30_9 ) : ( n2931 ) ;
assign n2933 =  ( n1952 ) ? ( VREG_30_10 ) : ( n2932 ) ;
assign n2934 =  ( n1951 ) ? ( VREG_30_11 ) : ( n2933 ) ;
assign n2935 =  ( n1950 ) ? ( VREG_30_12 ) : ( n2934 ) ;
assign n2936 =  ( n1949 ) ? ( VREG_30_13 ) : ( n2935 ) ;
assign n2937 =  ( n1948 ) ? ( VREG_30_14 ) : ( n2936 ) ;
assign n2938 =  ( n1947 ) ? ( VREG_30_15 ) : ( n2937 ) ;
assign n2939 =  ( n1946 ) ? ( VREG_31_0 ) : ( n2938 ) ;
assign n2940 =  ( n1945 ) ? ( VREG_31_1 ) : ( n2939 ) ;
assign n2941 =  ( n1944 ) ? ( VREG_31_2 ) : ( n2940 ) ;
assign n2942 =  ( n1943 ) ? ( VREG_31_3 ) : ( n2941 ) ;
assign n2943 =  ( n1942 ) ? ( VREG_31_4 ) : ( n2942 ) ;
assign n2944 =  ( n1941 ) ? ( VREG_31_5 ) : ( n2943 ) ;
assign n2945 =  ( n1940 ) ? ( VREG_31_6 ) : ( n2944 ) ;
assign n2946 =  ( n1939 ) ? ( VREG_31_7 ) : ( n2945 ) ;
assign n2947 =  ( n1938 ) ? ( VREG_31_8 ) : ( n2946 ) ;
assign n2948 =  ( n1937 ) ? ( VREG_31_9 ) : ( n2947 ) ;
assign n2949 =  ( n1936 ) ? ( VREG_31_10 ) : ( n2948 ) ;
assign n2950 =  ( n1935 ) ? ( VREG_31_11 ) : ( n2949 ) ;
assign n2951 =  ( n1934 ) ? ( VREG_31_12 ) : ( n2950 ) ;
assign n2952 =  ( n1933 ) ? ( VREG_31_13 ) : ( n2951 ) ;
assign n2953 =  ( n1932 ) ? ( VREG_31_14 ) : ( n2952 ) ;
assign n2954 =  ( n1931 ) ? ( VREG_31_15 ) : ( n2953 ) ;
assign n2955 =  ( n1919 ) + ( n2954 )  ;
assign n2956 =  ( n1919 ) - ( n2954 )  ;
assign n2957 =  ( n1919 ) & ( n2954 )  ;
assign n2958 =  ( n1919 ) | ( n2954 )  ;
assign n2959 =  ( ( n1919 ) * ( n2954 ))  ;
assign n2960 =  ( n148 ) ? ( n2959 ) : ( VREG_0_0 ) ;
assign n2961 =  ( n146 ) ? ( n2958 ) : ( n2960 ) ;
assign n2962 =  ( n144 ) ? ( n2957 ) : ( n2961 ) ;
assign n2963 =  ( n142 ) ? ( n2956 ) : ( n2962 ) ;
assign n2964 =  ( n10 ) ? ( n2955 ) : ( n2963 ) ;
assign n2965 =  ( n7 ) == ( 3'd2 )  ;
assign n2966 = n2[14:10] ;
assign n2967 =  ( n2966 ) == ( 5'd31 )  ;
assign n2968 =  ( n2966 ) == ( 5'd30 )  ;
assign n2969 =  ( n2966 ) == ( 5'd29 )  ;
assign n2970 =  ( n2966 ) == ( 5'd28 )  ;
assign n2971 =  ( n2966 ) == ( 5'd27 )  ;
assign n2972 =  ( n2966 ) == ( 5'd26 )  ;
assign n2973 =  ( n2966 ) == ( 5'd25 )  ;
assign n2974 =  ( n2966 ) == ( 5'd24 )  ;
assign n2975 =  ( n2966 ) == ( 5'd23 )  ;
assign n2976 =  ( n2966 ) == ( 5'd22 )  ;
assign n2977 =  ( n2966 ) == ( 5'd21 )  ;
assign n2978 =  ( n2966 ) == ( 5'd20 )  ;
assign n2979 =  ( n2966 ) == ( 5'd19 )  ;
assign n2980 =  ( n2966 ) == ( 5'd18 )  ;
assign n2981 =  ( n2966 ) == ( 5'd17 )  ;
assign n2982 =  ( n2966 ) == ( 5'd16 )  ;
assign n2983 =  ( n2966 ) == ( 5'd15 )  ;
assign n2984 =  ( n2966 ) == ( 5'd14 )  ;
assign n2985 =  ( n2966 ) == ( 5'd13 )  ;
assign n2986 =  ( n2966 ) == ( 5'd12 )  ;
assign n2987 =  ( n2966 ) == ( 5'd11 )  ;
assign n2988 =  ( n2966 ) == ( 5'd10 )  ;
assign n2989 =  ( n2966 ) == ( 5'd9 )  ;
assign n2990 =  ( n2966 ) == ( 5'd8 )  ;
assign n2991 =  ( n2966 ) == ( 5'd7 )  ;
assign n2992 =  ( n2966 ) == ( 5'd6 )  ;
assign n2993 =  ( n2966 ) == ( 5'd5 )  ;
assign n2994 =  ( n2966 ) == ( 5'd4 )  ;
assign n2995 =  ( n2966 ) == ( 5'd3 )  ;
assign n2996 =  ( n2966 ) == ( 5'd2 )  ;
assign n2997 =  ( n2966 ) == ( 5'd1 )  ;
assign n2998 =  ( n2966 ) == ( 5'd0 )  ;
assign n2999 =  ( n2998 ) ? ( SREG_0 ) : ( SREG_0 ) ;
assign n3000 =  ( n2997 ) ? ( SREG_1 ) : ( n2999 ) ;
assign n3001 =  ( n2996 ) ? ( SREG_2 ) : ( n3000 ) ;
assign n3002 =  ( n2995 ) ? ( SREG_3 ) : ( n3001 ) ;
assign n3003 =  ( n2994 ) ? ( SREG_4 ) : ( n3002 ) ;
assign n3004 =  ( n2993 ) ? ( SREG_5 ) : ( n3003 ) ;
assign n3005 =  ( n2992 ) ? ( SREG_6 ) : ( n3004 ) ;
assign n3006 =  ( n2991 ) ? ( SREG_7 ) : ( n3005 ) ;
assign n3007 =  ( n2990 ) ? ( SREG_8 ) : ( n3006 ) ;
assign n3008 =  ( n2989 ) ? ( SREG_9 ) : ( n3007 ) ;
assign n3009 =  ( n2988 ) ? ( SREG_10 ) : ( n3008 ) ;
assign n3010 =  ( n2987 ) ? ( SREG_11 ) : ( n3009 ) ;
assign n3011 =  ( n2986 ) ? ( SREG_12 ) : ( n3010 ) ;
assign n3012 =  ( n2985 ) ? ( SREG_13 ) : ( n3011 ) ;
assign n3013 =  ( n2984 ) ? ( SREG_14 ) : ( n3012 ) ;
assign n3014 =  ( n2983 ) ? ( SREG_15 ) : ( n3013 ) ;
assign n3015 =  ( n2982 ) ? ( SREG_16 ) : ( n3014 ) ;
assign n3016 =  ( n2981 ) ? ( SREG_17 ) : ( n3015 ) ;
assign n3017 =  ( n2980 ) ? ( SREG_18 ) : ( n3016 ) ;
assign n3018 =  ( n2979 ) ? ( SREG_19 ) : ( n3017 ) ;
assign n3019 =  ( n2978 ) ? ( SREG_20 ) : ( n3018 ) ;
assign n3020 =  ( n2977 ) ? ( SREG_21 ) : ( n3019 ) ;
assign n3021 =  ( n2976 ) ? ( SREG_22 ) : ( n3020 ) ;
assign n3022 =  ( n2975 ) ? ( SREG_23 ) : ( n3021 ) ;
assign n3023 =  ( n2974 ) ? ( SREG_24 ) : ( n3022 ) ;
assign n3024 =  ( n2973 ) ? ( SREG_25 ) : ( n3023 ) ;
assign n3025 =  ( n2972 ) ? ( SREG_26 ) : ( n3024 ) ;
assign n3026 =  ( n2971 ) ? ( SREG_27 ) : ( n3025 ) ;
assign n3027 =  ( n2970 ) ? ( SREG_28 ) : ( n3026 ) ;
assign n3028 =  ( n2969 ) ? ( SREG_29 ) : ( n3027 ) ;
assign n3029 =  ( n2968 ) ? ( SREG_30 ) : ( n3028 ) ;
assign n3030 =  ( n2967 ) ? ( SREG_31 ) : ( n3029 ) ;
assign n3031 = n3030[0:0] ;
assign n3032 =  ( n3031 ) == ( 1'd0 )  ;
assign n3033 =  ( n3032 ) ? ( VREG_0_0 ) : ( n1929 ) ;
assign n3034 =  ( n7 ) == ( 3'd5 )  ;
assign n3035 =  ( n3032 ) ? ( VREG_0_0 ) : ( n2964 ) ;
assign n3036 =  ( n3034 ) ? ( n3035 ) : ( VREG_0_0 ) ;
assign n3037 =  ( n2965 ) ? ( n3033 ) : ( n3036 ) ;
assign n3038 =  ( n1930 ) ? ( n2964 ) : ( n3037 ) ;
assign n3039 =  ( n879 ) ? ( n1929 ) : ( n3038 ) ;
assign n3040 =  ( n158 ) == ( 2'd1 )  ;
assign n3041 =  ( n1919 ) + ( n164 )  ;
assign n3042 =  ( n1919 ) - ( n164 )  ;
assign n3043 =  ( n1919 ) & ( n164 )  ;
assign n3044 =  ( n1919 ) | ( n164 )  ;
assign n3045 =  ( ( n1919 ) * ( n164 ))  ;
assign n3046 =  ( n172 ) ? ( n3045 ) : ( VREG_0_0 ) ;
assign n3047 =  ( n170 ) ? ( n3044 ) : ( n3046 ) ;
assign n3048 =  ( n168 ) ? ( n3043 ) : ( n3047 ) ;
assign n3049 =  ( n166 ) ? ( n3042 ) : ( n3048 ) ;
assign n3050 =  ( n162 ) ? ( n3041 ) : ( n3049 ) ;
assign n3051 =  ( n158 ) == ( 2'd3 )  ;
assign n3052 =  ( n1919 ) + ( n180 )  ;
assign n3053 =  ( n1919 ) - ( n180 )  ;
assign n3054 =  ( n1919 ) & ( n180 )  ;
assign n3055 =  ( n1919 ) | ( n180 )  ;
assign n3056 =  ( ( n1919 ) * ( n180 ))  ;
assign n3057 =  ( n172 ) ? ( n3056 ) : ( VREG_0_0 ) ;
assign n3058 =  ( n170 ) ? ( n3055 ) : ( n3057 ) ;
assign n3059 =  ( n168 ) ? ( n3054 ) : ( n3058 ) ;
assign n3060 =  ( n166 ) ? ( n3053 ) : ( n3059 ) ;
assign n3061 =  ( n162 ) ? ( n3052 ) : ( n3060 ) ;
assign n3062 =  ( n3032 ) ? ( VREG_0_0 ) : ( n3061 ) ;
assign n3063 =  ( n3051 ) ? ( n3062 ) : ( VREG_0_0 ) ;
assign n3064 =  ( n3040 ) ? ( n3050 ) : ( n3063 ) ;
assign n3065 =  ( n192 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n3066 =  ( n157 ) ? ( n3064 ) : ( n3065 ) ;
assign n3067 =  ( n6 ) ? ( n3039 ) : ( n3066 ) ;
assign n3068 =  ( n4 ) ? ( n3067 ) : ( VREG_0_0 ) ;
assign n3069 =  ( 32'd1 ) == ( 32'd15 )  ;
assign n3070 =  ( n12 ) & ( n3069 )  ;
assign n3071 =  ( 32'd1 ) == ( 32'd14 )  ;
assign n3072 =  ( n12 ) & ( n3071 )  ;
assign n3073 =  ( 32'd1 ) == ( 32'd13 )  ;
assign n3074 =  ( n12 ) & ( n3073 )  ;
assign n3075 =  ( 32'd1 ) == ( 32'd12 )  ;
assign n3076 =  ( n12 ) & ( n3075 )  ;
assign n3077 =  ( 32'd1 ) == ( 32'd11 )  ;
assign n3078 =  ( n12 ) & ( n3077 )  ;
assign n3079 =  ( 32'd1 ) == ( 32'd10 )  ;
assign n3080 =  ( n12 ) & ( n3079 )  ;
assign n3081 =  ( 32'd1 ) == ( 32'd9 )  ;
assign n3082 =  ( n12 ) & ( n3081 )  ;
assign n3083 =  ( 32'd1 ) == ( 32'd8 )  ;
assign n3084 =  ( n12 ) & ( n3083 )  ;
assign n3085 =  ( 32'd1 ) == ( 32'd7 )  ;
assign n3086 =  ( n12 ) & ( n3085 )  ;
assign n3087 =  ( 32'd1 ) == ( 32'd6 )  ;
assign n3088 =  ( n12 ) & ( n3087 )  ;
assign n3089 =  ( 32'd1 ) == ( 32'd5 )  ;
assign n3090 =  ( n12 ) & ( n3089 )  ;
assign n3091 =  ( 32'd1 ) == ( 32'd4 )  ;
assign n3092 =  ( n12 ) & ( n3091 )  ;
assign n3093 =  ( 32'd1 ) == ( 32'd3 )  ;
assign n3094 =  ( n12 ) & ( n3093 )  ;
assign n3095 =  ( 32'd1 ) == ( 32'd2 )  ;
assign n3096 =  ( n12 ) & ( n3095 )  ;
assign n3097 =  ( 32'd1 ) == ( 32'd1 )  ;
assign n3098 =  ( n12 ) & ( n3097 )  ;
assign n3099 =  ( 32'd1 ) == ( 32'd0 )  ;
assign n3100 =  ( n12 ) & ( n3099 )  ;
assign n3101 =  ( n13 ) & ( n3069 )  ;
assign n3102 =  ( n13 ) & ( n3071 )  ;
assign n3103 =  ( n13 ) & ( n3073 )  ;
assign n3104 =  ( n13 ) & ( n3075 )  ;
assign n3105 =  ( n13 ) & ( n3077 )  ;
assign n3106 =  ( n13 ) & ( n3079 )  ;
assign n3107 =  ( n13 ) & ( n3081 )  ;
assign n3108 =  ( n13 ) & ( n3083 )  ;
assign n3109 =  ( n13 ) & ( n3085 )  ;
assign n3110 =  ( n13 ) & ( n3087 )  ;
assign n3111 =  ( n13 ) & ( n3089 )  ;
assign n3112 =  ( n13 ) & ( n3091 )  ;
assign n3113 =  ( n13 ) & ( n3093 )  ;
assign n3114 =  ( n13 ) & ( n3095 )  ;
assign n3115 =  ( n13 ) & ( n3097 )  ;
assign n3116 =  ( n13 ) & ( n3099 )  ;
assign n3117 =  ( n14 ) & ( n3069 )  ;
assign n3118 =  ( n14 ) & ( n3071 )  ;
assign n3119 =  ( n14 ) & ( n3073 )  ;
assign n3120 =  ( n14 ) & ( n3075 )  ;
assign n3121 =  ( n14 ) & ( n3077 )  ;
assign n3122 =  ( n14 ) & ( n3079 )  ;
assign n3123 =  ( n14 ) & ( n3081 )  ;
assign n3124 =  ( n14 ) & ( n3083 )  ;
assign n3125 =  ( n14 ) & ( n3085 )  ;
assign n3126 =  ( n14 ) & ( n3087 )  ;
assign n3127 =  ( n14 ) & ( n3089 )  ;
assign n3128 =  ( n14 ) & ( n3091 )  ;
assign n3129 =  ( n14 ) & ( n3093 )  ;
assign n3130 =  ( n14 ) & ( n3095 )  ;
assign n3131 =  ( n14 ) & ( n3097 )  ;
assign n3132 =  ( n14 ) & ( n3099 )  ;
assign n3133 =  ( n15 ) & ( n3069 )  ;
assign n3134 =  ( n15 ) & ( n3071 )  ;
assign n3135 =  ( n15 ) & ( n3073 )  ;
assign n3136 =  ( n15 ) & ( n3075 )  ;
assign n3137 =  ( n15 ) & ( n3077 )  ;
assign n3138 =  ( n15 ) & ( n3079 )  ;
assign n3139 =  ( n15 ) & ( n3081 )  ;
assign n3140 =  ( n15 ) & ( n3083 )  ;
assign n3141 =  ( n15 ) & ( n3085 )  ;
assign n3142 =  ( n15 ) & ( n3087 )  ;
assign n3143 =  ( n15 ) & ( n3089 )  ;
assign n3144 =  ( n15 ) & ( n3091 )  ;
assign n3145 =  ( n15 ) & ( n3093 )  ;
assign n3146 =  ( n15 ) & ( n3095 )  ;
assign n3147 =  ( n15 ) & ( n3097 )  ;
assign n3148 =  ( n15 ) & ( n3099 )  ;
assign n3149 =  ( n16 ) & ( n3069 )  ;
assign n3150 =  ( n16 ) & ( n3071 )  ;
assign n3151 =  ( n16 ) & ( n3073 )  ;
assign n3152 =  ( n16 ) & ( n3075 )  ;
assign n3153 =  ( n16 ) & ( n3077 )  ;
assign n3154 =  ( n16 ) & ( n3079 )  ;
assign n3155 =  ( n16 ) & ( n3081 )  ;
assign n3156 =  ( n16 ) & ( n3083 )  ;
assign n3157 =  ( n16 ) & ( n3085 )  ;
assign n3158 =  ( n16 ) & ( n3087 )  ;
assign n3159 =  ( n16 ) & ( n3089 )  ;
assign n3160 =  ( n16 ) & ( n3091 )  ;
assign n3161 =  ( n16 ) & ( n3093 )  ;
assign n3162 =  ( n16 ) & ( n3095 )  ;
assign n3163 =  ( n16 ) & ( n3097 )  ;
assign n3164 =  ( n16 ) & ( n3099 )  ;
assign n3165 =  ( n17 ) & ( n3069 )  ;
assign n3166 =  ( n17 ) & ( n3071 )  ;
assign n3167 =  ( n17 ) & ( n3073 )  ;
assign n3168 =  ( n17 ) & ( n3075 )  ;
assign n3169 =  ( n17 ) & ( n3077 )  ;
assign n3170 =  ( n17 ) & ( n3079 )  ;
assign n3171 =  ( n17 ) & ( n3081 )  ;
assign n3172 =  ( n17 ) & ( n3083 )  ;
assign n3173 =  ( n17 ) & ( n3085 )  ;
assign n3174 =  ( n17 ) & ( n3087 )  ;
assign n3175 =  ( n17 ) & ( n3089 )  ;
assign n3176 =  ( n17 ) & ( n3091 )  ;
assign n3177 =  ( n17 ) & ( n3093 )  ;
assign n3178 =  ( n17 ) & ( n3095 )  ;
assign n3179 =  ( n17 ) & ( n3097 )  ;
assign n3180 =  ( n17 ) & ( n3099 )  ;
assign n3181 =  ( n18 ) & ( n3069 )  ;
assign n3182 =  ( n18 ) & ( n3071 )  ;
assign n3183 =  ( n18 ) & ( n3073 )  ;
assign n3184 =  ( n18 ) & ( n3075 )  ;
assign n3185 =  ( n18 ) & ( n3077 )  ;
assign n3186 =  ( n18 ) & ( n3079 )  ;
assign n3187 =  ( n18 ) & ( n3081 )  ;
assign n3188 =  ( n18 ) & ( n3083 )  ;
assign n3189 =  ( n18 ) & ( n3085 )  ;
assign n3190 =  ( n18 ) & ( n3087 )  ;
assign n3191 =  ( n18 ) & ( n3089 )  ;
assign n3192 =  ( n18 ) & ( n3091 )  ;
assign n3193 =  ( n18 ) & ( n3093 )  ;
assign n3194 =  ( n18 ) & ( n3095 )  ;
assign n3195 =  ( n18 ) & ( n3097 )  ;
assign n3196 =  ( n18 ) & ( n3099 )  ;
assign n3197 =  ( n19 ) & ( n3069 )  ;
assign n3198 =  ( n19 ) & ( n3071 )  ;
assign n3199 =  ( n19 ) & ( n3073 )  ;
assign n3200 =  ( n19 ) & ( n3075 )  ;
assign n3201 =  ( n19 ) & ( n3077 )  ;
assign n3202 =  ( n19 ) & ( n3079 )  ;
assign n3203 =  ( n19 ) & ( n3081 )  ;
assign n3204 =  ( n19 ) & ( n3083 )  ;
assign n3205 =  ( n19 ) & ( n3085 )  ;
assign n3206 =  ( n19 ) & ( n3087 )  ;
assign n3207 =  ( n19 ) & ( n3089 )  ;
assign n3208 =  ( n19 ) & ( n3091 )  ;
assign n3209 =  ( n19 ) & ( n3093 )  ;
assign n3210 =  ( n19 ) & ( n3095 )  ;
assign n3211 =  ( n19 ) & ( n3097 )  ;
assign n3212 =  ( n19 ) & ( n3099 )  ;
assign n3213 =  ( n20 ) & ( n3069 )  ;
assign n3214 =  ( n20 ) & ( n3071 )  ;
assign n3215 =  ( n20 ) & ( n3073 )  ;
assign n3216 =  ( n20 ) & ( n3075 )  ;
assign n3217 =  ( n20 ) & ( n3077 )  ;
assign n3218 =  ( n20 ) & ( n3079 )  ;
assign n3219 =  ( n20 ) & ( n3081 )  ;
assign n3220 =  ( n20 ) & ( n3083 )  ;
assign n3221 =  ( n20 ) & ( n3085 )  ;
assign n3222 =  ( n20 ) & ( n3087 )  ;
assign n3223 =  ( n20 ) & ( n3089 )  ;
assign n3224 =  ( n20 ) & ( n3091 )  ;
assign n3225 =  ( n20 ) & ( n3093 )  ;
assign n3226 =  ( n20 ) & ( n3095 )  ;
assign n3227 =  ( n20 ) & ( n3097 )  ;
assign n3228 =  ( n20 ) & ( n3099 )  ;
assign n3229 =  ( n21 ) & ( n3069 )  ;
assign n3230 =  ( n21 ) & ( n3071 )  ;
assign n3231 =  ( n21 ) & ( n3073 )  ;
assign n3232 =  ( n21 ) & ( n3075 )  ;
assign n3233 =  ( n21 ) & ( n3077 )  ;
assign n3234 =  ( n21 ) & ( n3079 )  ;
assign n3235 =  ( n21 ) & ( n3081 )  ;
assign n3236 =  ( n21 ) & ( n3083 )  ;
assign n3237 =  ( n21 ) & ( n3085 )  ;
assign n3238 =  ( n21 ) & ( n3087 )  ;
assign n3239 =  ( n21 ) & ( n3089 )  ;
assign n3240 =  ( n21 ) & ( n3091 )  ;
assign n3241 =  ( n21 ) & ( n3093 )  ;
assign n3242 =  ( n21 ) & ( n3095 )  ;
assign n3243 =  ( n21 ) & ( n3097 )  ;
assign n3244 =  ( n21 ) & ( n3099 )  ;
assign n3245 =  ( n22 ) & ( n3069 )  ;
assign n3246 =  ( n22 ) & ( n3071 )  ;
assign n3247 =  ( n22 ) & ( n3073 )  ;
assign n3248 =  ( n22 ) & ( n3075 )  ;
assign n3249 =  ( n22 ) & ( n3077 )  ;
assign n3250 =  ( n22 ) & ( n3079 )  ;
assign n3251 =  ( n22 ) & ( n3081 )  ;
assign n3252 =  ( n22 ) & ( n3083 )  ;
assign n3253 =  ( n22 ) & ( n3085 )  ;
assign n3254 =  ( n22 ) & ( n3087 )  ;
assign n3255 =  ( n22 ) & ( n3089 )  ;
assign n3256 =  ( n22 ) & ( n3091 )  ;
assign n3257 =  ( n22 ) & ( n3093 )  ;
assign n3258 =  ( n22 ) & ( n3095 )  ;
assign n3259 =  ( n22 ) & ( n3097 )  ;
assign n3260 =  ( n22 ) & ( n3099 )  ;
assign n3261 =  ( n23 ) & ( n3069 )  ;
assign n3262 =  ( n23 ) & ( n3071 )  ;
assign n3263 =  ( n23 ) & ( n3073 )  ;
assign n3264 =  ( n23 ) & ( n3075 )  ;
assign n3265 =  ( n23 ) & ( n3077 )  ;
assign n3266 =  ( n23 ) & ( n3079 )  ;
assign n3267 =  ( n23 ) & ( n3081 )  ;
assign n3268 =  ( n23 ) & ( n3083 )  ;
assign n3269 =  ( n23 ) & ( n3085 )  ;
assign n3270 =  ( n23 ) & ( n3087 )  ;
assign n3271 =  ( n23 ) & ( n3089 )  ;
assign n3272 =  ( n23 ) & ( n3091 )  ;
assign n3273 =  ( n23 ) & ( n3093 )  ;
assign n3274 =  ( n23 ) & ( n3095 )  ;
assign n3275 =  ( n23 ) & ( n3097 )  ;
assign n3276 =  ( n23 ) & ( n3099 )  ;
assign n3277 =  ( n24 ) & ( n3069 )  ;
assign n3278 =  ( n24 ) & ( n3071 )  ;
assign n3279 =  ( n24 ) & ( n3073 )  ;
assign n3280 =  ( n24 ) & ( n3075 )  ;
assign n3281 =  ( n24 ) & ( n3077 )  ;
assign n3282 =  ( n24 ) & ( n3079 )  ;
assign n3283 =  ( n24 ) & ( n3081 )  ;
assign n3284 =  ( n24 ) & ( n3083 )  ;
assign n3285 =  ( n24 ) & ( n3085 )  ;
assign n3286 =  ( n24 ) & ( n3087 )  ;
assign n3287 =  ( n24 ) & ( n3089 )  ;
assign n3288 =  ( n24 ) & ( n3091 )  ;
assign n3289 =  ( n24 ) & ( n3093 )  ;
assign n3290 =  ( n24 ) & ( n3095 )  ;
assign n3291 =  ( n24 ) & ( n3097 )  ;
assign n3292 =  ( n24 ) & ( n3099 )  ;
assign n3293 =  ( n25 ) & ( n3069 )  ;
assign n3294 =  ( n25 ) & ( n3071 )  ;
assign n3295 =  ( n25 ) & ( n3073 )  ;
assign n3296 =  ( n25 ) & ( n3075 )  ;
assign n3297 =  ( n25 ) & ( n3077 )  ;
assign n3298 =  ( n25 ) & ( n3079 )  ;
assign n3299 =  ( n25 ) & ( n3081 )  ;
assign n3300 =  ( n25 ) & ( n3083 )  ;
assign n3301 =  ( n25 ) & ( n3085 )  ;
assign n3302 =  ( n25 ) & ( n3087 )  ;
assign n3303 =  ( n25 ) & ( n3089 )  ;
assign n3304 =  ( n25 ) & ( n3091 )  ;
assign n3305 =  ( n25 ) & ( n3093 )  ;
assign n3306 =  ( n25 ) & ( n3095 )  ;
assign n3307 =  ( n25 ) & ( n3097 )  ;
assign n3308 =  ( n25 ) & ( n3099 )  ;
assign n3309 =  ( n26 ) & ( n3069 )  ;
assign n3310 =  ( n26 ) & ( n3071 )  ;
assign n3311 =  ( n26 ) & ( n3073 )  ;
assign n3312 =  ( n26 ) & ( n3075 )  ;
assign n3313 =  ( n26 ) & ( n3077 )  ;
assign n3314 =  ( n26 ) & ( n3079 )  ;
assign n3315 =  ( n26 ) & ( n3081 )  ;
assign n3316 =  ( n26 ) & ( n3083 )  ;
assign n3317 =  ( n26 ) & ( n3085 )  ;
assign n3318 =  ( n26 ) & ( n3087 )  ;
assign n3319 =  ( n26 ) & ( n3089 )  ;
assign n3320 =  ( n26 ) & ( n3091 )  ;
assign n3321 =  ( n26 ) & ( n3093 )  ;
assign n3322 =  ( n26 ) & ( n3095 )  ;
assign n3323 =  ( n26 ) & ( n3097 )  ;
assign n3324 =  ( n26 ) & ( n3099 )  ;
assign n3325 =  ( n27 ) & ( n3069 )  ;
assign n3326 =  ( n27 ) & ( n3071 )  ;
assign n3327 =  ( n27 ) & ( n3073 )  ;
assign n3328 =  ( n27 ) & ( n3075 )  ;
assign n3329 =  ( n27 ) & ( n3077 )  ;
assign n3330 =  ( n27 ) & ( n3079 )  ;
assign n3331 =  ( n27 ) & ( n3081 )  ;
assign n3332 =  ( n27 ) & ( n3083 )  ;
assign n3333 =  ( n27 ) & ( n3085 )  ;
assign n3334 =  ( n27 ) & ( n3087 )  ;
assign n3335 =  ( n27 ) & ( n3089 )  ;
assign n3336 =  ( n27 ) & ( n3091 )  ;
assign n3337 =  ( n27 ) & ( n3093 )  ;
assign n3338 =  ( n27 ) & ( n3095 )  ;
assign n3339 =  ( n27 ) & ( n3097 )  ;
assign n3340 =  ( n27 ) & ( n3099 )  ;
assign n3341 =  ( n28 ) & ( n3069 )  ;
assign n3342 =  ( n28 ) & ( n3071 )  ;
assign n3343 =  ( n28 ) & ( n3073 )  ;
assign n3344 =  ( n28 ) & ( n3075 )  ;
assign n3345 =  ( n28 ) & ( n3077 )  ;
assign n3346 =  ( n28 ) & ( n3079 )  ;
assign n3347 =  ( n28 ) & ( n3081 )  ;
assign n3348 =  ( n28 ) & ( n3083 )  ;
assign n3349 =  ( n28 ) & ( n3085 )  ;
assign n3350 =  ( n28 ) & ( n3087 )  ;
assign n3351 =  ( n28 ) & ( n3089 )  ;
assign n3352 =  ( n28 ) & ( n3091 )  ;
assign n3353 =  ( n28 ) & ( n3093 )  ;
assign n3354 =  ( n28 ) & ( n3095 )  ;
assign n3355 =  ( n28 ) & ( n3097 )  ;
assign n3356 =  ( n28 ) & ( n3099 )  ;
assign n3357 =  ( n29 ) & ( n3069 )  ;
assign n3358 =  ( n29 ) & ( n3071 )  ;
assign n3359 =  ( n29 ) & ( n3073 )  ;
assign n3360 =  ( n29 ) & ( n3075 )  ;
assign n3361 =  ( n29 ) & ( n3077 )  ;
assign n3362 =  ( n29 ) & ( n3079 )  ;
assign n3363 =  ( n29 ) & ( n3081 )  ;
assign n3364 =  ( n29 ) & ( n3083 )  ;
assign n3365 =  ( n29 ) & ( n3085 )  ;
assign n3366 =  ( n29 ) & ( n3087 )  ;
assign n3367 =  ( n29 ) & ( n3089 )  ;
assign n3368 =  ( n29 ) & ( n3091 )  ;
assign n3369 =  ( n29 ) & ( n3093 )  ;
assign n3370 =  ( n29 ) & ( n3095 )  ;
assign n3371 =  ( n29 ) & ( n3097 )  ;
assign n3372 =  ( n29 ) & ( n3099 )  ;
assign n3373 =  ( n30 ) & ( n3069 )  ;
assign n3374 =  ( n30 ) & ( n3071 )  ;
assign n3375 =  ( n30 ) & ( n3073 )  ;
assign n3376 =  ( n30 ) & ( n3075 )  ;
assign n3377 =  ( n30 ) & ( n3077 )  ;
assign n3378 =  ( n30 ) & ( n3079 )  ;
assign n3379 =  ( n30 ) & ( n3081 )  ;
assign n3380 =  ( n30 ) & ( n3083 )  ;
assign n3381 =  ( n30 ) & ( n3085 )  ;
assign n3382 =  ( n30 ) & ( n3087 )  ;
assign n3383 =  ( n30 ) & ( n3089 )  ;
assign n3384 =  ( n30 ) & ( n3091 )  ;
assign n3385 =  ( n30 ) & ( n3093 )  ;
assign n3386 =  ( n30 ) & ( n3095 )  ;
assign n3387 =  ( n30 ) & ( n3097 )  ;
assign n3388 =  ( n30 ) & ( n3099 )  ;
assign n3389 =  ( n31 ) & ( n3069 )  ;
assign n3390 =  ( n31 ) & ( n3071 )  ;
assign n3391 =  ( n31 ) & ( n3073 )  ;
assign n3392 =  ( n31 ) & ( n3075 )  ;
assign n3393 =  ( n31 ) & ( n3077 )  ;
assign n3394 =  ( n31 ) & ( n3079 )  ;
assign n3395 =  ( n31 ) & ( n3081 )  ;
assign n3396 =  ( n31 ) & ( n3083 )  ;
assign n3397 =  ( n31 ) & ( n3085 )  ;
assign n3398 =  ( n31 ) & ( n3087 )  ;
assign n3399 =  ( n31 ) & ( n3089 )  ;
assign n3400 =  ( n31 ) & ( n3091 )  ;
assign n3401 =  ( n31 ) & ( n3093 )  ;
assign n3402 =  ( n31 ) & ( n3095 )  ;
assign n3403 =  ( n31 ) & ( n3097 )  ;
assign n3404 =  ( n31 ) & ( n3099 )  ;
assign n3405 =  ( n32 ) & ( n3069 )  ;
assign n3406 =  ( n32 ) & ( n3071 )  ;
assign n3407 =  ( n32 ) & ( n3073 )  ;
assign n3408 =  ( n32 ) & ( n3075 )  ;
assign n3409 =  ( n32 ) & ( n3077 )  ;
assign n3410 =  ( n32 ) & ( n3079 )  ;
assign n3411 =  ( n32 ) & ( n3081 )  ;
assign n3412 =  ( n32 ) & ( n3083 )  ;
assign n3413 =  ( n32 ) & ( n3085 )  ;
assign n3414 =  ( n32 ) & ( n3087 )  ;
assign n3415 =  ( n32 ) & ( n3089 )  ;
assign n3416 =  ( n32 ) & ( n3091 )  ;
assign n3417 =  ( n32 ) & ( n3093 )  ;
assign n3418 =  ( n32 ) & ( n3095 )  ;
assign n3419 =  ( n32 ) & ( n3097 )  ;
assign n3420 =  ( n32 ) & ( n3099 )  ;
assign n3421 =  ( n33 ) & ( n3069 )  ;
assign n3422 =  ( n33 ) & ( n3071 )  ;
assign n3423 =  ( n33 ) & ( n3073 )  ;
assign n3424 =  ( n33 ) & ( n3075 )  ;
assign n3425 =  ( n33 ) & ( n3077 )  ;
assign n3426 =  ( n33 ) & ( n3079 )  ;
assign n3427 =  ( n33 ) & ( n3081 )  ;
assign n3428 =  ( n33 ) & ( n3083 )  ;
assign n3429 =  ( n33 ) & ( n3085 )  ;
assign n3430 =  ( n33 ) & ( n3087 )  ;
assign n3431 =  ( n33 ) & ( n3089 )  ;
assign n3432 =  ( n33 ) & ( n3091 )  ;
assign n3433 =  ( n33 ) & ( n3093 )  ;
assign n3434 =  ( n33 ) & ( n3095 )  ;
assign n3435 =  ( n33 ) & ( n3097 )  ;
assign n3436 =  ( n33 ) & ( n3099 )  ;
assign n3437 =  ( n34 ) & ( n3069 )  ;
assign n3438 =  ( n34 ) & ( n3071 )  ;
assign n3439 =  ( n34 ) & ( n3073 )  ;
assign n3440 =  ( n34 ) & ( n3075 )  ;
assign n3441 =  ( n34 ) & ( n3077 )  ;
assign n3442 =  ( n34 ) & ( n3079 )  ;
assign n3443 =  ( n34 ) & ( n3081 )  ;
assign n3444 =  ( n34 ) & ( n3083 )  ;
assign n3445 =  ( n34 ) & ( n3085 )  ;
assign n3446 =  ( n34 ) & ( n3087 )  ;
assign n3447 =  ( n34 ) & ( n3089 )  ;
assign n3448 =  ( n34 ) & ( n3091 )  ;
assign n3449 =  ( n34 ) & ( n3093 )  ;
assign n3450 =  ( n34 ) & ( n3095 )  ;
assign n3451 =  ( n34 ) & ( n3097 )  ;
assign n3452 =  ( n34 ) & ( n3099 )  ;
assign n3453 =  ( n35 ) & ( n3069 )  ;
assign n3454 =  ( n35 ) & ( n3071 )  ;
assign n3455 =  ( n35 ) & ( n3073 )  ;
assign n3456 =  ( n35 ) & ( n3075 )  ;
assign n3457 =  ( n35 ) & ( n3077 )  ;
assign n3458 =  ( n35 ) & ( n3079 )  ;
assign n3459 =  ( n35 ) & ( n3081 )  ;
assign n3460 =  ( n35 ) & ( n3083 )  ;
assign n3461 =  ( n35 ) & ( n3085 )  ;
assign n3462 =  ( n35 ) & ( n3087 )  ;
assign n3463 =  ( n35 ) & ( n3089 )  ;
assign n3464 =  ( n35 ) & ( n3091 )  ;
assign n3465 =  ( n35 ) & ( n3093 )  ;
assign n3466 =  ( n35 ) & ( n3095 )  ;
assign n3467 =  ( n35 ) & ( n3097 )  ;
assign n3468 =  ( n35 ) & ( n3099 )  ;
assign n3469 =  ( n36 ) & ( n3069 )  ;
assign n3470 =  ( n36 ) & ( n3071 )  ;
assign n3471 =  ( n36 ) & ( n3073 )  ;
assign n3472 =  ( n36 ) & ( n3075 )  ;
assign n3473 =  ( n36 ) & ( n3077 )  ;
assign n3474 =  ( n36 ) & ( n3079 )  ;
assign n3475 =  ( n36 ) & ( n3081 )  ;
assign n3476 =  ( n36 ) & ( n3083 )  ;
assign n3477 =  ( n36 ) & ( n3085 )  ;
assign n3478 =  ( n36 ) & ( n3087 )  ;
assign n3479 =  ( n36 ) & ( n3089 )  ;
assign n3480 =  ( n36 ) & ( n3091 )  ;
assign n3481 =  ( n36 ) & ( n3093 )  ;
assign n3482 =  ( n36 ) & ( n3095 )  ;
assign n3483 =  ( n36 ) & ( n3097 )  ;
assign n3484 =  ( n36 ) & ( n3099 )  ;
assign n3485 =  ( n37 ) & ( n3069 )  ;
assign n3486 =  ( n37 ) & ( n3071 )  ;
assign n3487 =  ( n37 ) & ( n3073 )  ;
assign n3488 =  ( n37 ) & ( n3075 )  ;
assign n3489 =  ( n37 ) & ( n3077 )  ;
assign n3490 =  ( n37 ) & ( n3079 )  ;
assign n3491 =  ( n37 ) & ( n3081 )  ;
assign n3492 =  ( n37 ) & ( n3083 )  ;
assign n3493 =  ( n37 ) & ( n3085 )  ;
assign n3494 =  ( n37 ) & ( n3087 )  ;
assign n3495 =  ( n37 ) & ( n3089 )  ;
assign n3496 =  ( n37 ) & ( n3091 )  ;
assign n3497 =  ( n37 ) & ( n3093 )  ;
assign n3498 =  ( n37 ) & ( n3095 )  ;
assign n3499 =  ( n37 ) & ( n3097 )  ;
assign n3500 =  ( n37 ) & ( n3099 )  ;
assign n3501 =  ( n38 ) & ( n3069 )  ;
assign n3502 =  ( n38 ) & ( n3071 )  ;
assign n3503 =  ( n38 ) & ( n3073 )  ;
assign n3504 =  ( n38 ) & ( n3075 )  ;
assign n3505 =  ( n38 ) & ( n3077 )  ;
assign n3506 =  ( n38 ) & ( n3079 )  ;
assign n3507 =  ( n38 ) & ( n3081 )  ;
assign n3508 =  ( n38 ) & ( n3083 )  ;
assign n3509 =  ( n38 ) & ( n3085 )  ;
assign n3510 =  ( n38 ) & ( n3087 )  ;
assign n3511 =  ( n38 ) & ( n3089 )  ;
assign n3512 =  ( n38 ) & ( n3091 )  ;
assign n3513 =  ( n38 ) & ( n3093 )  ;
assign n3514 =  ( n38 ) & ( n3095 )  ;
assign n3515 =  ( n38 ) & ( n3097 )  ;
assign n3516 =  ( n38 ) & ( n3099 )  ;
assign n3517 =  ( n39 ) & ( n3069 )  ;
assign n3518 =  ( n39 ) & ( n3071 )  ;
assign n3519 =  ( n39 ) & ( n3073 )  ;
assign n3520 =  ( n39 ) & ( n3075 )  ;
assign n3521 =  ( n39 ) & ( n3077 )  ;
assign n3522 =  ( n39 ) & ( n3079 )  ;
assign n3523 =  ( n39 ) & ( n3081 )  ;
assign n3524 =  ( n39 ) & ( n3083 )  ;
assign n3525 =  ( n39 ) & ( n3085 )  ;
assign n3526 =  ( n39 ) & ( n3087 )  ;
assign n3527 =  ( n39 ) & ( n3089 )  ;
assign n3528 =  ( n39 ) & ( n3091 )  ;
assign n3529 =  ( n39 ) & ( n3093 )  ;
assign n3530 =  ( n39 ) & ( n3095 )  ;
assign n3531 =  ( n39 ) & ( n3097 )  ;
assign n3532 =  ( n39 ) & ( n3099 )  ;
assign n3533 =  ( n40 ) & ( n3069 )  ;
assign n3534 =  ( n40 ) & ( n3071 )  ;
assign n3535 =  ( n40 ) & ( n3073 )  ;
assign n3536 =  ( n40 ) & ( n3075 )  ;
assign n3537 =  ( n40 ) & ( n3077 )  ;
assign n3538 =  ( n40 ) & ( n3079 )  ;
assign n3539 =  ( n40 ) & ( n3081 )  ;
assign n3540 =  ( n40 ) & ( n3083 )  ;
assign n3541 =  ( n40 ) & ( n3085 )  ;
assign n3542 =  ( n40 ) & ( n3087 )  ;
assign n3543 =  ( n40 ) & ( n3089 )  ;
assign n3544 =  ( n40 ) & ( n3091 )  ;
assign n3545 =  ( n40 ) & ( n3093 )  ;
assign n3546 =  ( n40 ) & ( n3095 )  ;
assign n3547 =  ( n40 ) & ( n3097 )  ;
assign n3548 =  ( n40 ) & ( n3099 )  ;
assign n3549 =  ( n41 ) & ( n3069 )  ;
assign n3550 =  ( n41 ) & ( n3071 )  ;
assign n3551 =  ( n41 ) & ( n3073 )  ;
assign n3552 =  ( n41 ) & ( n3075 )  ;
assign n3553 =  ( n41 ) & ( n3077 )  ;
assign n3554 =  ( n41 ) & ( n3079 )  ;
assign n3555 =  ( n41 ) & ( n3081 )  ;
assign n3556 =  ( n41 ) & ( n3083 )  ;
assign n3557 =  ( n41 ) & ( n3085 )  ;
assign n3558 =  ( n41 ) & ( n3087 )  ;
assign n3559 =  ( n41 ) & ( n3089 )  ;
assign n3560 =  ( n41 ) & ( n3091 )  ;
assign n3561 =  ( n41 ) & ( n3093 )  ;
assign n3562 =  ( n41 ) & ( n3095 )  ;
assign n3563 =  ( n41 ) & ( n3097 )  ;
assign n3564 =  ( n41 ) & ( n3099 )  ;
assign n3565 =  ( n42 ) & ( n3069 )  ;
assign n3566 =  ( n42 ) & ( n3071 )  ;
assign n3567 =  ( n42 ) & ( n3073 )  ;
assign n3568 =  ( n42 ) & ( n3075 )  ;
assign n3569 =  ( n42 ) & ( n3077 )  ;
assign n3570 =  ( n42 ) & ( n3079 )  ;
assign n3571 =  ( n42 ) & ( n3081 )  ;
assign n3572 =  ( n42 ) & ( n3083 )  ;
assign n3573 =  ( n42 ) & ( n3085 )  ;
assign n3574 =  ( n42 ) & ( n3087 )  ;
assign n3575 =  ( n42 ) & ( n3089 )  ;
assign n3576 =  ( n42 ) & ( n3091 )  ;
assign n3577 =  ( n42 ) & ( n3093 )  ;
assign n3578 =  ( n42 ) & ( n3095 )  ;
assign n3579 =  ( n42 ) & ( n3097 )  ;
assign n3580 =  ( n42 ) & ( n3099 )  ;
assign n3581 =  ( n43 ) & ( n3069 )  ;
assign n3582 =  ( n43 ) & ( n3071 )  ;
assign n3583 =  ( n43 ) & ( n3073 )  ;
assign n3584 =  ( n43 ) & ( n3075 )  ;
assign n3585 =  ( n43 ) & ( n3077 )  ;
assign n3586 =  ( n43 ) & ( n3079 )  ;
assign n3587 =  ( n43 ) & ( n3081 )  ;
assign n3588 =  ( n43 ) & ( n3083 )  ;
assign n3589 =  ( n43 ) & ( n3085 )  ;
assign n3590 =  ( n43 ) & ( n3087 )  ;
assign n3591 =  ( n43 ) & ( n3089 )  ;
assign n3592 =  ( n43 ) & ( n3091 )  ;
assign n3593 =  ( n43 ) & ( n3093 )  ;
assign n3594 =  ( n43 ) & ( n3095 )  ;
assign n3595 =  ( n43 ) & ( n3097 )  ;
assign n3596 =  ( n43 ) & ( n3099 )  ;
assign n3597 =  ( n3596 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n3598 =  ( n3595 ) ? ( VREG_0_1 ) : ( n3597 ) ;
assign n3599 =  ( n3594 ) ? ( VREG_0_2 ) : ( n3598 ) ;
assign n3600 =  ( n3593 ) ? ( VREG_0_3 ) : ( n3599 ) ;
assign n3601 =  ( n3592 ) ? ( VREG_0_4 ) : ( n3600 ) ;
assign n3602 =  ( n3591 ) ? ( VREG_0_5 ) : ( n3601 ) ;
assign n3603 =  ( n3590 ) ? ( VREG_0_6 ) : ( n3602 ) ;
assign n3604 =  ( n3589 ) ? ( VREG_0_7 ) : ( n3603 ) ;
assign n3605 =  ( n3588 ) ? ( VREG_0_8 ) : ( n3604 ) ;
assign n3606 =  ( n3587 ) ? ( VREG_0_9 ) : ( n3605 ) ;
assign n3607 =  ( n3586 ) ? ( VREG_0_10 ) : ( n3606 ) ;
assign n3608 =  ( n3585 ) ? ( VREG_0_11 ) : ( n3607 ) ;
assign n3609 =  ( n3584 ) ? ( VREG_0_12 ) : ( n3608 ) ;
assign n3610 =  ( n3583 ) ? ( VREG_0_13 ) : ( n3609 ) ;
assign n3611 =  ( n3582 ) ? ( VREG_0_14 ) : ( n3610 ) ;
assign n3612 =  ( n3581 ) ? ( VREG_0_15 ) : ( n3611 ) ;
assign n3613 =  ( n3580 ) ? ( VREG_1_0 ) : ( n3612 ) ;
assign n3614 =  ( n3579 ) ? ( VREG_1_1 ) : ( n3613 ) ;
assign n3615 =  ( n3578 ) ? ( VREG_1_2 ) : ( n3614 ) ;
assign n3616 =  ( n3577 ) ? ( VREG_1_3 ) : ( n3615 ) ;
assign n3617 =  ( n3576 ) ? ( VREG_1_4 ) : ( n3616 ) ;
assign n3618 =  ( n3575 ) ? ( VREG_1_5 ) : ( n3617 ) ;
assign n3619 =  ( n3574 ) ? ( VREG_1_6 ) : ( n3618 ) ;
assign n3620 =  ( n3573 ) ? ( VREG_1_7 ) : ( n3619 ) ;
assign n3621 =  ( n3572 ) ? ( VREG_1_8 ) : ( n3620 ) ;
assign n3622 =  ( n3571 ) ? ( VREG_1_9 ) : ( n3621 ) ;
assign n3623 =  ( n3570 ) ? ( VREG_1_10 ) : ( n3622 ) ;
assign n3624 =  ( n3569 ) ? ( VREG_1_11 ) : ( n3623 ) ;
assign n3625 =  ( n3568 ) ? ( VREG_1_12 ) : ( n3624 ) ;
assign n3626 =  ( n3567 ) ? ( VREG_1_13 ) : ( n3625 ) ;
assign n3627 =  ( n3566 ) ? ( VREG_1_14 ) : ( n3626 ) ;
assign n3628 =  ( n3565 ) ? ( VREG_1_15 ) : ( n3627 ) ;
assign n3629 =  ( n3564 ) ? ( VREG_2_0 ) : ( n3628 ) ;
assign n3630 =  ( n3563 ) ? ( VREG_2_1 ) : ( n3629 ) ;
assign n3631 =  ( n3562 ) ? ( VREG_2_2 ) : ( n3630 ) ;
assign n3632 =  ( n3561 ) ? ( VREG_2_3 ) : ( n3631 ) ;
assign n3633 =  ( n3560 ) ? ( VREG_2_4 ) : ( n3632 ) ;
assign n3634 =  ( n3559 ) ? ( VREG_2_5 ) : ( n3633 ) ;
assign n3635 =  ( n3558 ) ? ( VREG_2_6 ) : ( n3634 ) ;
assign n3636 =  ( n3557 ) ? ( VREG_2_7 ) : ( n3635 ) ;
assign n3637 =  ( n3556 ) ? ( VREG_2_8 ) : ( n3636 ) ;
assign n3638 =  ( n3555 ) ? ( VREG_2_9 ) : ( n3637 ) ;
assign n3639 =  ( n3554 ) ? ( VREG_2_10 ) : ( n3638 ) ;
assign n3640 =  ( n3553 ) ? ( VREG_2_11 ) : ( n3639 ) ;
assign n3641 =  ( n3552 ) ? ( VREG_2_12 ) : ( n3640 ) ;
assign n3642 =  ( n3551 ) ? ( VREG_2_13 ) : ( n3641 ) ;
assign n3643 =  ( n3550 ) ? ( VREG_2_14 ) : ( n3642 ) ;
assign n3644 =  ( n3549 ) ? ( VREG_2_15 ) : ( n3643 ) ;
assign n3645 =  ( n3548 ) ? ( VREG_3_0 ) : ( n3644 ) ;
assign n3646 =  ( n3547 ) ? ( VREG_3_1 ) : ( n3645 ) ;
assign n3647 =  ( n3546 ) ? ( VREG_3_2 ) : ( n3646 ) ;
assign n3648 =  ( n3545 ) ? ( VREG_3_3 ) : ( n3647 ) ;
assign n3649 =  ( n3544 ) ? ( VREG_3_4 ) : ( n3648 ) ;
assign n3650 =  ( n3543 ) ? ( VREG_3_5 ) : ( n3649 ) ;
assign n3651 =  ( n3542 ) ? ( VREG_3_6 ) : ( n3650 ) ;
assign n3652 =  ( n3541 ) ? ( VREG_3_7 ) : ( n3651 ) ;
assign n3653 =  ( n3540 ) ? ( VREG_3_8 ) : ( n3652 ) ;
assign n3654 =  ( n3539 ) ? ( VREG_3_9 ) : ( n3653 ) ;
assign n3655 =  ( n3538 ) ? ( VREG_3_10 ) : ( n3654 ) ;
assign n3656 =  ( n3537 ) ? ( VREG_3_11 ) : ( n3655 ) ;
assign n3657 =  ( n3536 ) ? ( VREG_3_12 ) : ( n3656 ) ;
assign n3658 =  ( n3535 ) ? ( VREG_3_13 ) : ( n3657 ) ;
assign n3659 =  ( n3534 ) ? ( VREG_3_14 ) : ( n3658 ) ;
assign n3660 =  ( n3533 ) ? ( VREG_3_15 ) : ( n3659 ) ;
assign n3661 =  ( n3532 ) ? ( VREG_4_0 ) : ( n3660 ) ;
assign n3662 =  ( n3531 ) ? ( VREG_4_1 ) : ( n3661 ) ;
assign n3663 =  ( n3530 ) ? ( VREG_4_2 ) : ( n3662 ) ;
assign n3664 =  ( n3529 ) ? ( VREG_4_3 ) : ( n3663 ) ;
assign n3665 =  ( n3528 ) ? ( VREG_4_4 ) : ( n3664 ) ;
assign n3666 =  ( n3527 ) ? ( VREG_4_5 ) : ( n3665 ) ;
assign n3667 =  ( n3526 ) ? ( VREG_4_6 ) : ( n3666 ) ;
assign n3668 =  ( n3525 ) ? ( VREG_4_7 ) : ( n3667 ) ;
assign n3669 =  ( n3524 ) ? ( VREG_4_8 ) : ( n3668 ) ;
assign n3670 =  ( n3523 ) ? ( VREG_4_9 ) : ( n3669 ) ;
assign n3671 =  ( n3522 ) ? ( VREG_4_10 ) : ( n3670 ) ;
assign n3672 =  ( n3521 ) ? ( VREG_4_11 ) : ( n3671 ) ;
assign n3673 =  ( n3520 ) ? ( VREG_4_12 ) : ( n3672 ) ;
assign n3674 =  ( n3519 ) ? ( VREG_4_13 ) : ( n3673 ) ;
assign n3675 =  ( n3518 ) ? ( VREG_4_14 ) : ( n3674 ) ;
assign n3676 =  ( n3517 ) ? ( VREG_4_15 ) : ( n3675 ) ;
assign n3677 =  ( n3516 ) ? ( VREG_5_0 ) : ( n3676 ) ;
assign n3678 =  ( n3515 ) ? ( VREG_5_1 ) : ( n3677 ) ;
assign n3679 =  ( n3514 ) ? ( VREG_5_2 ) : ( n3678 ) ;
assign n3680 =  ( n3513 ) ? ( VREG_5_3 ) : ( n3679 ) ;
assign n3681 =  ( n3512 ) ? ( VREG_5_4 ) : ( n3680 ) ;
assign n3682 =  ( n3511 ) ? ( VREG_5_5 ) : ( n3681 ) ;
assign n3683 =  ( n3510 ) ? ( VREG_5_6 ) : ( n3682 ) ;
assign n3684 =  ( n3509 ) ? ( VREG_5_7 ) : ( n3683 ) ;
assign n3685 =  ( n3508 ) ? ( VREG_5_8 ) : ( n3684 ) ;
assign n3686 =  ( n3507 ) ? ( VREG_5_9 ) : ( n3685 ) ;
assign n3687 =  ( n3506 ) ? ( VREG_5_10 ) : ( n3686 ) ;
assign n3688 =  ( n3505 ) ? ( VREG_5_11 ) : ( n3687 ) ;
assign n3689 =  ( n3504 ) ? ( VREG_5_12 ) : ( n3688 ) ;
assign n3690 =  ( n3503 ) ? ( VREG_5_13 ) : ( n3689 ) ;
assign n3691 =  ( n3502 ) ? ( VREG_5_14 ) : ( n3690 ) ;
assign n3692 =  ( n3501 ) ? ( VREG_5_15 ) : ( n3691 ) ;
assign n3693 =  ( n3500 ) ? ( VREG_6_0 ) : ( n3692 ) ;
assign n3694 =  ( n3499 ) ? ( VREG_6_1 ) : ( n3693 ) ;
assign n3695 =  ( n3498 ) ? ( VREG_6_2 ) : ( n3694 ) ;
assign n3696 =  ( n3497 ) ? ( VREG_6_3 ) : ( n3695 ) ;
assign n3697 =  ( n3496 ) ? ( VREG_6_4 ) : ( n3696 ) ;
assign n3698 =  ( n3495 ) ? ( VREG_6_5 ) : ( n3697 ) ;
assign n3699 =  ( n3494 ) ? ( VREG_6_6 ) : ( n3698 ) ;
assign n3700 =  ( n3493 ) ? ( VREG_6_7 ) : ( n3699 ) ;
assign n3701 =  ( n3492 ) ? ( VREG_6_8 ) : ( n3700 ) ;
assign n3702 =  ( n3491 ) ? ( VREG_6_9 ) : ( n3701 ) ;
assign n3703 =  ( n3490 ) ? ( VREG_6_10 ) : ( n3702 ) ;
assign n3704 =  ( n3489 ) ? ( VREG_6_11 ) : ( n3703 ) ;
assign n3705 =  ( n3488 ) ? ( VREG_6_12 ) : ( n3704 ) ;
assign n3706 =  ( n3487 ) ? ( VREG_6_13 ) : ( n3705 ) ;
assign n3707 =  ( n3486 ) ? ( VREG_6_14 ) : ( n3706 ) ;
assign n3708 =  ( n3485 ) ? ( VREG_6_15 ) : ( n3707 ) ;
assign n3709 =  ( n3484 ) ? ( VREG_7_0 ) : ( n3708 ) ;
assign n3710 =  ( n3483 ) ? ( VREG_7_1 ) : ( n3709 ) ;
assign n3711 =  ( n3482 ) ? ( VREG_7_2 ) : ( n3710 ) ;
assign n3712 =  ( n3481 ) ? ( VREG_7_3 ) : ( n3711 ) ;
assign n3713 =  ( n3480 ) ? ( VREG_7_4 ) : ( n3712 ) ;
assign n3714 =  ( n3479 ) ? ( VREG_7_5 ) : ( n3713 ) ;
assign n3715 =  ( n3478 ) ? ( VREG_7_6 ) : ( n3714 ) ;
assign n3716 =  ( n3477 ) ? ( VREG_7_7 ) : ( n3715 ) ;
assign n3717 =  ( n3476 ) ? ( VREG_7_8 ) : ( n3716 ) ;
assign n3718 =  ( n3475 ) ? ( VREG_7_9 ) : ( n3717 ) ;
assign n3719 =  ( n3474 ) ? ( VREG_7_10 ) : ( n3718 ) ;
assign n3720 =  ( n3473 ) ? ( VREG_7_11 ) : ( n3719 ) ;
assign n3721 =  ( n3472 ) ? ( VREG_7_12 ) : ( n3720 ) ;
assign n3722 =  ( n3471 ) ? ( VREG_7_13 ) : ( n3721 ) ;
assign n3723 =  ( n3470 ) ? ( VREG_7_14 ) : ( n3722 ) ;
assign n3724 =  ( n3469 ) ? ( VREG_7_15 ) : ( n3723 ) ;
assign n3725 =  ( n3468 ) ? ( VREG_8_0 ) : ( n3724 ) ;
assign n3726 =  ( n3467 ) ? ( VREG_8_1 ) : ( n3725 ) ;
assign n3727 =  ( n3466 ) ? ( VREG_8_2 ) : ( n3726 ) ;
assign n3728 =  ( n3465 ) ? ( VREG_8_3 ) : ( n3727 ) ;
assign n3729 =  ( n3464 ) ? ( VREG_8_4 ) : ( n3728 ) ;
assign n3730 =  ( n3463 ) ? ( VREG_8_5 ) : ( n3729 ) ;
assign n3731 =  ( n3462 ) ? ( VREG_8_6 ) : ( n3730 ) ;
assign n3732 =  ( n3461 ) ? ( VREG_8_7 ) : ( n3731 ) ;
assign n3733 =  ( n3460 ) ? ( VREG_8_8 ) : ( n3732 ) ;
assign n3734 =  ( n3459 ) ? ( VREG_8_9 ) : ( n3733 ) ;
assign n3735 =  ( n3458 ) ? ( VREG_8_10 ) : ( n3734 ) ;
assign n3736 =  ( n3457 ) ? ( VREG_8_11 ) : ( n3735 ) ;
assign n3737 =  ( n3456 ) ? ( VREG_8_12 ) : ( n3736 ) ;
assign n3738 =  ( n3455 ) ? ( VREG_8_13 ) : ( n3737 ) ;
assign n3739 =  ( n3454 ) ? ( VREG_8_14 ) : ( n3738 ) ;
assign n3740 =  ( n3453 ) ? ( VREG_8_15 ) : ( n3739 ) ;
assign n3741 =  ( n3452 ) ? ( VREG_9_0 ) : ( n3740 ) ;
assign n3742 =  ( n3451 ) ? ( VREG_9_1 ) : ( n3741 ) ;
assign n3743 =  ( n3450 ) ? ( VREG_9_2 ) : ( n3742 ) ;
assign n3744 =  ( n3449 ) ? ( VREG_9_3 ) : ( n3743 ) ;
assign n3745 =  ( n3448 ) ? ( VREG_9_4 ) : ( n3744 ) ;
assign n3746 =  ( n3447 ) ? ( VREG_9_5 ) : ( n3745 ) ;
assign n3747 =  ( n3446 ) ? ( VREG_9_6 ) : ( n3746 ) ;
assign n3748 =  ( n3445 ) ? ( VREG_9_7 ) : ( n3747 ) ;
assign n3749 =  ( n3444 ) ? ( VREG_9_8 ) : ( n3748 ) ;
assign n3750 =  ( n3443 ) ? ( VREG_9_9 ) : ( n3749 ) ;
assign n3751 =  ( n3442 ) ? ( VREG_9_10 ) : ( n3750 ) ;
assign n3752 =  ( n3441 ) ? ( VREG_9_11 ) : ( n3751 ) ;
assign n3753 =  ( n3440 ) ? ( VREG_9_12 ) : ( n3752 ) ;
assign n3754 =  ( n3439 ) ? ( VREG_9_13 ) : ( n3753 ) ;
assign n3755 =  ( n3438 ) ? ( VREG_9_14 ) : ( n3754 ) ;
assign n3756 =  ( n3437 ) ? ( VREG_9_15 ) : ( n3755 ) ;
assign n3757 =  ( n3436 ) ? ( VREG_10_0 ) : ( n3756 ) ;
assign n3758 =  ( n3435 ) ? ( VREG_10_1 ) : ( n3757 ) ;
assign n3759 =  ( n3434 ) ? ( VREG_10_2 ) : ( n3758 ) ;
assign n3760 =  ( n3433 ) ? ( VREG_10_3 ) : ( n3759 ) ;
assign n3761 =  ( n3432 ) ? ( VREG_10_4 ) : ( n3760 ) ;
assign n3762 =  ( n3431 ) ? ( VREG_10_5 ) : ( n3761 ) ;
assign n3763 =  ( n3430 ) ? ( VREG_10_6 ) : ( n3762 ) ;
assign n3764 =  ( n3429 ) ? ( VREG_10_7 ) : ( n3763 ) ;
assign n3765 =  ( n3428 ) ? ( VREG_10_8 ) : ( n3764 ) ;
assign n3766 =  ( n3427 ) ? ( VREG_10_9 ) : ( n3765 ) ;
assign n3767 =  ( n3426 ) ? ( VREG_10_10 ) : ( n3766 ) ;
assign n3768 =  ( n3425 ) ? ( VREG_10_11 ) : ( n3767 ) ;
assign n3769 =  ( n3424 ) ? ( VREG_10_12 ) : ( n3768 ) ;
assign n3770 =  ( n3423 ) ? ( VREG_10_13 ) : ( n3769 ) ;
assign n3771 =  ( n3422 ) ? ( VREG_10_14 ) : ( n3770 ) ;
assign n3772 =  ( n3421 ) ? ( VREG_10_15 ) : ( n3771 ) ;
assign n3773 =  ( n3420 ) ? ( VREG_11_0 ) : ( n3772 ) ;
assign n3774 =  ( n3419 ) ? ( VREG_11_1 ) : ( n3773 ) ;
assign n3775 =  ( n3418 ) ? ( VREG_11_2 ) : ( n3774 ) ;
assign n3776 =  ( n3417 ) ? ( VREG_11_3 ) : ( n3775 ) ;
assign n3777 =  ( n3416 ) ? ( VREG_11_4 ) : ( n3776 ) ;
assign n3778 =  ( n3415 ) ? ( VREG_11_5 ) : ( n3777 ) ;
assign n3779 =  ( n3414 ) ? ( VREG_11_6 ) : ( n3778 ) ;
assign n3780 =  ( n3413 ) ? ( VREG_11_7 ) : ( n3779 ) ;
assign n3781 =  ( n3412 ) ? ( VREG_11_8 ) : ( n3780 ) ;
assign n3782 =  ( n3411 ) ? ( VREG_11_9 ) : ( n3781 ) ;
assign n3783 =  ( n3410 ) ? ( VREG_11_10 ) : ( n3782 ) ;
assign n3784 =  ( n3409 ) ? ( VREG_11_11 ) : ( n3783 ) ;
assign n3785 =  ( n3408 ) ? ( VREG_11_12 ) : ( n3784 ) ;
assign n3786 =  ( n3407 ) ? ( VREG_11_13 ) : ( n3785 ) ;
assign n3787 =  ( n3406 ) ? ( VREG_11_14 ) : ( n3786 ) ;
assign n3788 =  ( n3405 ) ? ( VREG_11_15 ) : ( n3787 ) ;
assign n3789 =  ( n3404 ) ? ( VREG_12_0 ) : ( n3788 ) ;
assign n3790 =  ( n3403 ) ? ( VREG_12_1 ) : ( n3789 ) ;
assign n3791 =  ( n3402 ) ? ( VREG_12_2 ) : ( n3790 ) ;
assign n3792 =  ( n3401 ) ? ( VREG_12_3 ) : ( n3791 ) ;
assign n3793 =  ( n3400 ) ? ( VREG_12_4 ) : ( n3792 ) ;
assign n3794 =  ( n3399 ) ? ( VREG_12_5 ) : ( n3793 ) ;
assign n3795 =  ( n3398 ) ? ( VREG_12_6 ) : ( n3794 ) ;
assign n3796 =  ( n3397 ) ? ( VREG_12_7 ) : ( n3795 ) ;
assign n3797 =  ( n3396 ) ? ( VREG_12_8 ) : ( n3796 ) ;
assign n3798 =  ( n3395 ) ? ( VREG_12_9 ) : ( n3797 ) ;
assign n3799 =  ( n3394 ) ? ( VREG_12_10 ) : ( n3798 ) ;
assign n3800 =  ( n3393 ) ? ( VREG_12_11 ) : ( n3799 ) ;
assign n3801 =  ( n3392 ) ? ( VREG_12_12 ) : ( n3800 ) ;
assign n3802 =  ( n3391 ) ? ( VREG_12_13 ) : ( n3801 ) ;
assign n3803 =  ( n3390 ) ? ( VREG_12_14 ) : ( n3802 ) ;
assign n3804 =  ( n3389 ) ? ( VREG_12_15 ) : ( n3803 ) ;
assign n3805 =  ( n3388 ) ? ( VREG_13_0 ) : ( n3804 ) ;
assign n3806 =  ( n3387 ) ? ( VREG_13_1 ) : ( n3805 ) ;
assign n3807 =  ( n3386 ) ? ( VREG_13_2 ) : ( n3806 ) ;
assign n3808 =  ( n3385 ) ? ( VREG_13_3 ) : ( n3807 ) ;
assign n3809 =  ( n3384 ) ? ( VREG_13_4 ) : ( n3808 ) ;
assign n3810 =  ( n3383 ) ? ( VREG_13_5 ) : ( n3809 ) ;
assign n3811 =  ( n3382 ) ? ( VREG_13_6 ) : ( n3810 ) ;
assign n3812 =  ( n3381 ) ? ( VREG_13_7 ) : ( n3811 ) ;
assign n3813 =  ( n3380 ) ? ( VREG_13_8 ) : ( n3812 ) ;
assign n3814 =  ( n3379 ) ? ( VREG_13_9 ) : ( n3813 ) ;
assign n3815 =  ( n3378 ) ? ( VREG_13_10 ) : ( n3814 ) ;
assign n3816 =  ( n3377 ) ? ( VREG_13_11 ) : ( n3815 ) ;
assign n3817 =  ( n3376 ) ? ( VREG_13_12 ) : ( n3816 ) ;
assign n3818 =  ( n3375 ) ? ( VREG_13_13 ) : ( n3817 ) ;
assign n3819 =  ( n3374 ) ? ( VREG_13_14 ) : ( n3818 ) ;
assign n3820 =  ( n3373 ) ? ( VREG_13_15 ) : ( n3819 ) ;
assign n3821 =  ( n3372 ) ? ( VREG_14_0 ) : ( n3820 ) ;
assign n3822 =  ( n3371 ) ? ( VREG_14_1 ) : ( n3821 ) ;
assign n3823 =  ( n3370 ) ? ( VREG_14_2 ) : ( n3822 ) ;
assign n3824 =  ( n3369 ) ? ( VREG_14_3 ) : ( n3823 ) ;
assign n3825 =  ( n3368 ) ? ( VREG_14_4 ) : ( n3824 ) ;
assign n3826 =  ( n3367 ) ? ( VREG_14_5 ) : ( n3825 ) ;
assign n3827 =  ( n3366 ) ? ( VREG_14_6 ) : ( n3826 ) ;
assign n3828 =  ( n3365 ) ? ( VREG_14_7 ) : ( n3827 ) ;
assign n3829 =  ( n3364 ) ? ( VREG_14_8 ) : ( n3828 ) ;
assign n3830 =  ( n3363 ) ? ( VREG_14_9 ) : ( n3829 ) ;
assign n3831 =  ( n3362 ) ? ( VREG_14_10 ) : ( n3830 ) ;
assign n3832 =  ( n3361 ) ? ( VREG_14_11 ) : ( n3831 ) ;
assign n3833 =  ( n3360 ) ? ( VREG_14_12 ) : ( n3832 ) ;
assign n3834 =  ( n3359 ) ? ( VREG_14_13 ) : ( n3833 ) ;
assign n3835 =  ( n3358 ) ? ( VREG_14_14 ) : ( n3834 ) ;
assign n3836 =  ( n3357 ) ? ( VREG_14_15 ) : ( n3835 ) ;
assign n3837 =  ( n3356 ) ? ( VREG_15_0 ) : ( n3836 ) ;
assign n3838 =  ( n3355 ) ? ( VREG_15_1 ) : ( n3837 ) ;
assign n3839 =  ( n3354 ) ? ( VREG_15_2 ) : ( n3838 ) ;
assign n3840 =  ( n3353 ) ? ( VREG_15_3 ) : ( n3839 ) ;
assign n3841 =  ( n3352 ) ? ( VREG_15_4 ) : ( n3840 ) ;
assign n3842 =  ( n3351 ) ? ( VREG_15_5 ) : ( n3841 ) ;
assign n3843 =  ( n3350 ) ? ( VREG_15_6 ) : ( n3842 ) ;
assign n3844 =  ( n3349 ) ? ( VREG_15_7 ) : ( n3843 ) ;
assign n3845 =  ( n3348 ) ? ( VREG_15_8 ) : ( n3844 ) ;
assign n3846 =  ( n3347 ) ? ( VREG_15_9 ) : ( n3845 ) ;
assign n3847 =  ( n3346 ) ? ( VREG_15_10 ) : ( n3846 ) ;
assign n3848 =  ( n3345 ) ? ( VREG_15_11 ) : ( n3847 ) ;
assign n3849 =  ( n3344 ) ? ( VREG_15_12 ) : ( n3848 ) ;
assign n3850 =  ( n3343 ) ? ( VREG_15_13 ) : ( n3849 ) ;
assign n3851 =  ( n3342 ) ? ( VREG_15_14 ) : ( n3850 ) ;
assign n3852 =  ( n3341 ) ? ( VREG_15_15 ) : ( n3851 ) ;
assign n3853 =  ( n3340 ) ? ( VREG_16_0 ) : ( n3852 ) ;
assign n3854 =  ( n3339 ) ? ( VREG_16_1 ) : ( n3853 ) ;
assign n3855 =  ( n3338 ) ? ( VREG_16_2 ) : ( n3854 ) ;
assign n3856 =  ( n3337 ) ? ( VREG_16_3 ) : ( n3855 ) ;
assign n3857 =  ( n3336 ) ? ( VREG_16_4 ) : ( n3856 ) ;
assign n3858 =  ( n3335 ) ? ( VREG_16_5 ) : ( n3857 ) ;
assign n3859 =  ( n3334 ) ? ( VREG_16_6 ) : ( n3858 ) ;
assign n3860 =  ( n3333 ) ? ( VREG_16_7 ) : ( n3859 ) ;
assign n3861 =  ( n3332 ) ? ( VREG_16_8 ) : ( n3860 ) ;
assign n3862 =  ( n3331 ) ? ( VREG_16_9 ) : ( n3861 ) ;
assign n3863 =  ( n3330 ) ? ( VREG_16_10 ) : ( n3862 ) ;
assign n3864 =  ( n3329 ) ? ( VREG_16_11 ) : ( n3863 ) ;
assign n3865 =  ( n3328 ) ? ( VREG_16_12 ) : ( n3864 ) ;
assign n3866 =  ( n3327 ) ? ( VREG_16_13 ) : ( n3865 ) ;
assign n3867 =  ( n3326 ) ? ( VREG_16_14 ) : ( n3866 ) ;
assign n3868 =  ( n3325 ) ? ( VREG_16_15 ) : ( n3867 ) ;
assign n3869 =  ( n3324 ) ? ( VREG_17_0 ) : ( n3868 ) ;
assign n3870 =  ( n3323 ) ? ( VREG_17_1 ) : ( n3869 ) ;
assign n3871 =  ( n3322 ) ? ( VREG_17_2 ) : ( n3870 ) ;
assign n3872 =  ( n3321 ) ? ( VREG_17_3 ) : ( n3871 ) ;
assign n3873 =  ( n3320 ) ? ( VREG_17_4 ) : ( n3872 ) ;
assign n3874 =  ( n3319 ) ? ( VREG_17_5 ) : ( n3873 ) ;
assign n3875 =  ( n3318 ) ? ( VREG_17_6 ) : ( n3874 ) ;
assign n3876 =  ( n3317 ) ? ( VREG_17_7 ) : ( n3875 ) ;
assign n3877 =  ( n3316 ) ? ( VREG_17_8 ) : ( n3876 ) ;
assign n3878 =  ( n3315 ) ? ( VREG_17_9 ) : ( n3877 ) ;
assign n3879 =  ( n3314 ) ? ( VREG_17_10 ) : ( n3878 ) ;
assign n3880 =  ( n3313 ) ? ( VREG_17_11 ) : ( n3879 ) ;
assign n3881 =  ( n3312 ) ? ( VREG_17_12 ) : ( n3880 ) ;
assign n3882 =  ( n3311 ) ? ( VREG_17_13 ) : ( n3881 ) ;
assign n3883 =  ( n3310 ) ? ( VREG_17_14 ) : ( n3882 ) ;
assign n3884 =  ( n3309 ) ? ( VREG_17_15 ) : ( n3883 ) ;
assign n3885 =  ( n3308 ) ? ( VREG_18_0 ) : ( n3884 ) ;
assign n3886 =  ( n3307 ) ? ( VREG_18_1 ) : ( n3885 ) ;
assign n3887 =  ( n3306 ) ? ( VREG_18_2 ) : ( n3886 ) ;
assign n3888 =  ( n3305 ) ? ( VREG_18_3 ) : ( n3887 ) ;
assign n3889 =  ( n3304 ) ? ( VREG_18_4 ) : ( n3888 ) ;
assign n3890 =  ( n3303 ) ? ( VREG_18_5 ) : ( n3889 ) ;
assign n3891 =  ( n3302 ) ? ( VREG_18_6 ) : ( n3890 ) ;
assign n3892 =  ( n3301 ) ? ( VREG_18_7 ) : ( n3891 ) ;
assign n3893 =  ( n3300 ) ? ( VREG_18_8 ) : ( n3892 ) ;
assign n3894 =  ( n3299 ) ? ( VREG_18_9 ) : ( n3893 ) ;
assign n3895 =  ( n3298 ) ? ( VREG_18_10 ) : ( n3894 ) ;
assign n3896 =  ( n3297 ) ? ( VREG_18_11 ) : ( n3895 ) ;
assign n3897 =  ( n3296 ) ? ( VREG_18_12 ) : ( n3896 ) ;
assign n3898 =  ( n3295 ) ? ( VREG_18_13 ) : ( n3897 ) ;
assign n3899 =  ( n3294 ) ? ( VREG_18_14 ) : ( n3898 ) ;
assign n3900 =  ( n3293 ) ? ( VREG_18_15 ) : ( n3899 ) ;
assign n3901 =  ( n3292 ) ? ( VREG_19_0 ) : ( n3900 ) ;
assign n3902 =  ( n3291 ) ? ( VREG_19_1 ) : ( n3901 ) ;
assign n3903 =  ( n3290 ) ? ( VREG_19_2 ) : ( n3902 ) ;
assign n3904 =  ( n3289 ) ? ( VREG_19_3 ) : ( n3903 ) ;
assign n3905 =  ( n3288 ) ? ( VREG_19_4 ) : ( n3904 ) ;
assign n3906 =  ( n3287 ) ? ( VREG_19_5 ) : ( n3905 ) ;
assign n3907 =  ( n3286 ) ? ( VREG_19_6 ) : ( n3906 ) ;
assign n3908 =  ( n3285 ) ? ( VREG_19_7 ) : ( n3907 ) ;
assign n3909 =  ( n3284 ) ? ( VREG_19_8 ) : ( n3908 ) ;
assign n3910 =  ( n3283 ) ? ( VREG_19_9 ) : ( n3909 ) ;
assign n3911 =  ( n3282 ) ? ( VREG_19_10 ) : ( n3910 ) ;
assign n3912 =  ( n3281 ) ? ( VREG_19_11 ) : ( n3911 ) ;
assign n3913 =  ( n3280 ) ? ( VREG_19_12 ) : ( n3912 ) ;
assign n3914 =  ( n3279 ) ? ( VREG_19_13 ) : ( n3913 ) ;
assign n3915 =  ( n3278 ) ? ( VREG_19_14 ) : ( n3914 ) ;
assign n3916 =  ( n3277 ) ? ( VREG_19_15 ) : ( n3915 ) ;
assign n3917 =  ( n3276 ) ? ( VREG_20_0 ) : ( n3916 ) ;
assign n3918 =  ( n3275 ) ? ( VREG_20_1 ) : ( n3917 ) ;
assign n3919 =  ( n3274 ) ? ( VREG_20_2 ) : ( n3918 ) ;
assign n3920 =  ( n3273 ) ? ( VREG_20_3 ) : ( n3919 ) ;
assign n3921 =  ( n3272 ) ? ( VREG_20_4 ) : ( n3920 ) ;
assign n3922 =  ( n3271 ) ? ( VREG_20_5 ) : ( n3921 ) ;
assign n3923 =  ( n3270 ) ? ( VREG_20_6 ) : ( n3922 ) ;
assign n3924 =  ( n3269 ) ? ( VREG_20_7 ) : ( n3923 ) ;
assign n3925 =  ( n3268 ) ? ( VREG_20_8 ) : ( n3924 ) ;
assign n3926 =  ( n3267 ) ? ( VREG_20_9 ) : ( n3925 ) ;
assign n3927 =  ( n3266 ) ? ( VREG_20_10 ) : ( n3926 ) ;
assign n3928 =  ( n3265 ) ? ( VREG_20_11 ) : ( n3927 ) ;
assign n3929 =  ( n3264 ) ? ( VREG_20_12 ) : ( n3928 ) ;
assign n3930 =  ( n3263 ) ? ( VREG_20_13 ) : ( n3929 ) ;
assign n3931 =  ( n3262 ) ? ( VREG_20_14 ) : ( n3930 ) ;
assign n3932 =  ( n3261 ) ? ( VREG_20_15 ) : ( n3931 ) ;
assign n3933 =  ( n3260 ) ? ( VREG_21_0 ) : ( n3932 ) ;
assign n3934 =  ( n3259 ) ? ( VREG_21_1 ) : ( n3933 ) ;
assign n3935 =  ( n3258 ) ? ( VREG_21_2 ) : ( n3934 ) ;
assign n3936 =  ( n3257 ) ? ( VREG_21_3 ) : ( n3935 ) ;
assign n3937 =  ( n3256 ) ? ( VREG_21_4 ) : ( n3936 ) ;
assign n3938 =  ( n3255 ) ? ( VREG_21_5 ) : ( n3937 ) ;
assign n3939 =  ( n3254 ) ? ( VREG_21_6 ) : ( n3938 ) ;
assign n3940 =  ( n3253 ) ? ( VREG_21_7 ) : ( n3939 ) ;
assign n3941 =  ( n3252 ) ? ( VREG_21_8 ) : ( n3940 ) ;
assign n3942 =  ( n3251 ) ? ( VREG_21_9 ) : ( n3941 ) ;
assign n3943 =  ( n3250 ) ? ( VREG_21_10 ) : ( n3942 ) ;
assign n3944 =  ( n3249 ) ? ( VREG_21_11 ) : ( n3943 ) ;
assign n3945 =  ( n3248 ) ? ( VREG_21_12 ) : ( n3944 ) ;
assign n3946 =  ( n3247 ) ? ( VREG_21_13 ) : ( n3945 ) ;
assign n3947 =  ( n3246 ) ? ( VREG_21_14 ) : ( n3946 ) ;
assign n3948 =  ( n3245 ) ? ( VREG_21_15 ) : ( n3947 ) ;
assign n3949 =  ( n3244 ) ? ( VREG_22_0 ) : ( n3948 ) ;
assign n3950 =  ( n3243 ) ? ( VREG_22_1 ) : ( n3949 ) ;
assign n3951 =  ( n3242 ) ? ( VREG_22_2 ) : ( n3950 ) ;
assign n3952 =  ( n3241 ) ? ( VREG_22_3 ) : ( n3951 ) ;
assign n3953 =  ( n3240 ) ? ( VREG_22_4 ) : ( n3952 ) ;
assign n3954 =  ( n3239 ) ? ( VREG_22_5 ) : ( n3953 ) ;
assign n3955 =  ( n3238 ) ? ( VREG_22_6 ) : ( n3954 ) ;
assign n3956 =  ( n3237 ) ? ( VREG_22_7 ) : ( n3955 ) ;
assign n3957 =  ( n3236 ) ? ( VREG_22_8 ) : ( n3956 ) ;
assign n3958 =  ( n3235 ) ? ( VREG_22_9 ) : ( n3957 ) ;
assign n3959 =  ( n3234 ) ? ( VREG_22_10 ) : ( n3958 ) ;
assign n3960 =  ( n3233 ) ? ( VREG_22_11 ) : ( n3959 ) ;
assign n3961 =  ( n3232 ) ? ( VREG_22_12 ) : ( n3960 ) ;
assign n3962 =  ( n3231 ) ? ( VREG_22_13 ) : ( n3961 ) ;
assign n3963 =  ( n3230 ) ? ( VREG_22_14 ) : ( n3962 ) ;
assign n3964 =  ( n3229 ) ? ( VREG_22_15 ) : ( n3963 ) ;
assign n3965 =  ( n3228 ) ? ( VREG_23_0 ) : ( n3964 ) ;
assign n3966 =  ( n3227 ) ? ( VREG_23_1 ) : ( n3965 ) ;
assign n3967 =  ( n3226 ) ? ( VREG_23_2 ) : ( n3966 ) ;
assign n3968 =  ( n3225 ) ? ( VREG_23_3 ) : ( n3967 ) ;
assign n3969 =  ( n3224 ) ? ( VREG_23_4 ) : ( n3968 ) ;
assign n3970 =  ( n3223 ) ? ( VREG_23_5 ) : ( n3969 ) ;
assign n3971 =  ( n3222 ) ? ( VREG_23_6 ) : ( n3970 ) ;
assign n3972 =  ( n3221 ) ? ( VREG_23_7 ) : ( n3971 ) ;
assign n3973 =  ( n3220 ) ? ( VREG_23_8 ) : ( n3972 ) ;
assign n3974 =  ( n3219 ) ? ( VREG_23_9 ) : ( n3973 ) ;
assign n3975 =  ( n3218 ) ? ( VREG_23_10 ) : ( n3974 ) ;
assign n3976 =  ( n3217 ) ? ( VREG_23_11 ) : ( n3975 ) ;
assign n3977 =  ( n3216 ) ? ( VREG_23_12 ) : ( n3976 ) ;
assign n3978 =  ( n3215 ) ? ( VREG_23_13 ) : ( n3977 ) ;
assign n3979 =  ( n3214 ) ? ( VREG_23_14 ) : ( n3978 ) ;
assign n3980 =  ( n3213 ) ? ( VREG_23_15 ) : ( n3979 ) ;
assign n3981 =  ( n3212 ) ? ( VREG_24_0 ) : ( n3980 ) ;
assign n3982 =  ( n3211 ) ? ( VREG_24_1 ) : ( n3981 ) ;
assign n3983 =  ( n3210 ) ? ( VREG_24_2 ) : ( n3982 ) ;
assign n3984 =  ( n3209 ) ? ( VREG_24_3 ) : ( n3983 ) ;
assign n3985 =  ( n3208 ) ? ( VREG_24_4 ) : ( n3984 ) ;
assign n3986 =  ( n3207 ) ? ( VREG_24_5 ) : ( n3985 ) ;
assign n3987 =  ( n3206 ) ? ( VREG_24_6 ) : ( n3986 ) ;
assign n3988 =  ( n3205 ) ? ( VREG_24_7 ) : ( n3987 ) ;
assign n3989 =  ( n3204 ) ? ( VREG_24_8 ) : ( n3988 ) ;
assign n3990 =  ( n3203 ) ? ( VREG_24_9 ) : ( n3989 ) ;
assign n3991 =  ( n3202 ) ? ( VREG_24_10 ) : ( n3990 ) ;
assign n3992 =  ( n3201 ) ? ( VREG_24_11 ) : ( n3991 ) ;
assign n3993 =  ( n3200 ) ? ( VREG_24_12 ) : ( n3992 ) ;
assign n3994 =  ( n3199 ) ? ( VREG_24_13 ) : ( n3993 ) ;
assign n3995 =  ( n3198 ) ? ( VREG_24_14 ) : ( n3994 ) ;
assign n3996 =  ( n3197 ) ? ( VREG_24_15 ) : ( n3995 ) ;
assign n3997 =  ( n3196 ) ? ( VREG_25_0 ) : ( n3996 ) ;
assign n3998 =  ( n3195 ) ? ( VREG_25_1 ) : ( n3997 ) ;
assign n3999 =  ( n3194 ) ? ( VREG_25_2 ) : ( n3998 ) ;
assign n4000 =  ( n3193 ) ? ( VREG_25_3 ) : ( n3999 ) ;
assign n4001 =  ( n3192 ) ? ( VREG_25_4 ) : ( n4000 ) ;
assign n4002 =  ( n3191 ) ? ( VREG_25_5 ) : ( n4001 ) ;
assign n4003 =  ( n3190 ) ? ( VREG_25_6 ) : ( n4002 ) ;
assign n4004 =  ( n3189 ) ? ( VREG_25_7 ) : ( n4003 ) ;
assign n4005 =  ( n3188 ) ? ( VREG_25_8 ) : ( n4004 ) ;
assign n4006 =  ( n3187 ) ? ( VREG_25_9 ) : ( n4005 ) ;
assign n4007 =  ( n3186 ) ? ( VREG_25_10 ) : ( n4006 ) ;
assign n4008 =  ( n3185 ) ? ( VREG_25_11 ) : ( n4007 ) ;
assign n4009 =  ( n3184 ) ? ( VREG_25_12 ) : ( n4008 ) ;
assign n4010 =  ( n3183 ) ? ( VREG_25_13 ) : ( n4009 ) ;
assign n4011 =  ( n3182 ) ? ( VREG_25_14 ) : ( n4010 ) ;
assign n4012 =  ( n3181 ) ? ( VREG_25_15 ) : ( n4011 ) ;
assign n4013 =  ( n3180 ) ? ( VREG_26_0 ) : ( n4012 ) ;
assign n4014 =  ( n3179 ) ? ( VREG_26_1 ) : ( n4013 ) ;
assign n4015 =  ( n3178 ) ? ( VREG_26_2 ) : ( n4014 ) ;
assign n4016 =  ( n3177 ) ? ( VREG_26_3 ) : ( n4015 ) ;
assign n4017 =  ( n3176 ) ? ( VREG_26_4 ) : ( n4016 ) ;
assign n4018 =  ( n3175 ) ? ( VREG_26_5 ) : ( n4017 ) ;
assign n4019 =  ( n3174 ) ? ( VREG_26_6 ) : ( n4018 ) ;
assign n4020 =  ( n3173 ) ? ( VREG_26_7 ) : ( n4019 ) ;
assign n4021 =  ( n3172 ) ? ( VREG_26_8 ) : ( n4020 ) ;
assign n4022 =  ( n3171 ) ? ( VREG_26_9 ) : ( n4021 ) ;
assign n4023 =  ( n3170 ) ? ( VREG_26_10 ) : ( n4022 ) ;
assign n4024 =  ( n3169 ) ? ( VREG_26_11 ) : ( n4023 ) ;
assign n4025 =  ( n3168 ) ? ( VREG_26_12 ) : ( n4024 ) ;
assign n4026 =  ( n3167 ) ? ( VREG_26_13 ) : ( n4025 ) ;
assign n4027 =  ( n3166 ) ? ( VREG_26_14 ) : ( n4026 ) ;
assign n4028 =  ( n3165 ) ? ( VREG_26_15 ) : ( n4027 ) ;
assign n4029 =  ( n3164 ) ? ( VREG_27_0 ) : ( n4028 ) ;
assign n4030 =  ( n3163 ) ? ( VREG_27_1 ) : ( n4029 ) ;
assign n4031 =  ( n3162 ) ? ( VREG_27_2 ) : ( n4030 ) ;
assign n4032 =  ( n3161 ) ? ( VREG_27_3 ) : ( n4031 ) ;
assign n4033 =  ( n3160 ) ? ( VREG_27_4 ) : ( n4032 ) ;
assign n4034 =  ( n3159 ) ? ( VREG_27_5 ) : ( n4033 ) ;
assign n4035 =  ( n3158 ) ? ( VREG_27_6 ) : ( n4034 ) ;
assign n4036 =  ( n3157 ) ? ( VREG_27_7 ) : ( n4035 ) ;
assign n4037 =  ( n3156 ) ? ( VREG_27_8 ) : ( n4036 ) ;
assign n4038 =  ( n3155 ) ? ( VREG_27_9 ) : ( n4037 ) ;
assign n4039 =  ( n3154 ) ? ( VREG_27_10 ) : ( n4038 ) ;
assign n4040 =  ( n3153 ) ? ( VREG_27_11 ) : ( n4039 ) ;
assign n4041 =  ( n3152 ) ? ( VREG_27_12 ) : ( n4040 ) ;
assign n4042 =  ( n3151 ) ? ( VREG_27_13 ) : ( n4041 ) ;
assign n4043 =  ( n3150 ) ? ( VREG_27_14 ) : ( n4042 ) ;
assign n4044 =  ( n3149 ) ? ( VREG_27_15 ) : ( n4043 ) ;
assign n4045 =  ( n3148 ) ? ( VREG_28_0 ) : ( n4044 ) ;
assign n4046 =  ( n3147 ) ? ( VREG_28_1 ) : ( n4045 ) ;
assign n4047 =  ( n3146 ) ? ( VREG_28_2 ) : ( n4046 ) ;
assign n4048 =  ( n3145 ) ? ( VREG_28_3 ) : ( n4047 ) ;
assign n4049 =  ( n3144 ) ? ( VREG_28_4 ) : ( n4048 ) ;
assign n4050 =  ( n3143 ) ? ( VREG_28_5 ) : ( n4049 ) ;
assign n4051 =  ( n3142 ) ? ( VREG_28_6 ) : ( n4050 ) ;
assign n4052 =  ( n3141 ) ? ( VREG_28_7 ) : ( n4051 ) ;
assign n4053 =  ( n3140 ) ? ( VREG_28_8 ) : ( n4052 ) ;
assign n4054 =  ( n3139 ) ? ( VREG_28_9 ) : ( n4053 ) ;
assign n4055 =  ( n3138 ) ? ( VREG_28_10 ) : ( n4054 ) ;
assign n4056 =  ( n3137 ) ? ( VREG_28_11 ) : ( n4055 ) ;
assign n4057 =  ( n3136 ) ? ( VREG_28_12 ) : ( n4056 ) ;
assign n4058 =  ( n3135 ) ? ( VREG_28_13 ) : ( n4057 ) ;
assign n4059 =  ( n3134 ) ? ( VREG_28_14 ) : ( n4058 ) ;
assign n4060 =  ( n3133 ) ? ( VREG_28_15 ) : ( n4059 ) ;
assign n4061 =  ( n3132 ) ? ( VREG_29_0 ) : ( n4060 ) ;
assign n4062 =  ( n3131 ) ? ( VREG_29_1 ) : ( n4061 ) ;
assign n4063 =  ( n3130 ) ? ( VREG_29_2 ) : ( n4062 ) ;
assign n4064 =  ( n3129 ) ? ( VREG_29_3 ) : ( n4063 ) ;
assign n4065 =  ( n3128 ) ? ( VREG_29_4 ) : ( n4064 ) ;
assign n4066 =  ( n3127 ) ? ( VREG_29_5 ) : ( n4065 ) ;
assign n4067 =  ( n3126 ) ? ( VREG_29_6 ) : ( n4066 ) ;
assign n4068 =  ( n3125 ) ? ( VREG_29_7 ) : ( n4067 ) ;
assign n4069 =  ( n3124 ) ? ( VREG_29_8 ) : ( n4068 ) ;
assign n4070 =  ( n3123 ) ? ( VREG_29_9 ) : ( n4069 ) ;
assign n4071 =  ( n3122 ) ? ( VREG_29_10 ) : ( n4070 ) ;
assign n4072 =  ( n3121 ) ? ( VREG_29_11 ) : ( n4071 ) ;
assign n4073 =  ( n3120 ) ? ( VREG_29_12 ) : ( n4072 ) ;
assign n4074 =  ( n3119 ) ? ( VREG_29_13 ) : ( n4073 ) ;
assign n4075 =  ( n3118 ) ? ( VREG_29_14 ) : ( n4074 ) ;
assign n4076 =  ( n3117 ) ? ( VREG_29_15 ) : ( n4075 ) ;
assign n4077 =  ( n3116 ) ? ( VREG_30_0 ) : ( n4076 ) ;
assign n4078 =  ( n3115 ) ? ( VREG_30_1 ) : ( n4077 ) ;
assign n4079 =  ( n3114 ) ? ( VREG_30_2 ) : ( n4078 ) ;
assign n4080 =  ( n3113 ) ? ( VREG_30_3 ) : ( n4079 ) ;
assign n4081 =  ( n3112 ) ? ( VREG_30_4 ) : ( n4080 ) ;
assign n4082 =  ( n3111 ) ? ( VREG_30_5 ) : ( n4081 ) ;
assign n4083 =  ( n3110 ) ? ( VREG_30_6 ) : ( n4082 ) ;
assign n4084 =  ( n3109 ) ? ( VREG_30_7 ) : ( n4083 ) ;
assign n4085 =  ( n3108 ) ? ( VREG_30_8 ) : ( n4084 ) ;
assign n4086 =  ( n3107 ) ? ( VREG_30_9 ) : ( n4085 ) ;
assign n4087 =  ( n3106 ) ? ( VREG_30_10 ) : ( n4086 ) ;
assign n4088 =  ( n3105 ) ? ( VREG_30_11 ) : ( n4087 ) ;
assign n4089 =  ( n3104 ) ? ( VREG_30_12 ) : ( n4088 ) ;
assign n4090 =  ( n3103 ) ? ( VREG_30_13 ) : ( n4089 ) ;
assign n4091 =  ( n3102 ) ? ( VREG_30_14 ) : ( n4090 ) ;
assign n4092 =  ( n3101 ) ? ( VREG_30_15 ) : ( n4091 ) ;
assign n4093 =  ( n3100 ) ? ( VREG_31_0 ) : ( n4092 ) ;
assign n4094 =  ( n3098 ) ? ( VREG_31_1 ) : ( n4093 ) ;
assign n4095 =  ( n3096 ) ? ( VREG_31_2 ) : ( n4094 ) ;
assign n4096 =  ( n3094 ) ? ( VREG_31_3 ) : ( n4095 ) ;
assign n4097 =  ( n3092 ) ? ( VREG_31_4 ) : ( n4096 ) ;
assign n4098 =  ( n3090 ) ? ( VREG_31_5 ) : ( n4097 ) ;
assign n4099 =  ( n3088 ) ? ( VREG_31_6 ) : ( n4098 ) ;
assign n4100 =  ( n3086 ) ? ( VREG_31_7 ) : ( n4099 ) ;
assign n4101 =  ( n3084 ) ? ( VREG_31_8 ) : ( n4100 ) ;
assign n4102 =  ( n3082 ) ? ( VREG_31_9 ) : ( n4101 ) ;
assign n4103 =  ( n3080 ) ? ( VREG_31_10 ) : ( n4102 ) ;
assign n4104 =  ( n3078 ) ? ( VREG_31_11 ) : ( n4103 ) ;
assign n4105 =  ( n3076 ) ? ( VREG_31_12 ) : ( n4104 ) ;
assign n4106 =  ( n3074 ) ? ( VREG_31_13 ) : ( n4105 ) ;
assign n4107 =  ( n3072 ) ? ( VREG_31_14 ) : ( n4106 ) ;
assign n4108 =  ( n3070 ) ? ( VREG_31_15 ) : ( n4107 ) ;
assign n4109 =  ( n4108 ) + ( n140 )  ;
assign n4110 =  ( n4108 ) - ( n140 )  ;
assign n4111 =  ( n4108 ) & ( n140 )  ;
assign n4112 =  ( n4108 ) | ( n140 )  ;
assign n4113 =  ( ( n4108 ) * ( n140 ))  ;
assign n4114 =  ( n148 ) ? ( n4113 ) : ( VREG_0_1 ) ;
assign n4115 =  ( n146 ) ? ( n4112 ) : ( n4114 ) ;
assign n4116 =  ( n144 ) ? ( n4111 ) : ( n4115 ) ;
assign n4117 =  ( n142 ) ? ( n4110 ) : ( n4116 ) ;
assign n4118 =  ( n10 ) ? ( n4109 ) : ( n4117 ) ;
assign n4119 =  ( n77 ) & ( n3069 )  ;
assign n4120 =  ( n77 ) & ( n3071 )  ;
assign n4121 =  ( n77 ) & ( n3073 )  ;
assign n4122 =  ( n77 ) & ( n3075 )  ;
assign n4123 =  ( n77 ) & ( n3077 )  ;
assign n4124 =  ( n77 ) & ( n3079 )  ;
assign n4125 =  ( n77 ) & ( n3081 )  ;
assign n4126 =  ( n77 ) & ( n3083 )  ;
assign n4127 =  ( n77 ) & ( n3085 )  ;
assign n4128 =  ( n77 ) & ( n3087 )  ;
assign n4129 =  ( n77 ) & ( n3089 )  ;
assign n4130 =  ( n77 ) & ( n3091 )  ;
assign n4131 =  ( n77 ) & ( n3093 )  ;
assign n4132 =  ( n77 ) & ( n3095 )  ;
assign n4133 =  ( n77 ) & ( n3097 )  ;
assign n4134 =  ( n77 ) & ( n3099 )  ;
assign n4135 =  ( n78 ) & ( n3069 )  ;
assign n4136 =  ( n78 ) & ( n3071 )  ;
assign n4137 =  ( n78 ) & ( n3073 )  ;
assign n4138 =  ( n78 ) & ( n3075 )  ;
assign n4139 =  ( n78 ) & ( n3077 )  ;
assign n4140 =  ( n78 ) & ( n3079 )  ;
assign n4141 =  ( n78 ) & ( n3081 )  ;
assign n4142 =  ( n78 ) & ( n3083 )  ;
assign n4143 =  ( n78 ) & ( n3085 )  ;
assign n4144 =  ( n78 ) & ( n3087 )  ;
assign n4145 =  ( n78 ) & ( n3089 )  ;
assign n4146 =  ( n78 ) & ( n3091 )  ;
assign n4147 =  ( n78 ) & ( n3093 )  ;
assign n4148 =  ( n78 ) & ( n3095 )  ;
assign n4149 =  ( n78 ) & ( n3097 )  ;
assign n4150 =  ( n78 ) & ( n3099 )  ;
assign n4151 =  ( n79 ) & ( n3069 )  ;
assign n4152 =  ( n79 ) & ( n3071 )  ;
assign n4153 =  ( n79 ) & ( n3073 )  ;
assign n4154 =  ( n79 ) & ( n3075 )  ;
assign n4155 =  ( n79 ) & ( n3077 )  ;
assign n4156 =  ( n79 ) & ( n3079 )  ;
assign n4157 =  ( n79 ) & ( n3081 )  ;
assign n4158 =  ( n79 ) & ( n3083 )  ;
assign n4159 =  ( n79 ) & ( n3085 )  ;
assign n4160 =  ( n79 ) & ( n3087 )  ;
assign n4161 =  ( n79 ) & ( n3089 )  ;
assign n4162 =  ( n79 ) & ( n3091 )  ;
assign n4163 =  ( n79 ) & ( n3093 )  ;
assign n4164 =  ( n79 ) & ( n3095 )  ;
assign n4165 =  ( n79 ) & ( n3097 )  ;
assign n4166 =  ( n79 ) & ( n3099 )  ;
assign n4167 =  ( n80 ) & ( n3069 )  ;
assign n4168 =  ( n80 ) & ( n3071 )  ;
assign n4169 =  ( n80 ) & ( n3073 )  ;
assign n4170 =  ( n80 ) & ( n3075 )  ;
assign n4171 =  ( n80 ) & ( n3077 )  ;
assign n4172 =  ( n80 ) & ( n3079 )  ;
assign n4173 =  ( n80 ) & ( n3081 )  ;
assign n4174 =  ( n80 ) & ( n3083 )  ;
assign n4175 =  ( n80 ) & ( n3085 )  ;
assign n4176 =  ( n80 ) & ( n3087 )  ;
assign n4177 =  ( n80 ) & ( n3089 )  ;
assign n4178 =  ( n80 ) & ( n3091 )  ;
assign n4179 =  ( n80 ) & ( n3093 )  ;
assign n4180 =  ( n80 ) & ( n3095 )  ;
assign n4181 =  ( n80 ) & ( n3097 )  ;
assign n4182 =  ( n80 ) & ( n3099 )  ;
assign n4183 =  ( n81 ) & ( n3069 )  ;
assign n4184 =  ( n81 ) & ( n3071 )  ;
assign n4185 =  ( n81 ) & ( n3073 )  ;
assign n4186 =  ( n81 ) & ( n3075 )  ;
assign n4187 =  ( n81 ) & ( n3077 )  ;
assign n4188 =  ( n81 ) & ( n3079 )  ;
assign n4189 =  ( n81 ) & ( n3081 )  ;
assign n4190 =  ( n81 ) & ( n3083 )  ;
assign n4191 =  ( n81 ) & ( n3085 )  ;
assign n4192 =  ( n81 ) & ( n3087 )  ;
assign n4193 =  ( n81 ) & ( n3089 )  ;
assign n4194 =  ( n81 ) & ( n3091 )  ;
assign n4195 =  ( n81 ) & ( n3093 )  ;
assign n4196 =  ( n81 ) & ( n3095 )  ;
assign n4197 =  ( n81 ) & ( n3097 )  ;
assign n4198 =  ( n81 ) & ( n3099 )  ;
assign n4199 =  ( n82 ) & ( n3069 )  ;
assign n4200 =  ( n82 ) & ( n3071 )  ;
assign n4201 =  ( n82 ) & ( n3073 )  ;
assign n4202 =  ( n82 ) & ( n3075 )  ;
assign n4203 =  ( n82 ) & ( n3077 )  ;
assign n4204 =  ( n82 ) & ( n3079 )  ;
assign n4205 =  ( n82 ) & ( n3081 )  ;
assign n4206 =  ( n82 ) & ( n3083 )  ;
assign n4207 =  ( n82 ) & ( n3085 )  ;
assign n4208 =  ( n82 ) & ( n3087 )  ;
assign n4209 =  ( n82 ) & ( n3089 )  ;
assign n4210 =  ( n82 ) & ( n3091 )  ;
assign n4211 =  ( n82 ) & ( n3093 )  ;
assign n4212 =  ( n82 ) & ( n3095 )  ;
assign n4213 =  ( n82 ) & ( n3097 )  ;
assign n4214 =  ( n82 ) & ( n3099 )  ;
assign n4215 =  ( n83 ) & ( n3069 )  ;
assign n4216 =  ( n83 ) & ( n3071 )  ;
assign n4217 =  ( n83 ) & ( n3073 )  ;
assign n4218 =  ( n83 ) & ( n3075 )  ;
assign n4219 =  ( n83 ) & ( n3077 )  ;
assign n4220 =  ( n83 ) & ( n3079 )  ;
assign n4221 =  ( n83 ) & ( n3081 )  ;
assign n4222 =  ( n83 ) & ( n3083 )  ;
assign n4223 =  ( n83 ) & ( n3085 )  ;
assign n4224 =  ( n83 ) & ( n3087 )  ;
assign n4225 =  ( n83 ) & ( n3089 )  ;
assign n4226 =  ( n83 ) & ( n3091 )  ;
assign n4227 =  ( n83 ) & ( n3093 )  ;
assign n4228 =  ( n83 ) & ( n3095 )  ;
assign n4229 =  ( n83 ) & ( n3097 )  ;
assign n4230 =  ( n83 ) & ( n3099 )  ;
assign n4231 =  ( n84 ) & ( n3069 )  ;
assign n4232 =  ( n84 ) & ( n3071 )  ;
assign n4233 =  ( n84 ) & ( n3073 )  ;
assign n4234 =  ( n84 ) & ( n3075 )  ;
assign n4235 =  ( n84 ) & ( n3077 )  ;
assign n4236 =  ( n84 ) & ( n3079 )  ;
assign n4237 =  ( n84 ) & ( n3081 )  ;
assign n4238 =  ( n84 ) & ( n3083 )  ;
assign n4239 =  ( n84 ) & ( n3085 )  ;
assign n4240 =  ( n84 ) & ( n3087 )  ;
assign n4241 =  ( n84 ) & ( n3089 )  ;
assign n4242 =  ( n84 ) & ( n3091 )  ;
assign n4243 =  ( n84 ) & ( n3093 )  ;
assign n4244 =  ( n84 ) & ( n3095 )  ;
assign n4245 =  ( n84 ) & ( n3097 )  ;
assign n4246 =  ( n84 ) & ( n3099 )  ;
assign n4247 =  ( n85 ) & ( n3069 )  ;
assign n4248 =  ( n85 ) & ( n3071 )  ;
assign n4249 =  ( n85 ) & ( n3073 )  ;
assign n4250 =  ( n85 ) & ( n3075 )  ;
assign n4251 =  ( n85 ) & ( n3077 )  ;
assign n4252 =  ( n85 ) & ( n3079 )  ;
assign n4253 =  ( n85 ) & ( n3081 )  ;
assign n4254 =  ( n85 ) & ( n3083 )  ;
assign n4255 =  ( n85 ) & ( n3085 )  ;
assign n4256 =  ( n85 ) & ( n3087 )  ;
assign n4257 =  ( n85 ) & ( n3089 )  ;
assign n4258 =  ( n85 ) & ( n3091 )  ;
assign n4259 =  ( n85 ) & ( n3093 )  ;
assign n4260 =  ( n85 ) & ( n3095 )  ;
assign n4261 =  ( n85 ) & ( n3097 )  ;
assign n4262 =  ( n85 ) & ( n3099 )  ;
assign n4263 =  ( n86 ) & ( n3069 )  ;
assign n4264 =  ( n86 ) & ( n3071 )  ;
assign n4265 =  ( n86 ) & ( n3073 )  ;
assign n4266 =  ( n86 ) & ( n3075 )  ;
assign n4267 =  ( n86 ) & ( n3077 )  ;
assign n4268 =  ( n86 ) & ( n3079 )  ;
assign n4269 =  ( n86 ) & ( n3081 )  ;
assign n4270 =  ( n86 ) & ( n3083 )  ;
assign n4271 =  ( n86 ) & ( n3085 )  ;
assign n4272 =  ( n86 ) & ( n3087 )  ;
assign n4273 =  ( n86 ) & ( n3089 )  ;
assign n4274 =  ( n86 ) & ( n3091 )  ;
assign n4275 =  ( n86 ) & ( n3093 )  ;
assign n4276 =  ( n86 ) & ( n3095 )  ;
assign n4277 =  ( n86 ) & ( n3097 )  ;
assign n4278 =  ( n86 ) & ( n3099 )  ;
assign n4279 =  ( n87 ) & ( n3069 )  ;
assign n4280 =  ( n87 ) & ( n3071 )  ;
assign n4281 =  ( n87 ) & ( n3073 )  ;
assign n4282 =  ( n87 ) & ( n3075 )  ;
assign n4283 =  ( n87 ) & ( n3077 )  ;
assign n4284 =  ( n87 ) & ( n3079 )  ;
assign n4285 =  ( n87 ) & ( n3081 )  ;
assign n4286 =  ( n87 ) & ( n3083 )  ;
assign n4287 =  ( n87 ) & ( n3085 )  ;
assign n4288 =  ( n87 ) & ( n3087 )  ;
assign n4289 =  ( n87 ) & ( n3089 )  ;
assign n4290 =  ( n87 ) & ( n3091 )  ;
assign n4291 =  ( n87 ) & ( n3093 )  ;
assign n4292 =  ( n87 ) & ( n3095 )  ;
assign n4293 =  ( n87 ) & ( n3097 )  ;
assign n4294 =  ( n87 ) & ( n3099 )  ;
assign n4295 =  ( n88 ) & ( n3069 )  ;
assign n4296 =  ( n88 ) & ( n3071 )  ;
assign n4297 =  ( n88 ) & ( n3073 )  ;
assign n4298 =  ( n88 ) & ( n3075 )  ;
assign n4299 =  ( n88 ) & ( n3077 )  ;
assign n4300 =  ( n88 ) & ( n3079 )  ;
assign n4301 =  ( n88 ) & ( n3081 )  ;
assign n4302 =  ( n88 ) & ( n3083 )  ;
assign n4303 =  ( n88 ) & ( n3085 )  ;
assign n4304 =  ( n88 ) & ( n3087 )  ;
assign n4305 =  ( n88 ) & ( n3089 )  ;
assign n4306 =  ( n88 ) & ( n3091 )  ;
assign n4307 =  ( n88 ) & ( n3093 )  ;
assign n4308 =  ( n88 ) & ( n3095 )  ;
assign n4309 =  ( n88 ) & ( n3097 )  ;
assign n4310 =  ( n88 ) & ( n3099 )  ;
assign n4311 =  ( n89 ) & ( n3069 )  ;
assign n4312 =  ( n89 ) & ( n3071 )  ;
assign n4313 =  ( n89 ) & ( n3073 )  ;
assign n4314 =  ( n89 ) & ( n3075 )  ;
assign n4315 =  ( n89 ) & ( n3077 )  ;
assign n4316 =  ( n89 ) & ( n3079 )  ;
assign n4317 =  ( n89 ) & ( n3081 )  ;
assign n4318 =  ( n89 ) & ( n3083 )  ;
assign n4319 =  ( n89 ) & ( n3085 )  ;
assign n4320 =  ( n89 ) & ( n3087 )  ;
assign n4321 =  ( n89 ) & ( n3089 )  ;
assign n4322 =  ( n89 ) & ( n3091 )  ;
assign n4323 =  ( n89 ) & ( n3093 )  ;
assign n4324 =  ( n89 ) & ( n3095 )  ;
assign n4325 =  ( n89 ) & ( n3097 )  ;
assign n4326 =  ( n89 ) & ( n3099 )  ;
assign n4327 =  ( n90 ) & ( n3069 )  ;
assign n4328 =  ( n90 ) & ( n3071 )  ;
assign n4329 =  ( n90 ) & ( n3073 )  ;
assign n4330 =  ( n90 ) & ( n3075 )  ;
assign n4331 =  ( n90 ) & ( n3077 )  ;
assign n4332 =  ( n90 ) & ( n3079 )  ;
assign n4333 =  ( n90 ) & ( n3081 )  ;
assign n4334 =  ( n90 ) & ( n3083 )  ;
assign n4335 =  ( n90 ) & ( n3085 )  ;
assign n4336 =  ( n90 ) & ( n3087 )  ;
assign n4337 =  ( n90 ) & ( n3089 )  ;
assign n4338 =  ( n90 ) & ( n3091 )  ;
assign n4339 =  ( n90 ) & ( n3093 )  ;
assign n4340 =  ( n90 ) & ( n3095 )  ;
assign n4341 =  ( n90 ) & ( n3097 )  ;
assign n4342 =  ( n90 ) & ( n3099 )  ;
assign n4343 =  ( n91 ) & ( n3069 )  ;
assign n4344 =  ( n91 ) & ( n3071 )  ;
assign n4345 =  ( n91 ) & ( n3073 )  ;
assign n4346 =  ( n91 ) & ( n3075 )  ;
assign n4347 =  ( n91 ) & ( n3077 )  ;
assign n4348 =  ( n91 ) & ( n3079 )  ;
assign n4349 =  ( n91 ) & ( n3081 )  ;
assign n4350 =  ( n91 ) & ( n3083 )  ;
assign n4351 =  ( n91 ) & ( n3085 )  ;
assign n4352 =  ( n91 ) & ( n3087 )  ;
assign n4353 =  ( n91 ) & ( n3089 )  ;
assign n4354 =  ( n91 ) & ( n3091 )  ;
assign n4355 =  ( n91 ) & ( n3093 )  ;
assign n4356 =  ( n91 ) & ( n3095 )  ;
assign n4357 =  ( n91 ) & ( n3097 )  ;
assign n4358 =  ( n91 ) & ( n3099 )  ;
assign n4359 =  ( n92 ) & ( n3069 )  ;
assign n4360 =  ( n92 ) & ( n3071 )  ;
assign n4361 =  ( n92 ) & ( n3073 )  ;
assign n4362 =  ( n92 ) & ( n3075 )  ;
assign n4363 =  ( n92 ) & ( n3077 )  ;
assign n4364 =  ( n92 ) & ( n3079 )  ;
assign n4365 =  ( n92 ) & ( n3081 )  ;
assign n4366 =  ( n92 ) & ( n3083 )  ;
assign n4367 =  ( n92 ) & ( n3085 )  ;
assign n4368 =  ( n92 ) & ( n3087 )  ;
assign n4369 =  ( n92 ) & ( n3089 )  ;
assign n4370 =  ( n92 ) & ( n3091 )  ;
assign n4371 =  ( n92 ) & ( n3093 )  ;
assign n4372 =  ( n92 ) & ( n3095 )  ;
assign n4373 =  ( n92 ) & ( n3097 )  ;
assign n4374 =  ( n92 ) & ( n3099 )  ;
assign n4375 =  ( n93 ) & ( n3069 )  ;
assign n4376 =  ( n93 ) & ( n3071 )  ;
assign n4377 =  ( n93 ) & ( n3073 )  ;
assign n4378 =  ( n93 ) & ( n3075 )  ;
assign n4379 =  ( n93 ) & ( n3077 )  ;
assign n4380 =  ( n93 ) & ( n3079 )  ;
assign n4381 =  ( n93 ) & ( n3081 )  ;
assign n4382 =  ( n93 ) & ( n3083 )  ;
assign n4383 =  ( n93 ) & ( n3085 )  ;
assign n4384 =  ( n93 ) & ( n3087 )  ;
assign n4385 =  ( n93 ) & ( n3089 )  ;
assign n4386 =  ( n93 ) & ( n3091 )  ;
assign n4387 =  ( n93 ) & ( n3093 )  ;
assign n4388 =  ( n93 ) & ( n3095 )  ;
assign n4389 =  ( n93 ) & ( n3097 )  ;
assign n4390 =  ( n93 ) & ( n3099 )  ;
assign n4391 =  ( n94 ) & ( n3069 )  ;
assign n4392 =  ( n94 ) & ( n3071 )  ;
assign n4393 =  ( n94 ) & ( n3073 )  ;
assign n4394 =  ( n94 ) & ( n3075 )  ;
assign n4395 =  ( n94 ) & ( n3077 )  ;
assign n4396 =  ( n94 ) & ( n3079 )  ;
assign n4397 =  ( n94 ) & ( n3081 )  ;
assign n4398 =  ( n94 ) & ( n3083 )  ;
assign n4399 =  ( n94 ) & ( n3085 )  ;
assign n4400 =  ( n94 ) & ( n3087 )  ;
assign n4401 =  ( n94 ) & ( n3089 )  ;
assign n4402 =  ( n94 ) & ( n3091 )  ;
assign n4403 =  ( n94 ) & ( n3093 )  ;
assign n4404 =  ( n94 ) & ( n3095 )  ;
assign n4405 =  ( n94 ) & ( n3097 )  ;
assign n4406 =  ( n94 ) & ( n3099 )  ;
assign n4407 =  ( n95 ) & ( n3069 )  ;
assign n4408 =  ( n95 ) & ( n3071 )  ;
assign n4409 =  ( n95 ) & ( n3073 )  ;
assign n4410 =  ( n95 ) & ( n3075 )  ;
assign n4411 =  ( n95 ) & ( n3077 )  ;
assign n4412 =  ( n95 ) & ( n3079 )  ;
assign n4413 =  ( n95 ) & ( n3081 )  ;
assign n4414 =  ( n95 ) & ( n3083 )  ;
assign n4415 =  ( n95 ) & ( n3085 )  ;
assign n4416 =  ( n95 ) & ( n3087 )  ;
assign n4417 =  ( n95 ) & ( n3089 )  ;
assign n4418 =  ( n95 ) & ( n3091 )  ;
assign n4419 =  ( n95 ) & ( n3093 )  ;
assign n4420 =  ( n95 ) & ( n3095 )  ;
assign n4421 =  ( n95 ) & ( n3097 )  ;
assign n4422 =  ( n95 ) & ( n3099 )  ;
assign n4423 =  ( n96 ) & ( n3069 )  ;
assign n4424 =  ( n96 ) & ( n3071 )  ;
assign n4425 =  ( n96 ) & ( n3073 )  ;
assign n4426 =  ( n96 ) & ( n3075 )  ;
assign n4427 =  ( n96 ) & ( n3077 )  ;
assign n4428 =  ( n96 ) & ( n3079 )  ;
assign n4429 =  ( n96 ) & ( n3081 )  ;
assign n4430 =  ( n96 ) & ( n3083 )  ;
assign n4431 =  ( n96 ) & ( n3085 )  ;
assign n4432 =  ( n96 ) & ( n3087 )  ;
assign n4433 =  ( n96 ) & ( n3089 )  ;
assign n4434 =  ( n96 ) & ( n3091 )  ;
assign n4435 =  ( n96 ) & ( n3093 )  ;
assign n4436 =  ( n96 ) & ( n3095 )  ;
assign n4437 =  ( n96 ) & ( n3097 )  ;
assign n4438 =  ( n96 ) & ( n3099 )  ;
assign n4439 =  ( n97 ) & ( n3069 )  ;
assign n4440 =  ( n97 ) & ( n3071 )  ;
assign n4441 =  ( n97 ) & ( n3073 )  ;
assign n4442 =  ( n97 ) & ( n3075 )  ;
assign n4443 =  ( n97 ) & ( n3077 )  ;
assign n4444 =  ( n97 ) & ( n3079 )  ;
assign n4445 =  ( n97 ) & ( n3081 )  ;
assign n4446 =  ( n97 ) & ( n3083 )  ;
assign n4447 =  ( n97 ) & ( n3085 )  ;
assign n4448 =  ( n97 ) & ( n3087 )  ;
assign n4449 =  ( n97 ) & ( n3089 )  ;
assign n4450 =  ( n97 ) & ( n3091 )  ;
assign n4451 =  ( n97 ) & ( n3093 )  ;
assign n4452 =  ( n97 ) & ( n3095 )  ;
assign n4453 =  ( n97 ) & ( n3097 )  ;
assign n4454 =  ( n97 ) & ( n3099 )  ;
assign n4455 =  ( n98 ) & ( n3069 )  ;
assign n4456 =  ( n98 ) & ( n3071 )  ;
assign n4457 =  ( n98 ) & ( n3073 )  ;
assign n4458 =  ( n98 ) & ( n3075 )  ;
assign n4459 =  ( n98 ) & ( n3077 )  ;
assign n4460 =  ( n98 ) & ( n3079 )  ;
assign n4461 =  ( n98 ) & ( n3081 )  ;
assign n4462 =  ( n98 ) & ( n3083 )  ;
assign n4463 =  ( n98 ) & ( n3085 )  ;
assign n4464 =  ( n98 ) & ( n3087 )  ;
assign n4465 =  ( n98 ) & ( n3089 )  ;
assign n4466 =  ( n98 ) & ( n3091 )  ;
assign n4467 =  ( n98 ) & ( n3093 )  ;
assign n4468 =  ( n98 ) & ( n3095 )  ;
assign n4469 =  ( n98 ) & ( n3097 )  ;
assign n4470 =  ( n98 ) & ( n3099 )  ;
assign n4471 =  ( n99 ) & ( n3069 )  ;
assign n4472 =  ( n99 ) & ( n3071 )  ;
assign n4473 =  ( n99 ) & ( n3073 )  ;
assign n4474 =  ( n99 ) & ( n3075 )  ;
assign n4475 =  ( n99 ) & ( n3077 )  ;
assign n4476 =  ( n99 ) & ( n3079 )  ;
assign n4477 =  ( n99 ) & ( n3081 )  ;
assign n4478 =  ( n99 ) & ( n3083 )  ;
assign n4479 =  ( n99 ) & ( n3085 )  ;
assign n4480 =  ( n99 ) & ( n3087 )  ;
assign n4481 =  ( n99 ) & ( n3089 )  ;
assign n4482 =  ( n99 ) & ( n3091 )  ;
assign n4483 =  ( n99 ) & ( n3093 )  ;
assign n4484 =  ( n99 ) & ( n3095 )  ;
assign n4485 =  ( n99 ) & ( n3097 )  ;
assign n4486 =  ( n99 ) & ( n3099 )  ;
assign n4487 =  ( n100 ) & ( n3069 )  ;
assign n4488 =  ( n100 ) & ( n3071 )  ;
assign n4489 =  ( n100 ) & ( n3073 )  ;
assign n4490 =  ( n100 ) & ( n3075 )  ;
assign n4491 =  ( n100 ) & ( n3077 )  ;
assign n4492 =  ( n100 ) & ( n3079 )  ;
assign n4493 =  ( n100 ) & ( n3081 )  ;
assign n4494 =  ( n100 ) & ( n3083 )  ;
assign n4495 =  ( n100 ) & ( n3085 )  ;
assign n4496 =  ( n100 ) & ( n3087 )  ;
assign n4497 =  ( n100 ) & ( n3089 )  ;
assign n4498 =  ( n100 ) & ( n3091 )  ;
assign n4499 =  ( n100 ) & ( n3093 )  ;
assign n4500 =  ( n100 ) & ( n3095 )  ;
assign n4501 =  ( n100 ) & ( n3097 )  ;
assign n4502 =  ( n100 ) & ( n3099 )  ;
assign n4503 =  ( n101 ) & ( n3069 )  ;
assign n4504 =  ( n101 ) & ( n3071 )  ;
assign n4505 =  ( n101 ) & ( n3073 )  ;
assign n4506 =  ( n101 ) & ( n3075 )  ;
assign n4507 =  ( n101 ) & ( n3077 )  ;
assign n4508 =  ( n101 ) & ( n3079 )  ;
assign n4509 =  ( n101 ) & ( n3081 )  ;
assign n4510 =  ( n101 ) & ( n3083 )  ;
assign n4511 =  ( n101 ) & ( n3085 )  ;
assign n4512 =  ( n101 ) & ( n3087 )  ;
assign n4513 =  ( n101 ) & ( n3089 )  ;
assign n4514 =  ( n101 ) & ( n3091 )  ;
assign n4515 =  ( n101 ) & ( n3093 )  ;
assign n4516 =  ( n101 ) & ( n3095 )  ;
assign n4517 =  ( n101 ) & ( n3097 )  ;
assign n4518 =  ( n101 ) & ( n3099 )  ;
assign n4519 =  ( n102 ) & ( n3069 )  ;
assign n4520 =  ( n102 ) & ( n3071 )  ;
assign n4521 =  ( n102 ) & ( n3073 )  ;
assign n4522 =  ( n102 ) & ( n3075 )  ;
assign n4523 =  ( n102 ) & ( n3077 )  ;
assign n4524 =  ( n102 ) & ( n3079 )  ;
assign n4525 =  ( n102 ) & ( n3081 )  ;
assign n4526 =  ( n102 ) & ( n3083 )  ;
assign n4527 =  ( n102 ) & ( n3085 )  ;
assign n4528 =  ( n102 ) & ( n3087 )  ;
assign n4529 =  ( n102 ) & ( n3089 )  ;
assign n4530 =  ( n102 ) & ( n3091 )  ;
assign n4531 =  ( n102 ) & ( n3093 )  ;
assign n4532 =  ( n102 ) & ( n3095 )  ;
assign n4533 =  ( n102 ) & ( n3097 )  ;
assign n4534 =  ( n102 ) & ( n3099 )  ;
assign n4535 =  ( n103 ) & ( n3069 )  ;
assign n4536 =  ( n103 ) & ( n3071 )  ;
assign n4537 =  ( n103 ) & ( n3073 )  ;
assign n4538 =  ( n103 ) & ( n3075 )  ;
assign n4539 =  ( n103 ) & ( n3077 )  ;
assign n4540 =  ( n103 ) & ( n3079 )  ;
assign n4541 =  ( n103 ) & ( n3081 )  ;
assign n4542 =  ( n103 ) & ( n3083 )  ;
assign n4543 =  ( n103 ) & ( n3085 )  ;
assign n4544 =  ( n103 ) & ( n3087 )  ;
assign n4545 =  ( n103 ) & ( n3089 )  ;
assign n4546 =  ( n103 ) & ( n3091 )  ;
assign n4547 =  ( n103 ) & ( n3093 )  ;
assign n4548 =  ( n103 ) & ( n3095 )  ;
assign n4549 =  ( n103 ) & ( n3097 )  ;
assign n4550 =  ( n103 ) & ( n3099 )  ;
assign n4551 =  ( n104 ) & ( n3069 )  ;
assign n4552 =  ( n104 ) & ( n3071 )  ;
assign n4553 =  ( n104 ) & ( n3073 )  ;
assign n4554 =  ( n104 ) & ( n3075 )  ;
assign n4555 =  ( n104 ) & ( n3077 )  ;
assign n4556 =  ( n104 ) & ( n3079 )  ;
assign n4557 =  ( n104 ) & ( n3081 )  ;
assign n4558 =  ( n104 ) & ( n3083 )  ;
assign n4559 =  ( n104 ) & ( n3085 )  ;
assign n4560 =  ( n104 ) & ( n3087 )  ;
assign n4561 =  ( n104 ) & ( n3089 )  ;
assign n4562 =  ( n104 ) & ( n3091 )  ;
assign n4563 =  ( n104 ) & ( n3093 )  ;
assign n4564 =  ( n104 ) & ( n3095 )  ;
assign n4565 =  ( n104 ) & ( n3097 )  ;
assign n4566 =  ( n104 ) & ( n3099 )  ;
assign n4567 =  ( n105 ) & ( n3069 )  ;
assign n4568 =  ( n105 ) & ( n3071 )  ;
assign n4569 =  ( n105 ) & ( n3073 )  ;
assign n4570 =  ( n105 ) & ( n3075 )  ;
assign n4571 =  ( n105 ) & ( n3077 )  ;
assign n4572 =  ( n105 ) & ( n3079 )  ;
assign n4573 =  ( n105 ) & ( n3081 )  ;
assign n4574 =  ( n105 ) & ( n3083 )  ;
assign n4575 =  ( n105 ) & ( n3085 )  ;
assign n4576 =  ( n105 ) & ( n3087 )  ;
assign n4577 =  ( n105 ) & ( n3089 )  ;
assign n4578 =  ( n105 ) & ( n3091 )  ;
assign n4579 =  ( n105 ) & ( n3093 )  ;
assign n4580 =  ( n105 ) & ( n3095 )  ;
assign n4581 =  ( n105 ) & ( n3097 )  ;
assign n4582 =  ( n105 ) & ( n3099 )  ;
assign n4583 =  ( n106 ) & ( n3069 )  ;
assign n4584 =  ( n106 ) & ( n3071 )  ;
assign n4585 =  ( n106 ) & ( n3073 )  ;
assign n4586 =  ( n106 ) & ( n3075 )  ;
assign n4587 =  ( n106 ) & ( n3077 )  ;
assign n4588 =  ( n106 ) & ( n3079 )  ;
assign n4589 =  ( n106 ) & ( n3081 )  ;
assign n4590 =  ( n106 ) & ( n3083 )  ;
assign n4591 =  ( n106 ) & ( n3085 )  ;
assign n4592 =  ( n106 ) & ( n3087 )  ;
assign n4593 =  ( n106 ) & ( n3089 )  ;
assign n4594 =  ( n106 ) & ( n3091 )  ;
assign n4595 =  ( n106 ) & ( n3093 )  ;
assign n4596 =  ( n106 ) & ( n3095 )  ;
assign n4597 =  ( n106 ) & ( n3097 )  ;
assign n4598 =  ( n106 ) & ( n3099 )  ;
assign n4599 =  ( n107 ) & ( n3069 )  ;
assign n4600 =  ( n107 ) & ( n3071 )  ;
assign n4601 =  ( n107 ) & ( n3073 )  ;
assign n4602 =  ( n107 ) & ( n3075 )  ;
assign n4603 =  ( n107 ) & ( n3077 )  ;
assign n4604 =  ( n107 ) & ( n3079 )  ;
assign n4605 =  ( n107 ) & ( n3081 )  ;
assign n4606 =  ( n107 ) & ( n3083 )  ;
assign n4607 =  ( n107 ) & ( n3085 )  ;
assign n4608 =  ( n107 ) & ( n3087 )  ;
assign n4609 =  ( n107 ) & ( n3089 )  ;
assign n4610 =  ( n107 ) & ( n3091 )  ;
assign n4611 =  ( n107 ) & ( n3093 )  ;
assign n4612 =  ( n107 ) & ( n3095 )  ;
assign n4613 =  ( n107 ) & ( n3097 )  ;
assign n4614 =  ( n107 ) & ( n3099 )  ;
assign n4615 =  ( n108 ) & ( n3069 )  ;
assign n4616 =  ( n108 ) & ( n3071 )  ;
assign n4617 =  ( n108 ) & ( n3073 )  ;
assign n4618 =  ( n108 ) & ( n3075 )  ;
assign n4619 =  ( n108 ) & ( n3077 )  ;
assign n4620 =  ( n108 ) & ( n3079 )  ;
assign n4621 =  ( n108 ) & ( n3081 )  ;
assign n4622 =  ( n108 ) & ( n3083 )  ;
assign n4623 =  ( n108 ) & ( n3085 )  ;
assign n4624 =  ( n108 ) & ( n3087 )  ;
assign n4625 =  ( n108 ) & ( n3089 )  ;
assign n4626 =  ( n108 ) & ( n3091 )  ;
assign n4627 =  ( n108 ) & ( n3093 )  ;
assign n4628 =  ( n108 ) & ( n3095 )  ;
assign n4629 =  ( n108 ) & ( n3097 )  ;
assign n4630 =  ( n108 ) & ( n3099 )  ;
assign n4631 =  ( n4630 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n4632 =  ( n4629 ) ? ( VREG_0_1 ) : ( n4631 ) ;
assign n4633 =  ( n4628 ) ? ( VREG_0_2 ) : ( n4632 ) ;
assign n4634 =  ( n4627 ) ? ( VREG_0_3 ) : ( n4633 ) ;
assign n4635 =  ( n4626 ) ? ( VREG_0_4 ) : ( n4634 ) ;
assign n4636 =  ( n4625 ) ? ( VREG_0_5 ) : ( n4635 ) ;
assign n4637 =  ( n4624 ) ? ( VREG_0_6 ) : ( n4636 ) ;
assign n4638 =  ( n4623 ) ? ( VREG_0_7 ) : ( n4637 ) ;
assign n4639 =  ( n4622 ) ? ( VREG_0_8 ) : ( n4638 ) ;
assign n4640 =  ( n4621 ) ? ( VREG_0_9 ) : ( n4639 ) ;
assign n4641 =  ( n4620 ) ? ( VREG_0_10 ) : ( n4640 ) ;
assign n4642 =  ( n4619 ) ? ( VREG_0_11 ) : ( n4641 ) ;
assign n4643 =  ( n4618 ) ? ( VREG_0_12 ) : ( n4642 ) ;
assign n4644 =  ( n4617 ) ? ( VREG_0_13 ) : ( n4643 ) ;
assign n4645 =  ( n4616 ) ? ( VREG_0_14 ) : ( n4644 ) ;
assign n4646 =  ( n4615 ) ? ( VREG_0_15 ) : ( n4645 ) ;
assign n4647 =  ( n4614 ) ? ( VREG_1_0 ) : ( n4646 ) ;
assign n4648 =  ( n4613 ) ? ( VREG_1_1 ) : ( n4647 ) ;
assign n4649 =  ( n4612 ) ? ( VREG_1_2 ) : ( n4648 ) ;
assign n4650 =  ( n4611 ) ? ( VREG_1_3 ) : ( n4649 ) ;
assign n4651 =  ( n4610 ) ? ( VREG_1_4 ) : ( n4650 ) ;
assign n4652 =  ( n4609 ) ? ( VREG_1_5 ) : ( n4651 ) ;
assign n4653 =  ( n4608 ) ? ( VREG_1_6 ) : ( n4652 ) ;
assign n4654 =  ( n4607 ) ? ( VREG_1_7 ) : ( n4653 ) ;
assign n4655 =  ( n4606 ) ? ( VREG_1_8 ) : ( n4654 ) ;
assign n4656 =  ( n4605 ) ? ( VREG_1_9 ) : ( n4655 ) ;
assign n4657 =  ( n4604 ) ? ( VREG_1_10 ) : ( n4656 ) ;
assign n4658 =  ( n4603 ) ? ( VREG_1_11 ) : ( n4657 ) ;
assign n4659 =  ( n4602 ) ? ( VREG_1_12 ) : ( n4658 ) ;
assign n4660 =  ( n4601 ) ? ( VREG_1_13 ) : ( n4659 ) ;
assign n4661 =  ( n4600 ) ? ( VREG_1_14 ) : ( n4660 ) ;
assign n4662 =  ( n4599 ) ? ( VREG_1_15 ) : ( n4661 ) ;
assign n4663 =  ( n4598 ) ? ( VREG_2_0 ) : ( n4662 ) ;
assign n4664 =  ( n4597 ) ? ( VREG_2_1 ) : ( n4663 ) ;
assign n4665 =  ( n4596 ) ? ( VREG_2_2 ) : ( n4664 ) ;
assign n4666 =  ( n4595 ) ? ( VREG_2_3 ) : ( n4665 ) ;
assign n4667 =  ( n4594 ) ? ( VREG_2_4 ) : ( n4666 ) ;
assign n4668 =  ( n4593 ) ? ( VREG_2_5 ) : ( n4667 ) ;
assign n4669 =  ( n4592 ) ? ( VREG_2_6 ) : ( n4668 ) ;
assign n4670 =  ( n4591 ) ? ( VREG_2_7 ) : ( n4669 ) ;
assign n4671 =  ( n4590 ) ? ( VREG_2_8 ) : ( n4670 ) ;
assign n4672 =  ( n4589 ) ? ( VREG_2_9 ) : ( n4671 ) ;
assign n4673 =  ( n4588 ) ? ( VREG_2_10 ) : ( n4672 ) ;
assign n4674 =  ( n4587 ) ? ( VREG_2_11 ) : ( n4673 ) ;
assign n4675 =  ( n4586 ) ? ( VREG_2_12 ) : ( n4674 ) ;
assign n4676 =  ( n4585 ) ? ( VREG_2_13 ) : ( n4675 ) ;
assign n4677 =  ( n4584 ) ? ( VREG_2_14 ) : ( n4676 ) ;
assign n4678 =  ( n4583 ) ? ( VREG_2_15 ) : ( n4677 ) ;
assign n4679 =  ( n4582 ) ? ( VREG_3_0 ) : ( n4678 ) ;
assign n4680 =  ( n4581 ) ? ( VREG_3_1 ) : ( n4679 ) ;
assign n4681 =  ( n4580 ) ? ( VREG_3_2 ) : ( n4680 ) ;
assign n4682 =  ( n4579 ) ? ( VREG_3_3 ) : ( n4681 ) ;
assign n4683 =  ( n4578 ) ? ( VREG_3_4 ) : ( n4682 ) ;
assign n4684 =  ( n4577 ) ? ( VREG_3_5 ) : ( n4683 ) ;
assign n4685 =  ( n4576 ) ? ( VREG_3_6 ) : ( n4684 ) ;
assign n4686 =  ( n4575 ) ? ( VREG_3_7 ) : ( n4685 ) ;
assign n4687 =  ( n4574 ) ? ( VREG_3_8 ) : ( n4686 ) ;
assign n4688 =  ( n4573 ) ? ( VREG_3_9 ) : ( n4687 ) ;
assign n4689 =  ( n4572 ) ? ( VREG_3_10 ) : ( n4688 ) ;
assign n4690 =  ( n4571 ) ? ( VREG_3_11 ) : ( n4689 ) ;
assign n4691 =  ( n4570 ) ? ( VREG_3_12 ) : ( n4690 ) ;
assign n4692 =  ( n4569 ) ? ( VREG_3_13 ) : ( n4691 ) ;
assign n4693 =  ( n4568 ) ? ( VREG_3_14 ) : ( n4692 ) ;
assign n4694 =  ( n4567 ) ? ( VREG_3_15 ) : ( n4693 ) ;
assign n4695 =  ( n4566 ) ? ( VREG_4_0 ) : ( n4694 ) ;
assign n4696 =  ( n4565 ) ? ( VREG_4_1 ) : ( n4695 ) ;
assign n4697 =  ( n4564 ) ? ( VREG_4_2 ) : ( n4696 ) ;
assign n4698 =  ( n4563 ) ? ( VREG_4_3 ) : ( n4697 ) ;
assign n4699 =  ( n4562 ) ? ( VREG_4_4 ) : ( n4698 ) ;
assign n4700 =  ( n4561 ) ? ( VREG_4_5 ) : ( n4699 ) ;
assign n4701 =  ( n4560 ) ? ( VREG_4_6 ) : ( n4700 ) ;
assign n4702 =  ( n4559 ) ? ( VREG_4_7 ) : ( n4701 ) ;
assign n4703 =  ( n4558 ) ? ( VREG_4_8 ) : ( n4702 ) ;
assign n4704 =  ( n4557 ) ? ( VREG_4_9 ) : ( n4703 ) ;
assign n4705 =  ( n4556 ) ? ( VREG_4_10 ) : ( n4704 ) ;
assign n4706 =  ( n4555 ) ? ( VREG_4_11 ) : ( n4705 ) ;
assign n4707 =  ( n4554 ) ? ( VREG_4_12 ) : ( n4706 ) ;
assign n4708 =  ( n4553 ) ? ( VREG_4_13 ) : ( n4707 ) ;
assign n4709 =  ( n4552 ) ? ( VREG_4_14 ) : ( n4708 ) ;
assign n4710 =  ( n4551 ) ? ( VREG_4_15 ) : ( n4709 ) ;
assign n4711 =  ( n4550 ) ? ( VREG_5_0 ) : ( n4710 ) ;
assign n4712 =  ( n4549 ) ? ( VREG_5_1 ) : ( n4711 ) ;
assign n4713 =  ( n4548 ) ? ( VREG_5_2 ) : ( n4712 ) ;
assign n4714 =  ( n4547 ) ? ( VREG_5_3 ) : ( n4713 ) ;
assign n4715 =  ( n4546 ) ? ( VREG_5_4 ) : ( n4714 ) ;
assign n4716 =  ( n4545 ) ? ( VREG_5_5 ) : ( n4715 ) ;
assign n4717 =  ( n4544 ) ? ( VREG_5_6 ) : ( n4716 ) ;
assign n4718 =  ( n4543 ) ? ( VREG_5_7 ) : ( n4717 ) ;
assign n4719 =  ( n4542 ) ? ( VREG_5_8 ) : ( n4718 ) ;
assign n4720 =  ( n4541 ) ? ( VREG_5_9 ) : ( n4719 ) ;
assign n4721 =  ( n4540 ) ? ( VREG_5_10 ) : ( n4720 ) ;
assign n4722 =  ( n4539 ) ? ( VREG_5_11 ) : ( n4721 ) ;
assign n4723 =  ( n4538 ) ? ( VREG_5_12 ) : ( n4722 ) ;
assign n4724 =  ( n4537 ) ? ( VREG_5_13 ) : ( n4723 ) ;
assign n4725 =  ( n4536 ) ? ( VREG_5_14 ) : ( n4724 ) ;
assign n4726 =  ( n4535 ) ? ( VREG_5_15 ) : ( n4725 ) ;
assign n4727 =  ( n4534 ) ? ( VREG_6_0 ) : ( n4726 ) ;
assign n4728 =  ( n4533 ) ? ( VREG_6_1 ) : ( n4727 ) ;
assign n4729 =  ( n4532 ) ? ( VREG_6_2 ) : ( n4728 ) ;
assign n4730 =  ( n4531 ) ? ( VREG_6_3 ) : ( n4729 ) ;
assign n4731 =  ( n4530 ) ? ( VREG_6_4 ) : ( n4730 ) ;
assign n4732 =  ( n4529 ) ? ( VREG_6_5 ) : ( n4731 ) ;
assign n4733 =  ( n4528 ) ? ( VREG_6_6 ) : ( n4732 ) ;
assign n4734 =  ( n4527 ) ? ( VREG_6_7 ) : ( n4733 ) ;
assign n4735 =  ( n4526 ) ? ( VREG_6_8 ) : ( n4734 ) ;
assign n4736 =  ( n4525 ) ? ( VREG_6_9 ) : ( n4735 ) ;
assign n4737 =  ( n4524 ) ? ( VREG_6_10 ) : ( n4736 ) ;
assign n4738 =  ( n4523 ) ? ( VREG_6_11 ) : ( n4737 ) ;
assign n4739 =  ( n4522 ) ? ( VREG_6_12 ) : ( n4738 ) ;
assign n4740 =  ( n4521 ) ? ( VREG_6_13 ) : ( n4739 ) ;
assign n4741 =  ( n4520 ) ? ( VREG_6_14 ) : ( n4740 ) ;
assign n4742 =  ( n4519 ) ? ( VREG_6_15 ) : ( n4741 ) ;
assign n4743 =  ( n4518 ) ? ( VREG_7_0 ) : ( n4742 ) ;
assign n4744 =  ( n4517 ) ? ( VREG_7_1 ) : ( n4743 ) ;
assign n4745 =  ( n4516 ) ? ( VREG_7_2 ) : ( n4744 ) ;
assign n4746 =  ( n4515 ) ? ( VREG_7_3 ) : ( n4745 ) ;
assign n4747 =  ( n4514 ) ? ( VREG_7_4 ) : ( n4746 ) ;
assign n4748 =  ( n4513 ) ? ( VREG_7_5 ) : ( n4747 ) ;
assign n4749 =  ( n4512 ) ? ( VREG_7_6 ) : ( n4748 ) ;
assign n4750 =  ( n4511 ) ? ( VREG_7_7 ) : ( n4749 ) ;
assign n4751 =  ( n4510 ) ? ( VREG_7_8 ) : ( n4750 ) ;
assign n4752 =  ( n4509 ) ? ( VREG_7_9 ) : ( n4751 ) ;
assign n4753 =  ( n4508 ) ? ( VREG_7_10 ) : ( n4752 ) ;
assign n4754 =  ( n4507 ) ? ( VREG_7_11 ) : ( n4753 ) ;
assign n4755 =  ( n4506 ) ? ( VREG_7_12 ) : ( n4754 ) ;
assign n4756 =  ( n4505 ) ? ( VREG_7_13 ) : ( n4755 ) ;
assign n4757 =  ( n4504 ) ? ( VREG_7_14 ) : ( n4756 ) ;
assign n4758 =  ( n4503 ) ? ( VREG_7_15 ) : ( n4757 ) ;
assign n4759 =  ( n4502 ) ? ( VREG_8_0 ) : ( n4758 ) ;
assign n4760 =  ( n4501 ) ? ( VREG_8_1 ) : ( n4759 ) ;
assign n4761 =  ( n4500 ) ? ( VREG_8_2 ) : ( n4760 ) ;
assign n4762 =  ( n4499 ) ? ( VREG_8_3 ) : ( n4761 ) ;
assign n4763 =  ( n4498 ) ? ( VREG_8_4 ) : ( n4762 ) ;
assign n4764 =  ( n4497 ) ? ( VREG_8_5 ) : ( n4763 ) ;
assign n4765 =  ( n4496 ) ? ( VREG_8_6 ) : ( n4764 ) ;
assign n4766 =  ( n4495 ) ? ( VREG_8_7 ) : ( n4765 ) ;
assign n4767 =  ( n4494 ) ? ( VREG_8_8 ) : ( n4766 ) ;
assign n4768 =  ( n4493 ) ? ( VREG_8_9 ) : ( n4767 ) ;
assign n4769 =  ( n4492 ) ? ( VREG_8_10 ) : ( n4768 ) ;
assign n4770 =  ( n4491 ) ? ( VREG_8_11 ) : ( n4769 ) ;
assign n4771 =  ( n4490 ) ? ( VREG_8_12 ) : ( n4770 ) ;
assign n4772 =  ( n4489 ) ? ( VREG_8_13 ) : ( n4771 ) ;
assign n4773 =  ( n4488 ) ? ( VREG_8_14 ) : ( n4772 ) ;
assign n4774 =  ( n4487 ) ? ( VREG_8_15 ) : ( n4773 ) ;
assign n4775 =  ( n4486 ) ? ( VREG_9_0 ) : ( n4774 ) ;
assign n4776 =  ( n4485 ) ? ( VREG_9_1 ) : ( n4775 ) ;
assign n4777 =  ( n4484 ) ? ( VREG_9_2 ) : ( n4776 ) ;
assign n4778 =  ( n4483 ) ? ( VREG_9_3 ) : ( n4777 ) ;
assign n4779 =  ( n4482 ) ? ( VREG_9_4 ) : ( n4778 ) ;
assign n4780 =  ( n4481 ) ? ( VREG_9_5 ) : ( n4779 ) ;
assign n4781 =  ( n4480 ) ? ( VREG_9_6 ) : ( n4780 ) ;
assign n4782 =  ( n4479 ) ? ( VREG_9_7 ) : ( n4781 ) ;
assign n4783 =  ( n4478 ) ? ( VREG_9_8 ) : ( n4782 ) ;
assign n4784 =  ( n4477 ) ? ( VREG_9_9 ) : ( n4783 ) ;
assign n4785 =  ( n4476 ) ? ( VREG_9_10 ) : ( n4784 ) ;
assign n4786 =  ( n4475 ) ? ( VREG_9_11 ) : ( n4785 ) ;
assign n4787 =  ( n4474 ) ? ( VREG_9_12 ) : ( n4786 ) ;
assign n4788 =  ( n4473 ) ? ( VREG_9_13 ) : ( n4787 ) ;
assign n4789 =  ( n4472 ) ? ( VREG_9_14 ) : ( n4788 ) ;
assign n4790 =  ( n4471 ) ? ( VREG_9_15 ) : ( n4789 ) ;
assign n4791 =  ( n4470 ) ? ( VREG_10_0 ) : ( n4790 ) ;
assign n4792 =  ( n4469 ) ? ( VREG_10_1 ) : ( n4791 ) ;
assign n4793 =  ( n4468 ) ? ( VREG_10_2 ) : ( n4792 ) ;
assign n4794 =  ( n4467 ) ? ( VREG_10_3 ) : ( n4793 ) ;
assign n4795 =  ( n4466 ) ? ( VREG_10_4 ) : ( n4794 ) ;
assign n4796 =  ( n4465 ) ? ( VREG_10_5 ) : ( n4795 ) ;
assign n4797 =  ( n4464 ) ? ( VREG_10_6 ) : ( n4796 ) ;
assign n4798 =  ( n4463 ) ? ( VREG_10_7 ) : ( n4797 ) ;
assign n4799 =  ( n4462 ) ? ( VREG_10_8 ) : ( n4798 ) ;
assign n4800 =  ( n4461 ) ? ( VREG_10_9 ) : ( n4799 ) ;
assign n4801 =  ( n4460 ) ? ( VREG_10_10 ) : ( n4800 ) ;
assign n4802 =  ( n4459 ) ? ( VREG_10_11 ) : ( n4801 ) ;
assign n4803 =  ( n4458 ) ? ( VREG_10_12 ) : ( n4802 ) ;
assign n4804 =  ( n4457 ) ? ( VREG_10_13 ) : ( n4803 ) ;
assign n4805 =  ( n4456 ) ? ( VREG_10_14 ) : ( n4804 ) ;
assign n4806 =  ( n4455 ) ? ( VREG_10_15 ) : ( n4805 ) ;
assign n4807 =  ( n4454 ) ? ( VREG_11_0 ) : ( n4806 ) ;
assign n4808 =  ( n4453 ) ? ( VREG_11_1 ) : ( n4807 ) ;
assign n4809 =  ( n4452 ) ? ( VREG_11_2 ) : ( n4808 ) ;
assign n4810 =  ( n4451 ) ? ( VREG_11_3 ) : ( n4809 ) ;
assign n4811 =  ( n4450 ) ? ( VREG_11_4 ) : ( n4810 ) ;
assign n4812 =  ( n4449 ) ? ( VREG_11_5 ) : ( n4811 ) ;
assign n4813 =  ( n4448 ) ? ( VREG_11_6 ) : ( n4812 ) ;
assign n4814 =  ( n4447 ) ? ( VREG_11_7 ) : ( n4813 ) ;
assign n4815 =  ( n4446 ) ? ( VREG_11_8 ) : ( n4814 ) ;
assign n4816 =  ( n4445 ) ? ( VREG_11_9 ) : ( n4815 ) ;
assign n4817 =  ( n4444 ) ? ( VREG_11_10 ) : ( n4816 ) ;
assign n4818 =  ( n4443 ) ? ( VREG_11_11 ) : ( n4817 ) ;
assign n4819 =  ( n4442 ) ? ( VREG_11_12 ) : ( n4818 ) ;
assign n4820 =  ( n4441 ) ? ( VREG_11_13 ) : ( n4819 ) ;
assign n4821 =  ( n4440 ) ? ( VREG_11_14 ) : ( n4820 ) ;
assign n4822 =  ( n4439 ) ? ( VREG_11_15 ) : ( n4821 ) ;
assign n4823 =  ( n4438 ) ? ( VREG_12_0 ) : ( n4822 ) ;
assign n4824 =  ( n4437 ) ? ( VREG_12_1 ) : ( n4823 ) ;
assign n4825 =  ( n4436 ) ? ( VREG_12_2 ) : ( n4824 ) ;
assign n4826 =  ( n4435 ) ? ( VREG_12_3 ) : ( n4825 ) ;
assign n4827 =  ( n4434 ) ? ( VREG_12_4 ) : ( n4826 ) ;
assign n4828 =  ( n4433 ) ? ( VREG_12_5 ) : ( n4827 ) ;
assign n4829 =  ( n4432 ) ? ( VREG_12_6 ) : ( n4828 ) ;
assign n4830 =  ( n4431 ) ? ( VREG_12_7 ) : ( n4829 ) ;
assign n4831 =  ( n4430 ) ? ( VREG_12_8 ) : ( n4830 ) ;
assign n4832 =  ( n4429 ) ? ( VREG_12_9 ) : ( n4831 ) ;
assign n4833 =  ( n4428 ) ? ( VREG_12_10 ) : ( n4832 ) ;
assign n4834 =  ( n4427 ) ? ( VREG_12_11 ) : ( n4833 ) ;
assign n4835 =  ( n4426 ) ? ( VREG_12_12 ) : ( n4834 ) ;
assign n4836 =  ( n4425 ) ? ( VREG_12_13 ) : ( n4835 ) ;
assign n4837 =  ( n4424 ) ? ( VREG_12_14 ) : ( n4836 ) ;
assign n4838 =  ( n4423 ) ? ( VREG_12_15 ) : ( n4837 ) ;
assign n4839 =  ( n4422 ) ? ( VREG_13_0 ) : ( n4838 ) ;
assign n4840 =  ( n4421 ) ? ( VREG_13_1 ) : ( n4839 ) ;
assign n4841 =  ( n4420 ) ? ( VREG_13_2 ) : ( n4840 ) ;
assign n4842 =  ( n4419 ) ? ( VREG_13_3 ) : ( n4841 ) ;
assign n4843 =  ( n4418 ) ? ( VREG_13_4 ) : ( n4842 ) ;
assign n4844 =  ( n4417 ) ? ( VREG_13_5 ) : ( n4843 ) ;
assign n4845 =  ( n4416 ) ? ( VREG_13_6 ) : ( n4844 ) ;
assign n4846 =  ( n4415 ) ? ( VREG_13_7 ) : ( n4845 ) ;
assign n4847 =  ( n4414 ) ? ( VREG_13_8 ) : ( n4846 ) ;
assign n4848 =  ( n4413 ) ? ( VREG_13_9 ) : ( n4847 ) ;
assign n4849 =  ( n4412 ) ? ( VREG_13_10 ) : ( n4848 ) ;
assign n4850 =  ( n4411 ) ? ( VREG_13_11 ) : ( n4849 ) ;
assign n4851 =  ( n4410 ) ? ( VREG_13_12 ) : ( n4850 ) ;
assign n4852 =  ( n4409 ) ? ( VREG_13_13 ) : ( n4851 ) ;
assign n4853 =  ( n4408 ) ? ( VREG_13_14 ) : ( n4852 ) ;
assign n4854 =  ( n4407 ) ? ( VREG_13_15 ) : ( n4853 ) ;
assign n4855 =  ( n4406 ) ? ( VREG_14_0 ) : ( n4854 ) ;
assign n4856 =  ( n4405 ) ? ( VREG_14_1 ) : ( n4855 ) ;
assign n4857 =  ( n4404 ) ? ( VREG_14_2 ) : ( n4856 ) ;
assign n4858 =  ( n4403 ) ? ( VREG_14_3 ) : ( n4857 ) ;
assign n4859 =  ( n4402 ) ? ( VREG_14_4 ) : ( n4858 ) ;
assign n4860 =  ( n4401 ) ? ( VREG_14_5 ) : ( n4859 ) ;
assign n4861 =  ( n4400 ) ? ( VREG_14_6 ) : ( n4860 ) ;
assign n4862 =  ( n4399 ) ? ( VREG_14_7 ) : ( n4861 ) ;
assign n4863 =  ( n4398 ) ? ( VREG_14_8 ) : ( n4862 ) ;
assign n4864 =  ( n4397 ) ? ( VREG_14_9 ) : ( n4863 ) ;
assign n4865 =  ( n4396 ) ? ( VREG_14_10 ) : ( n4864 ) ;
assign n4866 =  ( n4395 ) ? ( VREG_14_11 ) : ( n4865 ) ;
assign n4867 =  ( n4394 ) ? ( VREG_14_12 ) : ( n4866 ) ;
assign n4868 =  ( n4393 ) ? ( VREG_14_13 ) : ( n4867 ) ;
assign n4869 =  ( n4392 ) ? ( VREG_14_14 ) : ( n4868 ) ;
assign n4870 =  ( n4391 ) ? ( VREG_14_15 ) : ( n4869 ) ;
assign n4871 =  ( n4390 ) ? ( VREG_15_0 ) : ( n4870 ) ;
assign n4872 =  ( n4389 ) ? ( VREG_15_1 ) : ( n4871 ) ;
assign n4873 =  ( n4388 ) ? ( VREG_15_2 ) : ( n4872 ) ;
assign n4874 =  ( n4387 ) ? ( VREG_15_3 ) : ( n4873 ) ;
assign n4875 =  ( n4386 ) ? ( VREG_15_4 ) : ( n4874 ) ;
assign n4876 =  ( n4385 ) ? ( VREG_15_5 ) : ( n4875 ) ;
assign n4877 =  ( n4384 ) ? ( VREG_15_6 ) : ( n4876 ) ;
assign n4878 =  ( n4383 ) ? ( VREG_15_7 ) : ( n4877 ) ;
assign n4879 =  ( n4382 ) ? ( VREG_15_8 ) : ( n4878 ) ;
assign n4880 =  ( n4381 ) ? ( VREG_15_9 ) : ( n4879 ) ;
assign n4881 =  ( n4380 ) ? ( VREG_15_10 ) : ( n4880 ) ;
assign n4882 =  ( n4379 ) ? ( VREG_15_11 ) : ( n4881 ) ;
assign n4883 =  ( n4378 ) ? ( VREG_15_12 ) : ( n4882 ) ;
assign n4884 =  ( n4377 ) ? ( VREG_15_13 ) : ( n4883 ) ;
assign n4885 =  ( n4376 ) ? ( VREG_15_14 ) : ( n4884 ) ;
assign n4886 =  ( n4375 ) ? ( VREG_15_15 ) : ( n4885 ) ;
assign n4887 =  ( n4374 ) ? ( VREG_16_0 ) : ( n4886 ) ;
assign n4888 =  ( n4373 ) ? ( VREG_16_1 ) : ( n4887 ) ;
assign n4889 =  ( n4372 ) ? ( VREG_16_2 ) : ( n4888 ) ;
assign n4890 =  ( n4371 ) ? ( VREG_16_3 ) : ( n4889 ) ;
assign n4891 =  ( n4370 ) ? ( VREG_16_4 ) : ( n4890 ) ;
assign n4892 =  ( n4369 ) ? ( VREG_16_5 ) : ( n4891 ) ;
assign n4893 =  ( n4368 ) ? ( VREG_16_6 ) : ( n4892 ) ;
assign n4894 =  ( n4367 ) ? ( VREG_16_7 ) : ( n4893 ) ;
assign n4895 =  ( n4366 ) ? ( VREG_16_8 ) : ( n4894 ) ;
assign n4896 =  ( n4365 ) ? ( VREG_16_9 ) : ( n4895 ) ;
assign n4897 =  ( n4364 ) ? ( VREG_16_10 ) : ( n4896 ) ;
assign n4898 =  ( n4363 ) ? ( VREG_16_11 ) : ( n4897 ) ;
assign n4899 =  ( n4362 ) ? ( VREG_16_12 ) : ( n4898 ) ;
assign n4900 =  ( n4361 ) ? ( VREG_16_13 ) : ( n4899 ) ;
assign n4901 =  ( n4360 ) ? ( VREG_16_14 ) : ( n4900 ) ;
assign n4902 =  ( n4359 ) ? ( VREG_16_15 ) : ( n4901 ) ;
assign n4903 =  ( n4358 ) ? ( VREG_17_0 ) : ( n4902 ) ;
assign n4904 =  ( n4357 ) ? ( VREG_17_1 ) : ( n4903 ) ;
assign n4905 =  ( n4356 ) ? ( VREG_17_2 ) : ( n4904 ) ;
assign n4906 =  ( n4355 ) ? ( VREG_17_3 ) : ( n4905 ) ;
assign n4907 =  ( n4354 ) ? ( VREG_17_4 ) : ( n4906 ) ;
assign n4908 =  ( n4353 ) ? ( VREG_17_5 ) : ( n4907 ) ;
assign n4909 =  ( n4352 ) ? ( VREG_17_6 ) : ( n4908 ) ;
assign n4910 =  ( n4351 ) ? ( VREG_17_7 ) : ( n4909 ) ;
assign n4911 =  ( n4350 ) ? ( VREG_17_8 ) : ( n4910 ) ;
assign n4912 =  ( n4349 ) ? ( VREG_17_9 ) : ( n4911 ) ;
assign n4913 =  ( n4348 ) ? ( VREG_17_10 ) : ( n4912 ) ;
assign n4914 =  ( n4347 ) ? ( VREG_17_11 ) : ( n4913 ) ;
assign n4915 =  ( n4346 ) ? ( VREG_17_12 ) : ( n4914 ) ;
assign n4916 =  ( n4345 ) ? ( VREG_17_13 ) : ( n4915 ) ;
assign n4917 =  ( n4344 ) ? ( VREG_17_14 ) : ( n4916 ) ;
assign n4918 =  ( n4343 ) ? ( VREG_17_15 ) : ( n4917 ) ;
assign n4919 =  ( n4342 ) ? ( VREG_18_0 ) : ( n4918 ) ;
assign n4920 =  ( n4341 ) ? ( VREG_18_1 ) : ( n4919 ) ;
assign n4921 =  ( n4340 ) ? ( VREG_18_2 ) : ( n4920 ) ;
assign n4922 =  ( n4339 ) ? ( VREG_18_3 ) : ( n4921 ) ;
assign n4923 =  ( n4338 ) ? ( VREG_18_4 ) : ( n4922 ) ;
assign n4924 =  ( n4337 ) ? ( VREG_18_5 ) : ( n4923 ) ;
assign n4925 =  ( n4336 ) ? ( VREG_18_6 ) : ( n4924 ) ;
assign n4926 =  ( n4335 ) ? ( VREG_18_7 ) : ( n4925 ) ;
assign n4927 =  ( n4334 ) ? ( VREG_18_8 ) : ( n4926 ) ;
assign n4928 =  ( n4333 ) ? ( VREG_18_9 ) : ( n4927 ) ;
assign n4929 =  ( n4332 ) ? ( VREG_18_10 ) : ( n4928 ) ;
assign n4930 =  ( n4331 ) ? ( VREG_18_11 ) : ( n4929 ) ;
assign n4931 =  ( n4330 ) ? ( VREG_18_12 ) : ( n4930 ) ;
assign n4932 =  ( n4329 ) ? ( VREG_18_13 ) : ( n4931 ) ;
assign n4933 =  ( n4328 ) ? ( VREG_18_14 ) : ( n4932 ) ;
assign n4934 =  ( n4327 ) ? ( VREG_18_15 ) : ( n4933 ) ;
assign n4935 =  ( n4326 ) ? ( VREG_19_0 ) : ( n4934 ) ;
assign n4936 =  ( n4325 ) ? ( VREG_19_1 ) : ( n4935 ) ;
assign n4937 =  ( n4324 ) ? ( VREG_19_2 ) : ( n4936 ) ;
assign n4938 =  ( n4323 ) ? ( VREG_19_3 ) : ( n4937 ) ;
assign n4939 =  ( n4322 ) ? ( VREG_19_4 ) : ( n4938 ) ;
assign n4940 =  ( n4321 ) ? ( VREG_19_5 ) : ( n4939 ) ;
assign n4941 =  ( n4320 ) ? ( VREG_19_6 ) : ( n4940 ) ;
assign n4942 =  ( n4319 ) ? ( VREG_19_7 ) : ( n4941 ) ;
assign n4943 =  ( n4318 ) ? ( VREG_19_8 ) : ( n4942 ) ;
assign n4944 =  ( n4317 ) ? ( VREG_19_9 ) : ( n4943 ) ;
assign n4945 =  ( n4316 ) ? ( VREG_19_10 ) : ( n4944 ) ;
assign n4946 =  ( n4315 ) ? ( VREG_19_11 ) : ( n4945 ) ;
assign n4947 =  ( n4314 ) ? ( VREG_19_12 ) : ( n4946 ) ;
assign n4948 =  ( n4313 ) ? ( VREG_19_13 ) : ( n4947 ) ;
assign n4949 =  ( n4312 ) ? ( VREG_19_14 ) : ( n4948 ) ;
assign n4950 =  ( n4311 ) ? ( VREG_19_15 ) : ( n4949 ) ;
assign n4951 =  ( n4310 ) ? ( VREG_20_0 ) : ( n4950 ) ;
assign n4952 =  ( n4309 ) ? ( VREG_20_1 ) : ( n4951 ) ;
assign n4953 =  ( n4308 ) ? ( VREG_20_2 ) : ( n4952 ) ;
assign n4954 =  ( n4307 ) ? ( VREG_20_3 ) : ( n4953 ) ;
assign n4955 =  ( n4306 ) ? ( VREG_20_4 ) : ( n4954 ) ;
assign n4956 =  ( n4305 ) ? ( VREG_20_5 ) : ( n4955 ) ;
assign n4957 =  ( n4304 ) ? ( VREG_20_6 ) : ( n4956 ) ;
assign n4958 =  ( n4303 ) ? ( VREG_20_7 ) : ( n4957 ) ;
assign n4959 =  ( n4302 ) ? ( VREG_20_8 ) : ( n4958 ) ;
assign n4960 =  ( n4301 ) ? ( VREG_20_9 ) : ( n4959 ) ;
assign n4961 =  ( n4300 ) ? ( VREG_20_10 ) : ( n4960 ) ;
assign n4962 =  ( n4299 ) ? ( VREG_20_11 ) : ( n4961 ) ;
assign n4963 =  ( n4298 ) ? ( VREG_20_12 ) : ( n4962 ) ;
assign n4964 =  ( n4297 ) ? ( VREG_20_13 ) : ( n4963 ) ;
assign n4965 =  ( n4296 ) ? ( VREG_20_14 ) : ( n4964 ) ;
assign n4966 =  ( n4295 ) ? ( VREG_20_15 ) : ( n4965 ) ;
assign n4967 =  ( n4294 ) ? ( VREG_21_0 ) : ( n4966 ) ;
assign n4968 =  ( n4293 ) ? ( VREG_21_1 ) : ( n4967 ) ;
assign n4969 =  ( n4292 ) ? ( VREG_21_2 ) : ( n4968 ) ;
assign n4970 =  ( n4291 ) ? ( VREG_21_3 ) : ( n4969 ) ;
assign n4971 =  ( n4290 ) ? ( VREG_21_4 ) : ( n4970 ) ;
assign n4972 =  ( n4289 ) ? ( VREG_21_5 ) : ( n4971 ) ;
assign n4973 =  ( n4288 ) ? ( VREG_21_6 ) : ( n4972 ) ;
assign n4974 =  ( n4287 ) ? ( VREG_21_7 ) : ( n4973 ) ;
assign n4975 =  ( n4286 ) ? ( VREG_21_8 ) : ( n4974 ) ;
assign n4976 =  ( n4285 ) ? ( VREG_21_9 ) : ( n4975 ) ;
assign n4977 =  ( n4284 ) ? ( VREG_21_10 ) : ( n4976 ) ;
assign n4978 =  ( n4283 ) ? ( VREG_21_11 ) : ( n4977 ) ;
assign n4979 =  ( n4282 ) ? ( VREG_21_12 ) : ( n4978 ) ;
assign n4980 =  ( n4281 ) ? ( VREG_21_13 ) : ( n4979 ) ;
assign n4981 =  ( n4280 ) ? ( VREG_21_14 ) : ( n4980 ) ;
assign n4982 =  ( n4279 ) ? ( VREG_21_15 ) : ( n4981 ) ;
assign n4983 =  ( n4278 ) ? ( VREG_22_0 ) : ( n4982 ) ;
assign n4984 =  ( n4277 ) ? ( VREG_22_1 ) : ( n4983 ) ;
assign n4985 =  ( n4276 ) ? ( VREG_22_2 ) : ( n4984 ) ;
assign n4986 =  ( n4275 ) ? ( VREG_22_3 ) : ( n4985 ) ;
assign n4987 =  ( n4274 ) ? ( VREG_22_4 ) : ( n4986 ) ;
assign n4988 =  ( n4273 ) ? ( VREG_22_5 ) : ( n4987 ) ;
assign n4989 =  ( n4272 ) ? ( VREG_22_6 ) : ( n4988 ) ;
assign n4990 =  ( n4271 ) ? ( VREG_22_7 ) : ( n4989 ) ;
assign n4991 =  ( n4270 ) ? ( VREG_22_8 ) : ( n4990 ) ;
assign n4992 =  ( n4269 ) ? ( VREG_22_9 ) : ( n4991 ) ;
assign n4993 =  ( n4268 ) ? ( VREG_22_10 ) : ( n4992 ) ;
assign n4994 =  ( n4267 ) ? ( VREG_22_11 ) : ( n4993 ) ;
assign n4995 =  ( n4266 ) ? ( VREG_22_12 ) : ( n4994 ) ;
assign n4996 =  ( n4265 ) ? ( VREG_22_13 ) : ( n4995 ) ;
assign n4997 =  ( n4264 ) ? ( VREG_22_14 ) : ( n4996 ) ;
assign n4998 =  ( n4263 ) ? ( VREG_22_15 ) : ( n4997 ) ;
assign n4999 =  ( n4262 ) ? ( VREG_23_0 ) : ( n4998 ) ;
assign n5000 =  ( n4261 ) ? ( VREG_23_1 ) : ( n4999 ) ;
assign n5001 =  ( n4260 ) ? ( VREG_23_2 ) : ( n5000 ) ;
assign n5002 =  ( n4259 ) ? ( VREG_23_3 ) : ( n5001 ) ;
assign n5003 =  ( n4258 ) ? ( VREG_23_4 ) : ( n5002 ) ;
assign n5004 =  ( n4257 ) ? ( VREG_23_5 ) : ( n5003 ) ;
assign n5005 =  ( n4256 ) ? ( VREG_23_6 ) : ( n5004 ) ;
assign n5006 =  ( n4255 ) ? ( VREG_23_7 ) : ( n5005 ) ;
assign n5007 =  ( n4254 ) ? ( VREG_23_8 ) : ( n5006 ) ;
assign n5008 =  ( n4253 ) ? ( VREG_23_9 ) : ( n5007 ) ;
assign n5009 =  ( n4252 ) ? ( VREG_23_10 ) : ( n5008 ) ;
assign n5010 =  ( n4251 ) ? ( VREG_23_11 ) : ( n5009 ) ;
assign n5011 =  ( n4250 ) ? ( VREG_23_12 ) : ( n5010 ) ;
assign n5012 =  ( n4249 ) ? ( VREG_23_13 ) : ( n5011 ) ;
assign n5013 =  ( n4248 ) ? ( VREG_23_14 ) : ( n5012 ) ;
assign n5014 =  ( n4247 ) ? ( VREG_23_15 ) : ( n5013 ) ;
assign n5015 =  ( n4246 ) ? ( VREG_24_0 ) : ( n5014 ) ;
assign n5016 =  ( n4245 ) ? ( VREG_24_1 ) : ( n5015 ) ;
assign n5017 =  ( n4244 ) ? ( VREG_24_2 ) : ( n5016 ) ;
assign n5018 =  ( n4243 ) ? ( VREG_24_3 ) : ( n5017 ) ;
assign n5019 =  ( n4242 ) ? ( VREG_24_4 ) : ( n5018 ) ;
assign n5020 =  ( n4241 ) ? ( VREG_24_5 ) : ( n5019 ) ;
assign n5021 =  ( n4240 ) ? ( VREG_24_6 ) : ( n5020 ) ;
assign n5022 =  ( n4239 ) ? ( VREG_24_7 ) : ( n5021 ) ;
assign n5023 =  ( n4238 ) ? ( VREG_24_8 ) : ( n5022 ) ;
assign n5024 =  ( n4237 ) ? ( VREG_24_9 ) : ( n5023 ) ;
assign n5025 =  ( n4236 ) ? ( VREG_24_10 ) : ( n5024 ) ;
assign n5026 =  ( n4235 ) ? ( VREG_24_11 ) : ( n5025 ) ;
assign n5027 =  ( n4234 ) ? ( VREG_24_12 ) : ( n5026 ) ;
assign n5028 =  ( n4233 ) ? ( VREG_24_13 ) : ( n5027 ) ;
assign n5029 =  ( n4232 ) ? ( VREG_24_14 ) : ( n5028 ) ;
assign n5030 =  ( n4231 ) ? ( VREG_24_15 ) : ( n5029 ) ;
assign n5031 =  ( n4230 ) ? ( VREG_25_0 ) : ( n5030 ) ;
assign n5032 =  ( n4229 ) ? ( VREG_25_1 ) : ( n5031 ) ;
assign n5033 =  ( n4228 ) ? ( VREG_25_2 ) : ( n5032 ) ;
assign n5034 =  ( n4227 ) ? ( VREG_25_3 ) : ( n5033 ) ;
assign n5035 =  ( n4226 ) ? ( VREG_25_4 ) : ( n5034 ) ;
assign n5036 =  ( n4225 ) ? ( VREG_25_5 ) : ( n5035 ) ;
assign n5037 =  ( n4224 ) ? ( VREG_25_6 ) : ( n5036 ) ;
assign n5038 =  ( n4223 ) ? ( VREG_25_7 ) : ( n5037 ) ;
assign n5039 =  ( n4222 ) ? ( VREG_25_8 ) : ( n5038 ) ;
assign n5040 =  ( n4221 ) ? ( VREG_25_9 ) : ( n5039 ) ;
assign n5041 =  ( n4220 ) ? ( VREG_25_10 ) : ( n5040 ) ;
assign n5042 =  ( n4219 ) ? ( VREG_25_11 ) : ( n5041 ) ;
assign n5043 =  ( n4218 ) ? ( VREG_25_12 ) : ( n5042 ) ;
assign n5044 =  ( n4217 ) ? ( VREG_25_13 ) : ( n5043 ) ;
assign n5045 =  ( n4216 ) ? ( VREG_25_14 ) : ( n5044 ) ;
assign n5046 =  ( n4215 ) ? ( VREG_25_15 ) : ( n5045 ) ;
assign n5047 =  ( n4214 ) ? ( VREG_26_0 ) : ( n5046 ) ;
assign n5048 =  ( n4213 ) ? ( VREG_26_1 ) : ( n5047 ) ;
assign n5049 =  ( n4212 ) ? ( VREG_26_2 ) : ( n5048 ) ;
assign n5050 =  ( n4211 ) ? ( VREG_26_3 ) : ( n5049 ) ;
assign n5051 =  ( n4210 ) ? ( VREG_26_4 ) : ( n5050 ) ;
assign n5052 =  ( n4209 ) ? ( VREG_26_5 ) : ( n5051 ) ;
assign n5053 =  ( n4208 ) ? ( VREG_26_6 ) : ( n5052 ) ;
assign n5054 =  ( n4207 ) ? ( VREG_26_7 ) : ( n5053 ) ;
assign n5055 =  ( n4206 ) ? ( VREG_26_8 ) : ( n5054 ) ;
assign n5056 =  ( n4205 ) ? ( VREG_26_9 ) : ( n5055 ) ;
assign n5057 =  ( n4204 ) ? ( VREG_26_10 ) : ( n5056 ) ;
assign n5058 =  ( n4203 ) ? ( VREG_26_11 ) : ( n5057 ) ;
assign n5059 =  ( n4202 ) ? ( VREG_26_12 ) : ( n5058 ) ;
assign n5060 =  ( n4201 ) ? ( VREG_26_13 ) : ( n5059 ) ;
assign n5061 =  ( n4200 ) ? ( VREG_26_14 ) : ( n5060 ) ;
assign n5062 =  ( n4199 ) ? ( VREG_26_15 ) : ( n5061 ) ;
assign n5063 =  ( n4198 ) ? ( VREG_27_0 ) : ( n5062 ) ;
assign n5064 =  ( n4197 ) ? ( VREG_27_1 ) : ( n5063 ) ;
assign n5065 =  ( n4196 ) ? ( VREG_27_2 ) : ( n5064 ) ;
assign n5066 =  ( n4195 ) ? ( VREG_27_3 ) : ( n5065 ) ;
assign n5067 =  ( n4194 ) ? ( VREG_27_4 ) : ( n5066 ) ;
assign n5068 =  ( n4193 ) ? ( VREG_27_5 ) : ( n5067 ) ;
assign n5069 =  ( n4192 ) ? ( VREG_27_6 ) : ( n5068 ) ;
assign n5070 =  ( n4191 ) ? ( VREG_27_7 ) : ( n5069 ) ;
assign n5071 =  ( n4190 ) ? ( VREG_27_8 ) : ( n5070 ) ;
assign n5072 =  ( n4189 ) ? ( VREG_27_9 ) : ( n5071 ) ;
assign n5073 =  ( n4188 ) ? ( VREG_27_10 ) : ( n5072 ) ;
assign n5074 =  ( n4187 ) ? ( VREG_27_11 ) : ( n5073 ) ;
assign n5075 =  ( n4186 ) ? ( VREG_27_12 ) : ( n5074 ) ;
assign n5076 =  ( n4185 ) ? ( VREG_27_13 ) : ( n5075 ) ;
assign n5077 =  ( n4184 ) ? ( VREG_27_14 ) : ( n5076 ) ;
assign n5078 =  ( n4183 ) ? ( VREG_27_15 ) : ( n5077 ) ;
assign n5079 =  ( n4182 ) ? ( VREG_28_0 ) : ( n5078 ) ;
assign n5080 =  ( n4181 ) ? ( VREG_28_1 ) : ( n5079 ) ;
assign n5081 =  ( n4180 ) ? ( VREG_28_2 ) : ( n5080 ) ;
assign n5082 =  ( n4179 ) ? ( VREG_28_3 ) : ( n5081 ) ;
assign n5083 =  ( n4178 ) ? ( VREG_28_4 ) : ( n5082 ) ;
assign n5084 =  ( n4177 ) ? ( VREG_28_5 ) : ( n5083 ) ;
assign n5085 =  ( n4176 ) ? ( VREG_28_6 ) : ( n5084 ) ;
assign n5086 =  ( n4175 ) ? ( VREG_28_7 ) : ( n5085 ) ;
assign n5087 =  ( n4174 ) ? ( VREG_28_8 ) : ( n5086 ) ;
assign n5088 =  ( n4173 ) ? ( VREG_28_9 ) : ( n5087 ) ;
assign n5089 =  ( n4172 ) ? ( VREG_28_10 ) : ( n5088 ) ;
assign n5090 =  ( n4171 ) ? ( VREG_28_11 ) : ( n5089 ) ;
assign n5091 =  ( n4170 ) ? ( VREG_28_12 ) : ( n5090 ) ;
assign n5092 =  ( n4169 ) ? ( VREG_28_13 ) : ( n5091 ) ;
assign n5093 =  ( n4168 ) ? ( VREG_28_14 ) : ( n5092 ) ;
assign n5094 =  ( n4167 ) ? ( VREG_28_15 ) : ( n5093 ) ;
assign n5095 =  ( n4166 ) ? ( VREG_29_0 ) : ( n5094 ) ;
assign n5096 =  ( n4165 ) ? ( VREG_29_1 ) : ( n5095 ) ;
assign n5097 =  ( n4164 ) ? ( VREG_29_2 ) : ( n5096 ) ;
assign n5098 =  ( n4163 ) ? ( VREG_29_3 ) : ( n5097 ) ;
assign n5099 =  ( n4162 ) ? ( VREG_29_4 ) : ( n5098 ) ;
assign n5100 =  ( n4161 ) ? ( VREG_29_5 ) : ( n5099 ) ;
assign n5101 =  ( n4160 ) ? ( VREG_29_6 ) : ( n5100 ) ;
assign n5102 =  ( n4159 ) ? ( VREG_29_7 ) : ( n5101 ) ;
assign n5103 =  ( n4158 ) ? ( VREG_29_8 ) : ( n5102 ) ;
assign n5104 =  ( n4157 ) ? ( VREG_29_9 ) : ( n5103 ) ;
assign n5105 =  ( n4156 ) ? ( VREG_29_10 ) : ( n5104 ) ;
assign n5106 =  ( n4155 ) ? ( VREG_29_11 ) : ( n5105 ) ;
assign n5107 =  ( n4154 ) ? ( VREG_29_12 ) : ( n5106 ) ;
assign n5108 =  ( n4153 ) ? ( VREG_29_13 ) : ( n5107 ) ;
assign n5109 =  ( n4152 ) ? ( VREG_29_14 ) : ( n5108 ) ;
assign n5110 =  ( n4151 ) ? ( VREG_29_15 ) : ( n5109 ) ;
assign n5111 =  ( n4150 ) ? ( VREG_30_0 ) : ( n5110 ) ;
assign n5112 =  ( n4149 ) ? ( VREG_30_1 ) : ( n5111 ) ;
assign n5113 =  ( n4148 ) ? ( VREG_30_2 ) : ( n5112 ) ;
assign n5114 =  ( n4147 ) ? ( VREG_30_3 ) : ( n5113 ) ;
assign n5115 =  ( n4146 ) ? ( VREG_30_4 ) : ( n5114 ) ;
assign n5116 =  ( n4145 ) ? ( VREG_30_5 ) : ( n5115 ) ;
assign n5117 =  ( n4144 ) ? ( VREG_30_6 ) : ( n5116 ) ;
assign n5118 =  ( n4143 ) ? ( VREG_30_7 ) : ( n5117 ) ;
assign n5119 =  ( n4142 ) ? ( VREG_30_8 ) : ( n5118 ) ;
assign n5120 =  ( n4141 ) ? ( VREG_30_9 ) : ( n5119 ) ;
assign n5121 =  ( n4140 ) ? ( VREG_30_10 ) : ( n5120 ) ;
assign n5122 =  ( n4139 ) ? ( VREG_30_11 ) : ( n5121 ) ;
assign n5123 =  ( n4138 ) ? ( VREG_30_12 ) : ( n5122 ) ;
assign n5124 =  ( n4137 ) ? ( VREG_30_13 ) : ( n5123 ) ;
assign n5125 =  ( n4136 ) ? ( VREG_30_14 ) : ( n5124 ) ;
assign n5126 =  ( n4135 ) ? ( VREG_30_15 ) : ( n5125 ) ;
assign n5127 =  ( n4134 ) ? ( VREG_31_0 ) : ( n5126 ) ;
assign n5128 =  ( n4133 ) ? ( VREG_31_1 ) : ( n5127 ) ;
assign n5129 =  ( n4132 ) ? ( VREG_31_2 ) : ( n5128 ) ;
assign n5130 =  ( n4131 ) ? ( VREG_31_3 ) : ( n5129 ) ;
assign n5131 =  ( n4130 ) ? ( VREG_31_4 ) : ( n5130 ) ;
assign n5132 =  ( n4129 ) ? ( VREG_31_5 ) : ( n5131 ) ;
assign n5133 =  ( n4128 ) ? ( VREG_31_6 ) : ( n5132 ) ;
assign n5134 =  ( n4127 ) ? ( VREG_31_7 ) : ( n5133 ) ;
assign n5135 =  ( n4126 ) ? ( VREG_31_8 ) : ( n5134 ) ;
assign n5136 =  ( n4125 ) ? ( VREG_31_9 ) : ( n5135 ) ;
assign n5137 =  ( n4124 ) ? ( VREG_31_10 ) : ( n5136 ) ;
assign n5138 =  ( n4123 ) ? ( VREG_31_11 ) : ( n5137 ) ;
assign n5139 =  ( n4122 ) ? ( VREG_31_12 ) : ( n5138 ) ;
assign n5140 =  ( n4121 ) ? ( VREG_31_13 ) : ( n5139 ) ;
assign n5141 =  ( n4120 ) ? ( VREG_31_14 ) : ( n5140 ) ;
assign n5142 =  ( n4119 ) ? ( VREG_31_15 ) : ( n5141 ) ;
assign n5143 =  ( n4108 ) + ( n5142 )  ;
assign n5144 =  ( n4108 ) - ( n5142 )  ;
assign n5145 =  ( n4108 ) & ( n5142 )  ;
assign n5146 =  ( n4108 ) | ( n5142 )  ;
assign n5147 =  ( ( n4108 ) * ( n5142 ))  ;
assign n5148 =  ( n148 ) ? ( n5147 ) : ( VREG_0_1 ) ;
assign n5149 =  ( n146 ) ? ( n5146 ) : ( n5148 ) ;
assign n5150 =  ( n144 ) ? ( n5145 ) : ( n5149 ) ;
assign n5151 =  ( n142 ) ? ( n5144 ) : ( n5150 ) ;
assign n5152 =  ( n10 ) ? ( n5143 ) : ( n5151 ) ;
assign n5153 = n3030[1:1] ;
assign n5154 =  ( n5153 ) == ( 1'd0 )  ;
assign n5155 =  ( n5154 ) ? ( VREG_0_1 ) : ( n4118 ) ;
assign n5156 =  ( n5154 ) ? ( VREG_0_1 ) : ( n5152 ) ;
assign n5157 =  ( n3034 ) ? ( n5156 ) : ( VREG_0_1 ) ;
assign n5158 =  ( n2965 ) ? ( n5155 ) : ( n5157 ) ;
assign n5159 =  ( n1930 ) ? ( n5152 ) : ( n5158 ) ;
assign n5160 =  ( n879 ) ? ( n4118 ) : ( n5159 ) ;
assign n5161 =  ( n4108 ) + ( n164 )  ;
assign n5162 =  ( n4108 ) - ( n164 )  ;
assign n5163 =  ( n4108 ) & ( n164 )  ;
assign n5164 =  ( n4108 ) | ( n164 )  ;
assign n5165 =  ( ( n4108 ) * ( n164 ))  ;
assign n5166 =  ( n172 ) ? ( n5165 ) : ( VREG_0_1 ) ;
assign n5167 =  ( n170 ) ? ( n5164 ) : ( n5166 ) ;
assign n5168 =  ( n168 ) ? ( n5163 ) : ( n5167 ) ;
assign n5169 =  ( n166 ) ? ( n5162 ) : ( n5168 ) ;
assign n5170 =  ( n162 ) ? ( n5161 ) : ( n5169 ) ;
assign n5171 =  ( n4108 ) + ( n180 )  ;
assign n5172 =  ( n4108 ) - ( n180 )  ;
assign n5173 =  ( n4108 ) & ( n180 )  ;
assign n5174 =  ( n4108 ) | ( n180 )  ;
assign n5175 =  ( ( n4108 ) * ( n180 ))  ;
assign n5176 =  ( n172 ) ? ( n5175 ) : ( VREG_0_1 ) ;
assign n5177 =  ( n170 ) ? ( n5174 ) : ( n5176 ) ;
assign n5178 =  ( n168 ) ? ( n5173 ) : ( n5177 ) ;
assign n5179 =  ( n166 ) ? ( n5172 ) : ( n5178 ) ;
assign n5180 =  ( n162 ) ? ( n5171 ) : ( n5179 ) ;
assign n5181 =  ( n5154 ) ? ( VREG_0_1 ) : ( n5180 ) ;
assign n5182 =  ( n3051 ) ? ( n5181 ) : ( VREG_0_1 ) ;
assign n5183 =  ( n3040 ) ? ( n5170 ) : ( n5182 ) ;
assign n5184 =  ( n192 ) ? ( VREG_0_1 ) : ( VREG_0_1 ) ;
assign n5185 =  ( n157 ) ? ( n5183 ) : ( n5184 ) ;
assign n5186 =  ( n6 ) ? ( n5160 ) : ( n5185 ) ;
assign n5187 =  ( n4 ) ? ( n5186 ) : ( VREG_0_1 ) ;
assign n5188 =  ( 32'd10 ) == ( 32'd15 )  ;
assign n5189 =  ( n12 ) & ( n5188 )  ;
assign n5190 =  ( 32'd10 ) == ( 32'd14 )  ;
assign n5191 =  ( n12 ) & ( n5190 )  ;
assign n5192 =  ( 32'd10 ) == ( 32'd13 )  ;
assign n5193 =  ( n12 ) & ( n5192 )  ;
assign n5194 =  ( 32'd10 ) == ( 32'd12 )  ;
assign n5195 =  ( n12 ) & ( n5194 )  ;
assign n5196 =  ( 32'd10 ) == ( 32'd11 )  ;
assign n5197 =  ( n12 ) & ( n5196 )  ;
assign n5198 =  ( 32'd10 ) == ( 32'd10 )  ;
assign n5199 =  ( n12 ) & ( n5198 )  ;
assign n5200 =  ( 32'd10 ) == ( 32'd9 )  ;
assign n5201 =  ( n12 ) & ( n5200 )  ;
assign n5202 =  ( 32'd10 ) == ( 32'd8 )  ;
assign n5203 =  ( n12 ) & ( n5202 )  ;
assign n5204 =  ( 32'd10 ) == ( 32'd7 )  ;
assign n5205 =  ( n12 ) & ( n5204 )  ;
assign n5206 =  ( 32'd10 ) == ( 32'd6 )  ;
assign n5207 =  ( n12 ) & ( n5206 )  ;
assign n5208 =  ( 32'd10 ) == ( 32'd5 )  ;
assign n5209 =  ( n12 ) & ( n5208 )  ;
assign n5210 =  ( 32'd10 ) == ( 32'd4 )  ;
assign n5211 =  ( n12 ) & ( n5210 )  ;
assign n5212 =  ( 32'd10 ) == ( 32'd3 )  ;
assign n5213 =  ( n12 ) & ( n5212 )  ;
assign n5214 =  ( 32'd10 ) == ( 32'd2 )  ;
assign n5215 =  ( n12 ) & ( n5214 )  ;
assign n5216 =  ( 32'd10 ) == ( 32'd1 )  ;
assign n5217 =  ( n12 ) & ( n5216 )  ;
assign n5218 =  ( 32'd10 ) == ( 32'd0 )  ;
assign n5219 =  ( n12 ) & ( n5218 )  ;
assign n5220 =  ( n13 ) & ( n5188 )  ;
assign n5221 =  ( n13 ) & ( n5190 )  ;
assign n5222 =  ( n13 ) & ( n5192 )  ;
assign n5223 =  ( n13 ) & ( n5194 )  ;
assign n5224 =  ( n13 ) & ( n5196 )  ;
assign n5225 =  ( n13 ) & ( n5198 )  ;
assign n5226 =  ( n13 ) & ( n5200 )  ;
assign n5227 =  ( n13 ) & ( n5202 )  ;
assign n5228 =  ( n13 ) & ( n5204 )  ;
assign n5229 =  ( n13 ) & ( n5206 )  ;
assign n5230 =  ( n13 ) & ( n5208 )  ;
assign n5231 =  ( n13 ) & ( n5210 )  ;
assign n5232 =  ( n13 ) & ( n5212 )  ;
assign n5233 =  ( n13 ) & ( n5214 )  ;
assign n5234 =  ( n13 ) & ( n5216 )  ;
assign n5235 =  ( n13 ) & ( n5218 )  ;
assign n5236 =  ( n14 ) & ( n5188 )  ;
assign n5237 =  ( n14 ) & ( n5190 )  ;
assign n5238 =  ( n14 ) & ( n5192 )  ;
assign n5239 =  ( n14 ) & ( n5194 )  ;
assign n5240 =  ( n14 ) & ( n5196 )  ;
assign n5241 =  ( n14 ) & ( n5198 )  ;
assign n5242 =  ( n14 ) & ( n5200 )  ;
assign n5243 =  ( n14 ) & ( n5202 )  ;
assign n5244 =  ( n14 ) & ( n5204 )  ;
assign n5245 =  ( n14 ) & ( n5206 )  ;
assign n5246 =  ( n14 ) & ( n5208 )  ;
assign n5247 =  ( n14 ) & ( n5210 )  ;
assign n5248 =  ( n14 ) & ( n5212 )  ;
assign n5249 =  ( n14 ) & ( n5214 )  ;
assign n5250 =  ( n14 ) & ( n5216 )  ;
assign n5251 =  ( n14 ) & ( n5218 )  ;
assign n5252 =  ( n15 ) & ( n5188 )  ;
assign n5253 =  ( n15 ) & ( n5190 )  ;
assign n5254 =  ( n15 ) & ( n5192 )  ;
assign n5255 =  ( n15 ) & ( n5194 )  ;
assign n5256 =  ( n15 ) & ( n5196 )  ;
assign n5257 =  ( n15 ) & ( n5198 )  ;
assign n5258 =  ( n15 ) & ( n5200 )  ;
assign n5259 =  ( n15 ) & ( n5202 )  ;
assign n5260 =  ( n15 ) & ( n5204 )  ;
assign n5261 =  ( n15 ) & ( n5206 )  ;
assign n5262 =  ( n15 ) & ( n5208 )  ;
assign n5263 =  ( n15 ) & ( n5210 )  ;
assign n5264 =  ( n15 ) & ( n5212 )  ;
assign n5265 =  ( n15 ) & ( n5214 )  ;
assign n5266 =  ( n15 ) & ( n5216 )  ;
assign n5267 =  ( n15 ) & ( n5218 )  ;
assign n5268 =  ( n16 ) & ( n5188 )  ;
assign n5269 =  ( n16 ) & ( n5190 )  ;
assign n5270 =  ( n16 ) & ( n5192 )  ;
assign n5271 =  ( n16 ) & ( n5194 )  ;
assign n5272 =  ( n16 ) & ( n5196 )  ;
assign n5273 =  ( n16 ) & ( n5198 )  ;
assign n5274 =  ( n16 ) & ( n5200 )  ;
assign n5275 =  ( n16 ) & ( n5202 )  ;
assign n5276 =  ( n16 ) & ( n5204 )  ;
assign n5277 =  ( n16 ) & ( n5206 )  ;
assign n5278 =  ( n16 ) & ( n5208 )  ;
assign n5279 =  ( n16 ) & ( n5210 )  ;
assign n5280 =  ( n16 ) & ( n5212 )  ;
assign n5281 =  ( n16 ) & ( n5214 )  ;
assign n5282 =  ( n16 ) & ( n5216 )  ;
assign n5283 =  ( n16 ) & ( n5218 )  ;
assign n5284 =  ( n17 ) & ( n5188 )  ;
assign n5285 =  ( n17 ) & ( n5190 )  ;
assign n5286 =  ( n17 ) & ( n5192 )  ;
assign n5287 =  ( n17 ) & ( n5194 )  ;
assign n5288 =  ( n17 ) & ( n5196 )  ;
assign n5289 =  ( n17 ) & ( n5198 )  ;
assign n5290 =  ( n17 ) & ( n5200 )  ;
assign n5291 =  ( n17 ) & ( n5202 )  ;
assign n5292 =  ( n17 ) & ( n5204 )  ;
assign n5293 =  ( n17 ) & ( n5206 )  ;
assign n5294 =  ( n17 ) & ( n5208 )  ;
assign n5295 =  ( n17 ) & ( n5210 )  ;
assign n5296 =  ( n17 ) & ( n5212 )  ;
assign n5297 =  ( n17 ) & ( n5214 )  ;
assign n5298 =  ( n17 ) & ( n5216 )  ;
assign n5299 =  ( n17 ) & ( n5218 )  ;
assign n5300 =  ( n18 ) & ( n5188 )  ;
assign n5301 =  ( n18 ) & ( n5190 )  ;
assign n5302 =  ( n18 ) & ( n5192 )  ;
assign n5303 =  ( n18 ) & ( n5194 )  ;
assign n5304 =  ( n18 ) & ( n5196 )  ;
assign n5305 =  ( n18 ) & ( n5198 )  ;
assign n5306 =  ( n18 ) & ( n5200 )  ;
assign n5307 =  ( n18 ) & ( n5202 )  ;
assign n5308 =  ( n18 ) & ( n5204 )  ;
assign n5309 =  ( n18 ) & ( n5206 )  ;
assign n5310 =  ( n18 ) & ( n5208 )  ;
assign n5311 =  ( n18 ) & ( n5210 )  ;
assign n5312 =  ( n18 ) & ( n5212 )  ;
assign n5313 =  ( n18 ) & ( n5214 )  ;
assign n5314 =  ( n18 ) & ( n5216 )  ;
assign n5315 =  ( n18 ) & ( n5218 )  ;
assign n5316 =  ( n19 ) & ( n5188 )  ;
assign n5317 =  ( n19 ) & ( n5190 )  ;
assign n5318 =  ( n19 ) & ( n5192 )  ;
assign n5319 =  ( n19 ) & ( n5194 )  ;
assign n5320 =  ( n19 ) & ( n5196 )  ;
assign n5321 =  ( n19 ) & ( n5198 )  ;
assign n5322 =  ( n19 ) & ( n5200 )  ;
assign n5323 =  ( n19 ) & ( n5202 )  ;
assign n5324 =  ( n19 ) & ( n5204 )  ;
assign n5325 =  ( n19 ) & ( n5206 )  ;
assign n5326 =  ( n19 ) & ( n5208 )  ;
assign n5327 =  ( n19 ) & ( n5210 )  ;
assign n5328 =  ( n19 ) & ( n5212 )  ;
assign n5329 =  ( n19 ) & ( n5214 )  ;
assign n5330 =  ( n19 ) & ( n5216 )  ;
assign n5331 =  ( n19 ) & ( n5218 )  ;
assign n5332 =  ( n20 ) & ( n5188 )  ;
assign n5333 =  ( n20 ) & ( n5190 )  ;
assign n5334 =  ( n20 ) & ( n5192 )  ;
assign n5335 =  ( n20 ) & ( n5194 )  ;
assign n5336 =  ( n20 ) & ( n5196 )  ;
assign n5337 =  ( n20 ) & ( n5198 )  ;
assign n5338 =  ( n20 ) & ( n5200 )  ;
assign n5339 =  ( n20 ) & ( n5202 )  ;
assign n5340 =  ( n20 ) & ( n5204 )  ;
assign n5341 =  ( n20 ) & ( n5206 )  ;
assign n5342 =  ( n20 ) & ( n5208 )  ;
assign n5343 =  ( n20 ) & ( n5210 )  ;
assign n5344 =  ( n20 ) & ( n5212 )  ;
assign n5345 =  ( n20 ) & ( n5214 )  ;
assign n5346 =  ( n20 ) & ( n5216 )  ;
assign n5347 =  ( n20 ) & ( n5218 )  ;
assign n5348 =  ( n21 ) & ( n5188 )  ;
assign n5349 =  ( n21 ) & ( n5190 )  ;
assign n5350 =  ( n21 ) & ( n5192 )  ;
assign n5351 =  ( n21 ) & ( n5194 )  ;
assign n5352 =  ( n21 ) & ( n5196 )  ;
assign n5353 =  ( n21 ) & ( n5198 )  ;
assign n5354 =  ( n21 ) & ( n5200 )  ;
assign n5355 =  ( n21 ) & ( n5202 )  ;
assign n5356 =  ( n21 ) & ( n5204 )  ;
assign n5357 =  ( n21 ) & ( n5206 )  ;
assign n5358 =  ( n21 ) & ( n5208 )  ;
assign n5359 =  ( n21 ) & ( n5210 )  ;
assign n5360 =  ( n21 ) & ( n5212 )  ;
assign n5361 =  ( n21 ) & ( n5214 )  ;
assign n5362 =  ( n21 ) & ( n5216 )  ;
assign n5363 =  ( n21 ) & ( n5218 )  ;
assign n5364 =  ( n22 ) & ( n5188 )  ;
assign n5365 =  ( n22 ) & ( n5190 )  ;
assign n5366 =  ( n22 ) & ( n5192 )  ;
assign n5367 =  ( n22 ) & ( n5194 )  ;
assign n5368 =  ( n22 ) & ( n5196 )  ;
assign n5369 =  ( n22 ) & ( n5198 )  ;
assign n5370 =  ( n22 ) & ( n5200 )  ;
assign n5371 =  ( n22 ) & ( n5202 )  ;
assign n5372 =  ( n22 ) & ( n5204 )  ;
assign n5373 =  ( n22 ) & ( n5206 )  ;
assign n5374 =  ( n22 ) & ( n5208 )  ;
assign n5375 =  ( n22 ) & ( n5210 )  ;
assign n5376 =  ( n22 ) & ( n5212 )  ;
assign n5377 =  ( n22 ) & ( n5214 )  ;
assign n5378 =  ( n22 ) & ( n5216 )  ;
assign n5379 =  ( n22 ) & ( n5218 )  ;
assign n5380 =  ( n23 ) & ( n5188 )  ;
assign n5381 =  ( n23 ) & ( n5190 )  ;
assign n5382 =  ( n23 ) & ( n5192 )  ;
assign n5383 =  ( n23 ) & ( n5194 )  ;
assign n5384 =  ( n23 ) & ( n5196 )  ;
assign n5385 =  ( n23 ) & ( n5198 )  ;
assign n5386 =  ( n23 ) & ( n5200 )  ;
assign n5387 =  ( n23 ) & ( n5202 )  ;
assign n5388 =  ( n23 ) & ( n5204 )  ;
assign n5389 =  ( n23 ) & ( n5206 )  ;
assign n5390 =  ( n23 ) & ( n5208 )  ;
assign n5391 =  ( n23 ) & ( n5210 )  ;
assign n5392 =  ( n23 ) & ( n5212 )  ;
assign n5393 =  ( n23 ) & ( n5214 )  ;
assign n5394 =  ( n23 ) & ( n5216 )  ;
assign n5395 =  ( n23 ) & ( n5218 )  ;
assign n5396 =  ( n24 ) & ( n5188 )  ;
assign n5397 =  ( n24 ) & ( n5190 )  ;
assign n5398 =  ( n24 ) & ( n5192 )  ;
assign n5399 =  ( n24 ) & ( n5194 )  ;
assign n5400 =  ( n24 ) & ( n5196 )  ;
assign n5401 =  ( n24 ) & ( n5198 )  ;
assign n5402 =  ( n24 ) & ( n5200 )  ;
assign n5403 =  ( n24 ) & ( n5202 )  ;
assign n5404 =  ( n24 ) & ( n5204 )  ;
assign n5405 =  ( n24 ) & ( n5206 )  ;
assign n5406 =  ( n24 ) & ( n5208 )  ;
assign n5407 =  ( n24 ) & ( n5210 )  ;
assign n5408 =  ( n24 ) & ( n5212 )  ;
assign n5409 =  ( n24 ) & ( n5214 )  ;
assign n5410 =  ( n24 ) & ( n5216 )  ;
assign n5411 =  ( n24 ) & ( n5218 )  ;
assign n5412 =  ( n25 ) & ( n5188 )  ;
assign n5413 =  ( n25 ) & ( n5190 )  ;
assign n5414 =  ( n25 ) & ( n5192 )  ;
assign n5415 =  ( n25 ) & ( n5194 )  ;
assign n5416 =  ( n25 ) & ( n5196 )  ;
assign n5417 =  ( n25 ) & ( n5198 )  ;
assign n5418 =  ( n25 ) & ( n5200 )  ;
assign n5419 =  ( n25 ) & ( n5202 )  ;
assign n5420 =  ( n25 ) & ( n5204 )  ;
assign n5421 =  ( n25 ) & ( n5206 )  ;
assign n5422 =  ( n25 ) & ( n5208 )  ;
assign n5423 =  ( n25 ) & ( n5210 )  ;
assign n5424 =  ( n25 ) & ( n5212 )  ;
assign n5425 =  ( n25 ) & ( n5214 )  ;
assign n5426 =  ( n25 ) & ( n5216 )  ;
assign n5427 =  ( n25 ) & ( n5218 )  ;
assign n5428 =  ( n26 ) & ( n5188 )  ;
assign n5429 =  ( n26 ) & ( n5190 )  ;
assign n5430 =  ( n26 ) & ( n5192 )  ;
assign n5431 =  ( n26 ) & ( n5194 )  ;
assign n5432 =  ( n26 ) & ( n5196 )  ;
assign n5433 =  ( n26 ) & ( n5198 )  ;
assign n5434 =  ( n26 ) & ( n5200 )  ;
assign n5435 =  ( n26 ) & ( n5202 )  ;
assign n5436 =  ( n26 ) & ( n5204 )  ;
assign n5437 =  ( n26 ) & ( n5206 )  ;
assign n5438 =  ( n26 ) & ( n5208 )  ;
assign n5439 =  ( n26 ) & ( n5210 )  ;
assign n5440 =  ( n26 ) & ( n5212 )  ;
assign n5441 =  ( n26 ) & ( n5214 )  ;
assign n5442 =  ( n26 ) & ( n5216 )  ;
assign n5443 =  ( n26 ) & ( n5218 )  ;
assign n5444 =  ( n27 ) & ( n5188 )  ;
assign n5445 =  ( n27 ) & ( n5190 )  ;
assign n5446 =  ( n27 ) & ( n5192 )  ;
assign n5447 =  ( n27 ) & ( n5194 )  ;
assign n5448 =  ( n27 ) & ( n5196 )  ;
assign n5449 =  ( n27 ) & ( n5198 )  ;
assign n5450 =  ( n27 ) & ( n5200 )  ;
assign n5451 =  ( n27 ) & ( n5202 )  ;
assign n5452 =  ( n27 ) & ( n5204 )  ;
assign n5453 =  ( n27 ) & ( n5206 )  ;
assign n5454 =  ( n27 ) & ( n5208 )  ;
assign n5455 =  ( n27 ) & ( n5210 )  ;
assign n5456 =  ( n27 ) & ( n5212 )  ;
assign n5457 =  ( n27 ) & ( n5214 )  ;
assign n5458 =  ( n27 ) & ( n5216 )  ;
assign n5459 =  ( n27 ) & ( n5218 )  ;
assign n5460 =  ( n28 ) & ( n5188 )  ;
assign n5461 =  ( n28 ) & ( n5190 )  ;
assign n5462 =  ( n28 ) & ( n5192 )  ;
assign n5463 =  ( n28 ) & ( n5194 )  ;
assign n5464 =  ( n28 ) & ( n5196 )  ;
assign n5465 =  ( n28 ) & ( n5198 )  ;
assign n5466 =  ( n28 ) & ( n5200 )  ;
assign n5467 =  ( n28 ) & ( n5202 )  ;
assign n5468 =  ( n28 ) & ( n5204 )  ;
assign n5469 =  ( n28 ) & ( n5206 )  ;
assign n5470 =  ( n28 ) & ( n5208 )  ;
assign n5471 =  ( n28 ) & ( n5210 )  ;
assign n5472 =  ( n28 ) & ( n5212 )  ;
assign n5473 =  ( n28 ) & ( n5214 )  ;
assign n5474 =  ( n28 ) & ( n5216 )  ;
assign n5475 =  ( n28 ) & ( n5218 )  ;
assign n5476 =  ( n29 ) & ( n5188 )  ;
assign n5477 =  ( n29 ) & ( n5190 )  ;
assign n5478 =  ( n29 ) & ( n5192 )  ;
assign n5479 =  ( n29 ) & ( n5194 )  ;
assign n5480 =  ( n29 ) & ( n5196 )  ;
assign n5481 =  ( n29 ) & ( n5198 )  ;
assign n5482 =  ( n29 ) & ( n5200 )  ;
assign n5483 =  ( n29 ) & ( n5202 )  ;
assign n5484 =  ( n29 ) & ( n5204 )  ;
assign n5485 =  ( n29 ) & ( n5206 )  ;
assign n5486 =  ( n29 ) & ( n5208 )  ;
assign n5487 =  ( n29 ) & ( n5210 )  ;
assign n5488 =  ( n29 ) & ( n5212 )  ;
assign n5489 =  ( n29 ) & ( n5214 )  ;
assign n5490 =  ( n29 ) & ( n5216 )  ;
assign n5491 =  ( n29 ) & ( n5218 )  ;
assign n5492 =  ( n30 ) & ( n5188 )  ;
assign n5493 =  ( n30 ) & ( n5190 )  ;
assign n5494 =  ( n30 ) & ( n5192 )  ;
assign n5495 =  ( n30 ) & ( n5194 )  ;
assign n5496 =  ( n30 ) & ( n5196 )  ;
assign n5497 =  ( n30 ) & ( n5198 )  ;
assign n5498 =  ( n30 ) & ( n5200 )  ;
assign n5499 =  ( n30 ) & ( n5202 )  ;
assign n5500 =  ( n30 ) & ( n5204 )  ;
assign n5501 =  ( n30 ) & ( n5206 )  ;
assign n5502 =  ( n30 ) & ( n5208 )  ;
assign n5503 =  ( n30 ) & ( n5210 )  ;
assign n5504 =  ( n30 ) & ( n5212 )  ;
assign n5505 =  ( n30 ) & ( n5214 )  ;
assign n5506 =  ( n30 ) & ( n5216 )  ;
assign n5507 =  ( n30 ) & ( n5218 )  ;
assign n5508 =  ( n31 ) & ( n5188 )  ;
assign n5509 =  ( n31 ) & ( n5190 )  ;
assign n5510 =  ( n31 ) & ( n5192 )  ;
assign n5511 =  ( n31 ) & ( n5194 )  ;
assign n5512 =  ( n31 ) & ( n5196 )  ;
assign n5513 =  ( n31 ) & ( n5198 )  ;
assign n5514 =  ( n31 ) & ( n5200 )  ;
assign n5515 =  ( n31 ) & ( n5202 )  ;
assign n5516 =  ( n31 ) & ( n5204 )  ;
assign n5517 =  ( n31 ) & ( n5206 )  ;
assign n5518 =  ( n31 ) & ( n5208 )  ;
assign n5519 =  ( n31 ) & ( n5210 )  ;
assign n5520 =  ( n31 ) & ( n5212 )  ;
assign n5521 =  ( n31 ) & ( n5214 )  ;
assign n5522 =  ( n31 ) & ( n5216 )  ;
assign n5523 =  ( n31 ) & ( n5218 )  ;
assign n5524 =  ( n32 ) & ( n5188 )  ;
assign n5525 =  ( n32 ) & ( n5190 )  ;
assign n5526 =  ( n32 ) & ( n5192 )  ;
assign n5527 =  ( n32 ) & ( n5194 )  ;
assign n5528 =  ( n32 ) & ( n5196 )  ;
assign n5529 =  ( n32 ) & ( n5198 )  ;
assign n5530 =  ( n32 ) & ( n5200 )  ;
assign n5531 =  ( n32 ) & ( n5202 )  ;
assign n5532 =  ( n32 ) & ( n5204 )  ;
assign n5533 =  ( n32 ) & ( n5206 )  ;
assign n5534 =  ( n32 ) & ( n5208 )  ;
assign n5535 =  ( n32 ) & ( n5210 )  ;
assign n5536 =  ( n32 ) & ( n5212 )  ;
assign n5537 =  ( n32 ) & ( n5214 )  ;
assign n5538 =  ( n32 ) & ( n5216 )  ;
assign n5539 =  ( n32 ) & ( n5218 )  ;
assign n5540 =  ( n33 ) & ( n5188 )  ;
assign n5541 =  ( n33 ) & ( n5190 )  ;
assign n5542 =  ( n33 ) & ( n5192 )  ;
assign n5543 =  ( n33 ) & ( n5194 )  ;
assign n5544 =  ( n33 ) & ( n5196 )  ;
assign n5545 =  ( n33 ) & ( n5198 )  ;
assign n5546 =  ( n33 ) & ( n5200 )  ;
assign n5547 =  ( n33 ) & ( n5202 )  ;
assign n5548 =  ( n33 ) & ( n5204 )  ;
assign n5549 =  ( n33 ) & ( n5206 )  ;
assign n5550 =  ( n33 ) & ( n5208 )  ;
assign n5551 =  ( n33 ) & ( n5210 )  ;
assign n5552 =  ( n33 ) & ( n5212 )  ;
assign n5553 =  ( n33 ) & ( n5214 )  ;
assign n5554 =  ( n33 ) & ( n5216 )  ;
assign n5555 =  ( n33 ) & ( n5218 )  ;
assign n5556 =  ( n34 ) & ( n5188 )  ;
assign n5557 =  ( n34 ) & ( n5190 )  ;
assign n5558 =  ( n34 ) & ( n5192 )  ;
assign n5559 =  ( n34 ) & ( n5194 )  ;
assign n5560 =  ( n34 ) & ( n5196 )  ;
assign n5561 =  ( n34 ) & ( n5198 )  ;
assign n5562 =  ( n34 ) & ( n5200 )  ;
assign n5563 =  ( n34 ) & ( n5202 )  ;
assign n5564 =  ( n34 ) & ( n5204 )  ;
assign n5565 =  ( n34 ) & ( n5206 )  ;
assign n5566 =  ( n34 ) & ( n5208 )  ;
assign n5567 =  ( n34 ) & ( n5210 )  ;
assign n5568 =  ( n34 ) & ( n5212 )  ;
assign n5569 =  ( n34 ) & ( n5214 )  ;
assign n5570 =  ( n34 ) & ( n5216 )  ;
assign n5571 =  ( n34 ) & ( n5218 )  ;
assign n5572 =  ( n35 ) & ( n5188 )  ;
assign n5573 =  ( n35 ) & ( n5190 )  ;
assign n5574 =  ( n35 ) & ( n5192 )  ;
assign n5575 =  ( n35 ) & ( n5194 )  ;
assign n5576 =  ( n35 ) & ( n5196 )  ;
assign n5577 =  ( n35 ) & ( n5198 )  ;
assign n5578 =  ( n35 ) & ( n5200 )  ;
assign n5579 =  ( n35 ) & ( n5202 )  ;
assign n5580 =  ( n35 ) & ( n5204 )  ;
assign n5581 =  ( n35 ) & ( n5206 )  ;
assign n5582 =  ( n35 ) & ( n5208 )  ;
assign n5583 =  ( n35 ) & ( n5210 )  ;
assign n5584 =  ( n35 ) & ( n5212 )  ;
assign n5585 =  ( n35 ) & ( n5214 )  ;
assign n5586 =  ( n35 ) & ( n5216 )  ;
assign n5587 =  ( n35 ) & ( n5218 )  ;
assign n5588 =  ( n36 ) & ( n5188 )  ;
assign n5589 =  ( n36 ) & ( n5190 )  ;
assign n5590 =  ( n36 ) & ( n5192 )  ;
assign n5591 =  ( n36 ) & ( n5194 )  ;
assign n5592 =  ( n36 ) & ( n5196 )  ;
assign n5593 =  ( n36 ) & ( n5198 )  ;
assign n5594 =  ( n36 ) & ( n5200 )  ;
assign n5595 =  ( n36 ) & ( n5202 )  ;
assign n5596 =  ( n36 ) & ( n5204 )  ;
assign n5597 =  ( n36 ) & ( n5206 )  ;
assign n5598 =  ( n36 ) & ( n5208 )  ;
assign n5599 =  ( n36 ) & ( n5210 )  ;
assign n5600 =  ( n36 ) & ( n5212 )  ;
assign n5601 =  ( n36 ) & ( n5214 )  ;
assign n5602 =  ( n36 ) & ( n5216 )  ;
assign n5603 =  ( n36 ) & ( n5218 )  ;
assign n5604 =  ( n37 ) & ( n5188 )  ;
assign n5605 =  ( n37 ) & ( n5190 )  ;
assign n5606 =  ( n37 ) & ( n5192 )  ;
assign n5607 =  ( n37 ) & ( n5194 )  ;
assign n5608 =  ( n37 ) & ( n5196 )  ;
assign n5609 =  ( n37 ) & ( n5198 )  ;
assign n5610 =  ( n37 ) & ( n5200 )  ;
assign n5611 =  ( n37 ) & ( n5202 )  ;
assign n5612 =  ( n37 ) & ( n5204 )  ;
assign n5613 =  ( n37 ) & ( n5206 )  ;
assign n5614 =  ( n37 ) & ( n5208 )  ;
assign n5615 =  ( n37 ) & ( n5210 )  ;
assign n5616 =  ( n37 ) & ( n5212 )  ;
assign n5617 =  ( n37 ) & ( n5214 )  ;
assign n5618 =  ( n37 ) & ( n5216 )  ;
assign n5619 =  ( n37 ) & ( n5218 )  ;
assign n5620 =  ( n38 ) & ( n5188 )  ;
assign n5621 =  ( n38 ) & ( n5190 )  ;
assign n5622 =  ( n38 ) & ( n5192 )  ;
assign n5623 =  ( n38 ) & ( n5194 )  ;
assign n5624 =  ( n38 ) & ( n5196 )  ;
assign n5625 =  ( n38 ) & ( n5198 )  ;
assign n5626 =  ( n38 ) & ( n5200 )  ;
assign n5627 =  ( n38 ) & ( n5202 )  ;
assign n5628 =  ( n38 ) & ( n5204 )  ;
assign n5629 =  ( n38 ) & ( n5206 )  ;
assign n5630 =  ( n38 ) & ( n5208 )  ;
assign n5631 =  ( n38 ) & ( n5210 )  ;
assign n5632 =  ( n38 ) & ( n5212 )  ;
assign n5633 =  ( n38 ) & ( n5214 )  ;
assign n5634 =  ( n38 ) & ( n5216 )  ;
assign n5635 =  ( n38 ) & ( n5218 )  ;
assign n5636 =  ( n39 ) & ( n5188 )  ;
assign n5637 =  ( n39 ) & ( n5190 )  ;
assign n5638 =  ( n39 ) & ( n5192 )  ;
assign n5639 =  ( n39 ) & ( n5194 )  ;
assign n5640 =  ( n39 ) & ( n5196 )  ;
assign n5641 =  ( n39 ) & ( n5198 )  ;
assign n5642 =  ( n39 ) & ( n5200 )  ;
assign n5643 =  ( n39 ) & ( n5202 )  ;
assign n5644 =  ( n39 ) & ( n5204 )  ;
assign n5645 =  ( n39 ) & ( n5206 )  ;
assign n5646 =  ( n39 ) & ( n5208 )  ;
assign n5647 =  ( n39 ) & ( n5210 )  ;
assign n5648 =  ( n39 ) & ( n5212 )  ;
assign n5649 =  ( n39 ) & ( n5214 )  ;
assign n5650 =  ( n39 ) & ( n5216 )  ;
assign n5651 =  ( n39 ) & ( n5218 )  ;
assign n5652 =  ( n40 ) & ( n5188 )  ;
assign n5653 =  ( n40 ) & ( n5190 )  ;
assign n5654 =  ( n40 ) & ( n5192 )  ;
assign n5655 =  ( n40 ) & ( n5194 )  ;
assign n5656 =  ( n40 ) & ( n5196 )  ;
assign n5657 =  ( n40 ) & ( n5198 )  ;
assign n5658 =  ( n40 ) & ( n5200 )  ;
assign n5659 =  ( n40 ) & ( n5202 )  ;
assign n5660 =  ( n40 ) & ( n5204 )  ;
assign n5661 =  ( n40 ) & ( n5206 )  ;
assign n5662 =  ( n40 ) & ( n5208 )  ;
assign n5663 =  ( n40 ) & ( n5210 )  ;
assign n5664 =  ( n40 ) & ( n5212 )  ;
assign n5665 =  ( n40 ) & ( n5214 )  ;
assign n5666 =  ( n40 ) & ( n5216 )  ;
assign n5667 =  ( n40 ) & ( n5218 )  ;
assign n5668 =  ( n41 ) & ( n5188 )  ;
assign n5669 =  ( n41 ) & ( n5190 )  ;
assign n5670 =  ( n41 ) & ( n5192 )  ;
assign n5671 =  ( n41 ) & ( n5194 )  ;
assign n5672 =  ( n41 ) & ( n5196 )  ;
assign n5673 =  ( n41 ) & ( n5198 )  ;
assign n5674 =  ( n41 ) & ( n5200 )  ;
assign n5675 =  ( n41 ) & ( n5202 )  ;
assign n5676 =  ( n41 ) & ( n5204 )  ;
assign n5677 =  ( n41 ) & ( n5206 )  ;
assign n5678 =  ( n41 ) & ( n5208 )  ;
assign n5679 =  ( n41 ) & ( n5210 )  ;
assign n5680 =  ( n41 ) & ( n5212 )  ;
assign n5681 =  ( n41 ) & ( n5214 )  ;
assign n5682 =  ( n41 ) & ( n5216 )  ;
assign n5683 =  ( n41 ) & ( n5218 )  ;
assign n5684 =  ( n42 ) & ( n5188 )  ;
assign n5685 =  ( n42 ) & ( n5190 )  ;
assign n5686 =  ( n42 ) & ( n5192 )  ;
assign n5687 =  ( n42 ) & ( n5194 )  ;
assign n5688 =  ( n42 ) & ( n5196 )  ;
assign n5689 =  ( n42 ) & ( n5198 )  ;
assign n5690 =  ( n42 ) & ( n5200 )  ;
assign n5691 =  ( n42 ) & ( n5202 )  ;
assign n5692 =  ( n42 ) & ( n5204 )  ;
assign n5693 =  ( n42 ) & ( n5206 )  ;
assign n5694 =  ( n42 ) & ( n5208 )  ;
assign n5695 =  ( n42 ) & ( n5210 )  ;
assign n5696 =  ( n42 ) & ( n5212 )  ;
assign n5697 =  ( n42 ) & ( n5214 )  ;
assign n5698 =  ( n42 ) & ( n5216 )  ;
assign n5699 =  ( n42 ) & ( n5218 )  ;
assign n5700 =  ( n43 ) & ( n5188 )  ;
assign n5701 =  ( n43 ) & ( n5190 )  ;
assign n5702 =  ( n43 ) & ( n5192 )  ;
assign n5703 =  ( n43 ) & ( n5194 )  ;
assign n5704 =  ( n43 ) & ( n5196 )  ;
assign n5705 =  ( n43 ) & ( n5198 )  ;
assign n5706 =  ( n43 ) & ( n5200 )  ;
assign n5707 =  ( n43 ) & ( n5202 )  ;
assign n5708 =  ( n43 ) & ( n5204 )  ;
assign n5709 =  ( n43 ) & ( n5206 )  ;
assign n5710 =  ( n43 ) & ( n5208 )  ;
assign n5711 =  ( n43 ) & ( n5210 )  ;
assign n5712 =  ( n43 ) & ( n5212 )  ;
assign n5713 =  ( n43 ) & ( n5214 )  ;
assign n5714 =  ( n43 ) & ( n5216 )  ;
assign n5715 =  ( n43 ) & ( n5218 )  ;
assign n5716 =  ( n5715 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n5717 =  ( n5714 ) ? ( VREG_0_1 ) : ( n5716 ) ;
assign n5718 =  ( n5713 ) ? ( VREG_0_2 ) : ( n5717 ) ;
assign n5719 =  ( n5712 ) ? ( VREG_0_3 ) : ( n5718 ) ;
assign n5720 =  ( n5711 ) ? ( VREG_0_4 ) : ( n5719 ) ;
assign n5721 =  ( n5710 ) ? ( VREG_0_5 ) : ( n5720 ) ;
assign n5722 =  ( n5709 ) ? ( VREG_0_6 ) : ( n5721 ) ;
assign n5723 =  ( n5708 ) ? ( VREG_0_7 ) : ( n5722 ) ;
assign n5724 =  ( n5707 ) ? ( VREG_0_8 ) : ( n5723 ) ;
assign n5725 =  ( n5706 ) ? ( VREG_0_9 ) : ( n5724 ) ;
assign n5726 =  ( n5705 ) ? ( VREG_0_10 ) : ( n5725 ) ;
assign n5727 =  ( n5704 ) ? ( VREG_0_11 ) : ( n5726 ) ;
assign n5728 =  ( n5703 ) ? ( VREG_0_12 ) : ( n5727 ) ;
assign n5729 =  ( n5702 ) ? ( VREG_0_13 ) : ( n5728 ) ;
assign n5730 =  ( n5701 ) ? ( VREG_0_14 ) : ( n5729 ) ;
assign n5731 =  ( n5700 ) ? ( VREG_0_15 ) : ( n5730 ) ;
assign n5732 =  ( n5699 ) ? ( VREG_1_0 ) : ( n5731 ) ;
assign n5733 =  ( n5698 ) ? ( VREG_1_1 ) : ( n5732 ) ;
assign n5734 =  ( n5697 ) ? ( VREG_1_2 ) : ( n5733 ) ;
assign n5735 =  ( n5696 ) ? ( VREG_1_3 ) : ( n5734 ) ;
assign n5736 =  ( n5695 ) ? ( VREG_1_4 ) : ( n5735 ) ;
assign n5737 =  ( n5694 ) ? ( VREG_1_5 ) : ( n5736 ) ;
assign n5738 =  ( n5693 ) ? ( VREG_1_6 ) : ( n5737 ) ;
assign n5739 =  ( n5692 ) ? ( VREG_1_7 ) : ( n5738 ) ;
assign n5740 =  ( n5691 ) ? ( VREG_1_8 ) : ( n5739 ) ;
assign n5741 =  ( n5690 ) ? ( VREG_1_9 ) : ( n5740 ) ;
assign n5742 =  ( n5689 ) ? ( VREG_1_10 ) : ( n5741 ) ;
assign n5743 =  ( n5688 ) ? ( VREG_1_11 ) : ( n5742 ) ;
assign n5744 =  ( n5687 ) ? ( VREG_1_12 ) : ( n5743 ) ;
assign n5745 =  ( n5686 ) ? ( VREG_1_13 ) : ( n5744 ) ;
assign n5746 =  ( n5685 ) ? ( VREG_1_14 ) : ( n5745 ) ;
assign n5747 =  ( n5684 ) ? ( VREG_1_15 ) : ( n5746 ) ;
assign n5748 =  ( n5683 ) ? ( VREG_2_0 ) : ( n5747 ) ;
assign n5749 =  ( n5682 ) ? ( VREG_2_1 ) : ( n5748 ) ;
assign n5750 =  ( n5681 ) ? ( VREG_2_2 ) : ( n5749 ) ;
assign n5751 =  ( n5680 ) ? ( VREG_2_3 ) : ( n5750 ) ;
assign n5752 =  ( n5679 ) ? ( VREG_2_4 ) : ( n5751 ) ;
assign n5753 =  ( n5678 ) ? ( VREG_2_5 ) : ( n5752 ) ;
assign n5754 =  ( n5677 ) ? ( VREG_2_6 ) : ( n5753 ) ;
assign n5755 =  ( n5676 ) ? ( VREG_2_7 ) : ( n5754 ) ;
assign n5756 =  ( n5675 ) ? ( VREG_2_8 ) : ( n5755 ) ;
assign n5757 =  ( n5674 ) ? ( VREG_2_9 ) : ( n5756 ) ;
assign n5758 =  ( n5673 ) ? ( VREG_2_10 ) : ( n5757 ) ;
assign n5759 =  ( n5672 ) ? ( VREG_2_11 ) : ( n5758 ) ;
assign n5760 =  ( n5671 ) ? ( VREG_2_12 ) : ( n5759 ) ;
assign n5761 =  ( n5670 ) ? ( VREG_2_13 ) : ( n5760 ) ;
assign n5762 =  ( n5669 ) ? ( VREG_2_14 ) : ( n5761 ) ;
assign n5763 =  ( n5668 ) ? ( VREG_2_15 ) : ( n5762 ) ;
assign n5764 =  ( n5667 ) ? ( VREG_3_0 ) : ( n5763 ) ;
assign n5765 =  ( n5666 ) ? ( VREG_3_1 ) : ( n5764 ) ;
assign n5766 =  ( n5665 ) ? ( VREG_3_2 ) : ( n5765 ) ;
assign n5767 =  ( n5664 ) ? ( VREG_3_3 ) : ( n5766 ) ;
assign n5768 =  ( n5663 ) ? ( VREG_3_4 ) : ( n5767 ) ;
assign n5769 =  ( n5662 ) ? ( VREG_3_5 ) : ( n5768 ) ;
assign n5770 =  ( n5661 ) ? ( VREG_3_6 ) : ( n5769 ) ;
assign n5771 =  ( n5660 ) ? ( VREG_3_7 ) : ( n5770 ) ;
assign n5772 =  ( n5659 ) ? ( VREG_3_8 ) : ( n5771 ) ;
assign n5773 =  ( n5658 ) ? ( VREG_3_9 ) : ( n5772 ) ;
assign n5774 =  ( n5657 ) ? ( VREG_3_10 ) : ( n5773 ) ;
assign n5775 =  ( n5656 ) ? ( VREG_3_11 ) : ( n5774 ) ;
assign n5776 =  ( n5655 ) ? ( VREG_3_12 ) : ( n5775 ) ;
assign n5777 =  ( n5654 ) ? ( VREG_3_13 ) : ( n5776 ) ;
assign n5778 =  ( n5653 ) ? ( VREG_3_14 ) : ( n5777 ) ;
assign n5779 =  ( n5652 ) ? ( VREG_3_15 ) : ( n5778 ) ;
assign n5780 =  ( n5651 ) ? ( VREG_4_0 ) : ( n5779 ) ;
assign n5781 =  ( n5650 ) ? ( VREG_4_1 ) : ( n5780 ) ;
assign n5782 =  ( n5649 ) ? ( VREG_4_2 ) : ( n5781 ) ;
assign n5783 =  ( n5648 ) ? ( VREG_4_3 ) : ( n5782 ) ;
assign n5784 =  ( n5647 ) ? ( VREG_4_4 ) : ( n5783 ) ;
assign n5785 =  ( n5646 ) ? ( VREG_4_5 ) : ( n5784 ) ;
assign n5786 =  ( n5645 ) ? ( VREG_4_6 ) : ( n5785 ) ;
assign n5787 =  ( n5644 ) ? ( VREG_4_7 ) : ( n5786 ) ;
assign n5788 =  ( n5643 ) ? ( VREG_4_8 ) : ( n5787 ) ;
assign n5789 =  ( n5642 ) ? ( VREG_4_9 ) : ( n5788 ) ;
assign n5790 =  ( n5641 ) ? ( VREG_4_10 ) : ( n5789 ) ;
assign n5791 =  ( n5640 ) ? ( VREG_4_11 ) : ( n5790 ) ;
assign n5792 =  ( n5639 ) ? ( VREG_4_12 ) : ( n5791 ) ;
assign n5793 =  ( n5638 ) ? ( VREG_4_13 ) : ( n5792 ) ;
assign n5794 =  ( n5637 ) ? ( VREG_4_14 ) : ( n5793 ) ;
assign n5795 =  ( n5636 ) ? ( VREG_4_15 ) : ( n5794 ) ;
assign n5796 =  ( n5635 ) ? ( VREG_5_0 ) : ( n5795 ) ;
assign n5797 =  ( n5634 ) ? ( VREG_5_1 ) : ( n5796 ) ;
assign n5798 =  ( n5633 ) ? ( VREG_5_2 ) : ( n5797 ) ;
assign n5799 =  ( n5632 ) ? ( VREG_5_3 ) : ( n5798 ) ;
assign n5800 =  ( n5631 ) ? ( VREG_5_4 ) : ( n5799 ) ;
assign n5801 =  ( n5630 ) ? ( VREG_5_5 ) : ( n5800 ) ;
assign n5802 =  ( n5629 ) ? ( VREG_5_6 ) : ( n5801 ) ;
assign n5803 =  ( n5628 ) ? ( VREG_5_7 ) : ( n5802 ) ;
assign n5804 =  ( n5627 ) ? ( VREG_5_8 ) : ( n5803 ) ;
assign n5805 =  ( n5626 ) ? ( VREG_5_9 ) : ( n5804 ) ;
assign n5806 =  ( n5625 ) ? ( VREG_5_10 ) : ( n5805 ) ;
assign n5807 =  ( n5624 ) ? ( VREG_5_11 ) : ( n5806 ) ;
assign n5808 =  ( n5623 ) ? ( VREG_5_12 ) : ( n5807 ) ;
assign n5809 =  ( n5622 ) ? ( VREG_5_13 ) : ( n5808 ) ;
assign n5810 =  ( n5621 ) ? ( VREG_5_14 ) : ( n5809 ) ;
assign n5811 =  ( n5620 ) ? ( VREG_5_15 ) : ( n5810 ) ;
assign n5812 =  ( n5619 ) ? ( VREG_6_0 ) : ( n5811 ) ;
assign n5813 =  ( n5618 ) ? ( VREG_6_1 ) : ( n5812 ) ;
assign n5814 =  ( n5617 ) ? ( VREG_6_2 ) : ( n5813 ) ;
assign n5815 =  ( n5616 ) ? ( VREG_6_3 ) : ( n5814 ) ;
assign n5816 =  ( n5615 ) ? ( VREG_6_4 ) : ( n5815 ) ;
assign n5817 =  ( n5614 ) ? ( VREG_6_5 ) : ( n5816 ) ;
assign n5818 =  ( n5613 ) ? ( VREG_6_6 ) : ( n5817 ) ;
assign n5819 =  ( n5612 ) ? ( VREG_6_7 ) : ( n5818 ) ;
assign n5820 =  ( n5611 ) ? ( VREG_6_8 ) : ( n5819 ) ;
assign n5821 =  ( n5610 ) ? ( VREG_6_9 ) : ( n5820 ) ;
assign n5822 =  ( n5609 ) ? ( VREG_6_10 ) : ( n5821 ) ;
assign n5823 =  ( n5608 ) ? ( VREG_6_11 ) : ( n5822 ) ;
assign n5824 =  ( n5607 ) ? ( VREG_6_12 ) : ( n5823 ) ;
assign n5825 =  ( n5606 ) ? ( VREG_6_13 ) : ( n5824 ) ;
assign n5826 =  ( n5605 ) ? ( VREG_6_14 ) : ( n5825 ) ;
assign n5827 =  ( n5604 ) ? ( VREG_6_15 ) : ( n5826 ) ;
assign n5828 =  ( n5603 ) ? ( VREG_7_0 ) : ( n5827 ) ;
assign n5829 =  ( n5602 ) ? ( VREG_7_1 ) : ( n5828 ) ;
assign n5830 =  ( n5601 ) ? ( VREG_7_2 ) : ( n5829 ) ;
assign n5831 =  ( n5600 ) ? ( VREG_7_3 ) : ( n5830 ) ;
assign n5832 =  ( n5599 ) ? ( VREG_7_4 ) : ( n5831 ) ;
assign n5833 =  ( n5598 ) ? ( VREG_7_5 ) : ( n5832 ) ;
assign n5834 =  ( n5597 ) ? ( VREG_7_6 ) : ( n5833 ) ;
assign n5835 =  ( n5596 ) ? ( VREG_7_7 ) : ( n5834 ) ;
assign n5836 =  ( n5595 ) ? ( VREG_7_8 ) : ( n5835 ) ;
assign n5837 =  ( n5594 ) ? ( VREG_7_9 ) : ( n5836 ) ;
assign n5838 =  ( n5593 ) ? ( VREG_7_10 ) : ( n5837 ) ;
assign n5839 =  ( n5592 ) ? ( VREG_7_11 ) : ( n5838 ) ;
assign n5840 =  ( n5591 ) ? ( VREG_7_12 ) : ( n5839 ) ;
assign n5841 =  ( n5590 ) ? ( VREG_7_13 ) : ( n5840 ) ;
assign n5842 =  ( n5589 ) ? ( VREG_7_14 ) : ( n5841 ) ;
assign n5843 =  ( n5588 ) ? ( VREG_7_15 ) : ( n5842 ) ;
assign n5844 =  ( n5587 ) ? ( VREG_8_0 ) : ( n5843 ) ;
assign n5845 =  ( n5586 ) ? ( VREG_8_1 ) : ( n5844 ) ;
assign n5846 =  ( n5585 ) ? ( VREG_8_2 ) : ( n5845 ) ;
assign n5847 =  ( n5584 ) ? ( VREG_8_3 ) : ( n5846 ) ;
assign n5848 =  ( n5583 ) ? ( VREG_8_4 ) : ( n5847 ) ;
assign n5849 =  ( n5582 ) ? ( VREG_8_5 ) : ( n5848 ) ;
assign n5850 =  ( n5581 ) ? ( VREG_8_6 ) : ( n5849 ) ;
assign n5851 =  ( n5580 ) ? ( VREG_8_7 ) : ( n5850 ) ;
assign n5852 =  ( n5579 ) ? ( VREG_8_8 ) : ( n5851 ) ;
assign n5853 =  ( n5578 ) ? ( VREG_8_9 ) : ( n5852 ) ;
assign n5854 =  ( n5577 ) ? ( VREG_8_10 ) : ( n5853 ) ;
assign n5855 =  ( n5576 ) ? ( VREG_8_11 ) : ( n5854 ) ;
assign n5856 =  ( n5575 ) ? ( VREG_8_12 ) : ( n5855 ) ;
assign n5857 =  ( n5574 ) ? ( VREG_8_13 ) : ( n5856 ) ;
assign n5858 =  ( n5573 ) ? ( VREG_8_14 ) : ( n5857 ) ;
assign n5859 =  ( n5572 ) ? ( VREG_8_15 ) : ( n5858 ) ;
assign n5860 =  ( n5571 ) ? ( VREG_9_0 ) : ( n5859 ) ;
assign n5861 =  ( n5570 ) ? ( VREG_9_1 ) : ( n5860 ) ;
assign n5862 =  ( n5569 ) ? ( VREG_9_2 ) : ( n5861 ) ;
assign n5863 =  ( n5568 ) ? ( VREG_9_3 ) : ( n5862 ) ;
assign n5864 =  ( n5567 ) ? ( VREG_9_4 ) : ( n5863 ) ;
assign n5865 =  ( n5566 ) ? ( VREG_9_5 ) : ( n5864 ) ;
assign n5866 =  ( n5565 ) ? ( VREG_9_6 ) : ( n5865 ) ;
assign n5867 =  ( n5564 ) ? ( VREG_9_7 ) : ( n5866 ) ;
assign n5868 =  ( n5563 ) ? ( VREG_9_8 ) : ( n5867 ) ;
assign n5869 =  ( n5562 ) ? ( VREG_9_9 ) : ( n5868 ) ;
assign n5870 =  ( n5561 ) ? ( VREG_9_10 ) : ( n5869 ) ;
assign n5871 =  ( n5560 ) ? ( VREG_9_11 ) : ( n5870 ) ;
assign n5872 =  ( n5559 ) ? ( VREG_9_12 ) : ( n5871 ) ;
assign n5873 =  ( n5558 ) ? ( VREG_9_13 ) : ( n5872 ) ;
assign n5874 =  ( n5557 ) ? ( VREG_9_14 ) : ( n5873 ) ;
assign n5875 =  ( n5556 ) ? ( VREG_9_15 ) : ( n5874 ) ;
assign n5876 =  ( n5555 ) ? ( VREG_10_0 ) : ( n5875 ) ;
assign n5877 =  ( n5554 ) ? ( VREG_10_1 ) : ( n5876 ) ;
assign n5878 =  ( n5553 ) ? ( VREG_10_2 ) : ( n5877 ) ;
assign n5879 =  ( n5552 ) ? ( VREG_10_3 ) : ( n5878 ) ;
assign n5880 =  ( n5551 ) ? ( VREG_10_4 ) : ( n5879 ) ;
assign n5881 =  ( n5550 ) ? ( VREG_10_5 ) : ( n5880 ) ;
assign n5882 =  ( n5549 ) ? ( VREG_10_6 ) : ( n5881 ) ;
assign n5883 =  ( n5548 ) ? ( VREG_10_7 ) : ( n5882 ) ;
assign n5884 =  ( n5547 ) ? ( VREG_10_8 ) : ( n5883 ) ;
assign n5885 =  ( n5546 ) ? ( VREG_10_9 ) : ( n5884 ) ;
assign n5886 =  ( n5545 ) ? ( VREG_10_10 ) : ( n5885 ) ;
assign n5887 =  ( n5544 ) ? ( VREG_10_11 ) : ( n5886 ) ;
assign n5888 =  ( n5543 ) ? ( VREG_10_12 ) : ( n5887 ) ;
assign n5889 =  ( n5542 ) ? ( VREG_10_13 ) : ( n5888 ) ;
assign n5890 =  ( n5541 ) ? ( VREG_10_14 ) : ( n5889 ) ;
assign n5891 =  ( n5540 ) ? ( VREG_10_15 ) : ( n5890 ) ;
assign n5892 =  ( n5539 ) ? ( VREG_11_0 ) : ( n5891 ) ;
assign n5893 =  ( n5538 ) ? ( VREG_11_1 ) : ( n5892 ) ;
assign n5894 =  ( n5537 ) ? ( VREG_11_2 ) : ( n5893 ) ;
assign n5895 =  ( n5536 ) ? ( VREG_11_3 ) : ( n5894 ) ;
assign n5896 =  ( n5535 ) ? ( VREG_11_4 ) : ( n5895 ) ;
assign n5897 =  ( n5534 ) ? ( VREG_11_5 ) : ( n5896 ) ;
assign n5898 =  ( n5533 ) ? ( VREG_11_6 ) : ( n5897 ) ;
assign n5899 =  ( n5532 ) ? ( VREG_11_7 ) : ( n5898 ) ;
assign n5900 =  ( n5531 ) ? ( VREG_11_8 ) : ( n5899 ) ;
assign n5901 =  ( n5530 ) ? ( VREG_11_9 ) : ( n5900 ) ;
assign n5902 =  ( n5529 ) ? ( VREG_11_10 ) : ( n5901 ) ;
assign n5903 =  ( n5528 ) ? ( VREG_11_11 ) : ( n5902 ) ;
assign n5904 =  ( n5527 ) ? ( VREG_11_12 ) : ( n5903 ) ;
assign n5905 =  ( n5526 ) ? ( VREG_11_13 ) : ( n5904 ) ;
assign n5906 =  ( n5525 ) ? ( VREG_11_14 ) : ( n5905 ) ;
assign n5907 =  ( n5524 ) ? ( VREG_11_15 ) : ( n5906 ) ;
assign n5908 =  ( n5523 ) ? ( VREG_12_0 ) : ( n5907 ) ;
assign n5909 =  ( n5522 ) ? ( VREG_12_1 ) : ( n5908 ) ;
assign n5910 =  ( n5521 ) ? ( VREG_12_2 ) : ( n5909 ) ;
assign n5911 =  ( n5520 ) ? ( VREG_12_3 ) : ( n5910 ) ;
assign n5912 =  ( n5519 ) ? ( VREG_12_4 ) : ( n5911 ) ;
assign n5913 =  ( n5518 ) ? ( VREG_12_5 ) : ( n5912 ) ;
assign n5914 =  ( n5517 ) ? ( VREG_12_6 ) : ( n5913 ) ;
assign n5915 =  ( n5516 ) ? ( VREG_12_7 ) : ( n5914 ) ;
assign n5916 =  ( n5515 ) ? ( VREG_12_8 ) : ( n5915 ) ;
assign n5917 =  ( n5514 ) ? ( VREG_12_9 ) : ( n5916 ) ;
assign n5918 =  ( n5513 ) ? ( VREG_12_10 ) : ( n5917 ) ;
assign n5919 =  ( n5512 ) ? ( VREG_12_11 ) : ( n5918 ) ;
assign n5920 =  ( n5511 ) ? ( VREG_12_12 ) : ( n5919 ) ;
assign n5921 =  ( n5510 ) ? ( VREG_12_13 ) : ( n5920 ) ;
assign n5922 =  ( n5509 ) ? ( VREG_12_14 ) : ( n5921 ) ;
assign n5923 =  ( n5508 ) ? ( VREG_12_15 ) : ( n5922 ) ;
assign n5924 =  ( n5507 ) ? ( VREG_13_0 ) : ( n5923 ) ;
assign n5925 =  ( n5506 ) ? ( VREG_13_1 ) : ( n5924 ) ;
assign n5926 =  ( n5505 ) ? ( VREG_13_2 ) : ( n5925 ) ;
assign n5927 =  ( n5504 ) ? ( VREG_13_3 ) : ( n5926 ) ;
assign n5928 =  ( n5503 ) ? ( VREG_13_4 ) : ( n5927 ) ;
assign n5929 =  ( n5502 ) ? ( VREG_13_5 ) : ( n5928 ) ;
assign n5930 =  ( n5501 ) ? ( VREG_13_6 ) : ( n5929 ) ;
assign n5931 =  ( n5500 ) ? ( VREG_13_7 ) : ( n5930 ) ;
assign n5932 =  ( n5499 ) ? ( VREG_13_8 ) : ( n5931 ) ;
assign n5933 =  ( n5498 ) ? ( VREG_13_9 ) : ( n5932 ) ;
assign n5934 =  ( n5497 ) ? ( VREG_13_10 ) : ( n5933 ) ;
assign n5935 =  ( n5496 ) ? ( VREG_13_11 ) : ( n5934 ) ;
assign n5936 =  ( n5495 ) ? ( VREG_13_12 ) : ( n5935 ) ;
assign n5937 =  ( n5494 ) ? ( VREG_13_13 ) : ( n5936 ) ;
assign n5938 =  ( n5493 ) ? ( VREG_13_14 ) : ( n5937 ) ;
assign n5939 =  ( n5492 ) ? ( VREG_13_15 ) : ( n5938 ) ;
assign n5940 =  ( n5491 ) ? ( VREG_14_0 ) : ( n5939 ) ;
assign n5941 =  ( n5490 ) ? ( VREG_14_1 ) : ( n5940 ) ;
assign n5942 =  ( n5489 ) ? ( VREG_14_2 ) : ( n5941 ) ;
assign n5943 =  ( n5488 ) ? ( VREG_14_3 ) : ( n5942 ) ;
assign n5944 =  ( n5487 ) ? ( VREG_14_4 ) : ( n5943 ) ;
assign n5945 =  ( n5486 ) ? ( VREG_14_5 ) : ( n5944 ) ;
assign n5946 =  ( n5485 ) ? ( VREG_14_6 ) : ( n5945 ) ;
assign n5947 =  ( n5484 ) ? ( VREG_14_7 ) : ( n5946 ) ;
assign n5948 =  ( n5483 ) ? ( VREG_14_8 ) : ( n5947 ) ;
assign n5949 =  ( n5482 ) ? ( VREG_14_9 ) : ( n5948 ) ;
assign n5950 =  ( n5481 ) ? ( VREG_14_10 ) : ( n5949 ) ;
assign n5951 =  ( n5480 ) ? ( VREG_14_11 ) : ( n5950 ) ;
assign n5952 =  ( n5479 ) ? ( VREG_14_12 ) : ( n5951 ) ;
assign n5953 =  ( n5478 ) ? ( VREG_14_13 ) : ( n5952 ) ;
assign n5954 =  ( n5477 ) ? ( VREG_14_14 ) : ( n5953 ) ;
assign n5955 =  ( n5476 ) ? ( VREG_14_15 ) : ( n5954 ) ;
assign n5956 =  ( n5475 ) ? ( VREG_15_0 ) : ( n5955 ) ;
assign n5957 =  ( n5474 ) ? ( VREG_15_1 ) : ( n5956 ) ;
assign n5958 =  ( n5473 ) ? ( VREG_15_2 ) : ( n5957 ) ;
assign n5959 =  ( n5472 ) ? ( VREG_15_3 ) : ( n5958 ) ;
assign n5960 =  ( n5471 ) ? ( VREG_15_4 ) : ( n5959 ) ;
assign n5961 =  ( n5470 ) ? ( VREG_15_5 ) : ( n5960 ) ;
assign n5962 =  ( n5469 ) ? ( VREG_15_6 ) : ( n5961 ) ;
assign n5963 =  ( n5468 ) ? ( VREG_15_7 ) : ( n5962 ) ;
assign n5964 =  ( n5467 ) ? ( VREG_15_8 ) : ( n5963 ) ;
assign n5965 =  ( n5466 ) ? ( VREG_15_9 ) : ( n5964 ) ;
assign n5966 =  ( n5465 ) ? ( VREG_15_10 ) : ( n5965 ) ;
assign n5967 =  ( n5464 ) ? ( VREG_15_11 ) : ( n5966 ) ;
assign n5968 =  ( n5463 ) ? ( VREG_15_12 ) : ( n5967 ) ;
assign n5969 =  ( n5462 ) ? ( VREG_15_13 ) : ( n5968 ) ;
assign n5970 =  ( n5461 ) ? ( VREG_15_14 ) : ( n5969 ) ;
assign n5971 =  ( n5460 ) ? ( VREG_15_15 ) : ( n5970 ) ;
assign n5972 =  ( n5459 ) ? ( VREG_16_0 ) : ( n5971 ) ;
assign n5973 =  ( n5458 ) ? ( VREG_16_1 ) : ( n5972 ) ;
assign n5974 =  ( n5457 ) ? ( VREG_16_2 ) : ( n5973 ) ;
assign n5975 =  ( n5456 ) ? ( VREG_16_3 ) : ( n5974 ) ;
assign n5976 =  ( n5455 ) ? ( VREG_16_4 ) : ( n5975 ) ;
assign n5977 =  ( n5454 ) ? ( VREG_16_5 ) : ( n5976 ) ;
assign n5978 =  ( n5453 ) ? ( VREG_16_6 ) : ( n5977 ) ;
assign n5979 =  ( n5452 ) ? ( VREG_16_7 ) : ( n5978 ) ;
assign n5980 =  ( n5451 ) ? ( VREG_16_8 ) : ( n5979 ) ;
assign n5981 =  ( n5450 ) ? ( VREG_16_9 ) : ( n5980 ) ;
assign n5982 =  ( n5449 ) ? ( VREG_16_10 ) : ( n5981 ) ;
assign n5983 =  ( n5448 ) ? ( VREG_16_11 ) : ( n5982 ) ;
assign n5984 =  ( n5447 ) ? ( VREG_16_12 ) : ( n5983 ) ;
assign n5985 =  ( n5446 ) ? ( VREG_16_13 ) : ( n5984 ) ;
assign n5986 =  ( n5445 ) ? ( VREG_16_14 ) : ( n5985 ) ;
assign n5987 =  ( n5444 ) ? ( VREG_16_15 ) : ( n5986 ) ;
assign n5988 =  ( n5443 ) ? ( VREG_17_0 ) : ( n5987 ) ;
assign n5989 =  ( n5442 ) ? ( VREG_17_1 ) : ( n5988 ) ;
assign n5990 =  ( n5441 ) ? ( VREG_17_2 ) : ( n5989 ) ;
assign n5991 =  ( n5440 ) ? ( VREG_17_3 ) : ( n5990 ) ;
assign n5992 =  ( n5439 ) ? ( VREG_17_4 ) : ( n5991 ) ;
assign n5993 =  ( n5438 ) ? ( VREG_17_5 ) : ( n5992 ) ;
assign n5994 =  ( n5437 ) ? ( VREG_17_6 ) : ( n5993 ) ;
assign n5995 =  ( n5436 ) ? ( VREG_17_7 ) : ( n5994 ) ;
assign n5996 =  ( n5435 ) ? ( VREG_17_8 ) : ( n5995 ) ;
assign n5997 =  ( n5434 ) ? ( VREG_17_9 ) : ( n5996 ) ;
assign n5998 =  ( n5433 ) ? ( VREG_17_10 ) : ( n5997 ) ;
assign n5999 =  ( n5432 ) ? ( VREG_17_11 ) : ( n5998 ) ;
assign n6000 =  ( n5431 ) ? ( VREG_17_12 ) : ( n5999 ) ;
assign n6001 =  ( n5430 ) ? ( VREG_17_13 ) : ( n6000 ) ;
assign n6002 =  ( n5429 ) ? ( VREG_17_14 ) : ( n6001 ) ;
assign n6003 =  ( n5428 ) ? ( VREG_17_15 ) : ( n6002 ) ;
assign n6004 =  ( n5427 ) ? ( VREG_18_0 ) : ( n6003 ) ;
assign n6005 =  ( n5426 ) ? ( VREG_18_1 ) : ( n6004 ) ;
assign n6006 =  ( n5425 ) ? ( VREG_18_2 ) : ( n6005 ) ;
assign n6007 =  ( n5424 ) ? ( VREG_18_3 ) : ( n6006 ) ;
assign n6008 =  ( n5423 ) ? ( VREG_18_4 ) : ( n6007 ) ;
assign n6009 =  ( n5422 ) ? ( VREG_18_5 ) : ( n6008 ) ;
assign n6010 =  ( n5421 ) ? ( VREG_18_6 ) : ( n6009 ) ;
assign n6011 =  ( n5420 ) ? ( VREG_18_7 ) : ( n6010 ) ;
assign n6012 =  ( n5419 ) ? ( VREG_18_8 ) : ( n6011 ) ;
assign n6013 =  ( n5418 ) ? ( VREG_18_9 ) : ( n6012 ) ;
assign n6014 =  ( n5417 ) ? ( VREG_18_10 ) : ( n6013 ) ;
assign n6015 =  ( n5416 ) ? ( VREG_18_11 ) : ( n6014 ) ;
assign n6016 =  ( n5415 ) ? ( VREG_18_12 ) : ( n6015 ) ;
assign n6017 =  ( n5414 ) ? ( VREG_18_13 ) : ( n6016 ) ;
assign n6018 =  ( n5413 ) ? ( VREG_18_14 ) : ( n6017 ) ;
assign n6019 =  ( n5412 ) ? ( VREG_18_15 ) : ( n6018 ) ;
assign n6020 =  ( n5411 ) ? ( VREG_19_0 ) : ( n6019 ) ;
assign n6021 =  ( n5410 ) ? ( VREG_19_1 ) : ( n6020 ) ;
assign n6022 =  ( n5409 ) ? ( VREG_19_2 ) : ( n6021 ) ;
assign n6023 =  ( n5408 ) ? ( VREG_19_3 ) : ( n6022 ) ;
assign n6024 =  ( n5407 ) ? ( VREG_19_4 ) : ( n6023 ) ;
assign n6025 =  ( n5406 ) ? ( VREG_19_5 ) : ( n6024 ) ;
assign n6026 =  ( n5405 ) ? ( VREG_19_6 ) : ( n6025 ) ;
assign n6027 =  ( n5404 ) ? ( VREG_19_7 ) : ( n6026 ) ;
assign n6028 =  ( n5403 ) ? ( VREG_19_8 ) : ( n6027 ) ;
assign n6029 =  ( n5402 ) ? ( VREG_19_9 ) : ( n6028 ) ;
assign n6030 =  ( n5401 ) ? ( VREG_19_10 ) : ( n6029 ) ;
assign n6031 =  ( n5400 ) ? ( VREG_19_11 ) : ( n6030 ) ;
assign n6032 =  ( n5399 ) ? ( VREG_19_12 ) : ( n6031 ) ;
assign n6033 =  ( n5398 ) ? ( VREG_19_13 ) : ( n6032 ) ;
assign n6034 =  ( n5397 ) ? ( VREG_19_14 ) : ( n6033 ) ;
assign n6035 =  ( n5396 ) ? ( VREG_19_15 ) : ( n6034 ) ;
assign n6036 =  ( n5395 ) ? ( VREG_20_0 ) : ( n6035 ) ;
assign n6037 =  ( n5394 ) ? ( VREG_20_1 ) : ( n6036 ) ;
assign n6038 =  ( n5393 ) ? ( VREG_20_2 ) : ( n6037 ) ;
assign n6039 =  ( n5392 ) ? ( VREG_20_3 ) : ( n6038 ) ;
assign n6040 =  ( n5391 ) ? ( VREG_20_4 ) : ( n6039 ) ;
assign n6041 =  ( n5390 ) ? ( VREG_20_5 ) : ( n6040 ) ;
assign n6042 =  ( n5389 ) ? ( VREG_20_6 ) : ( n6041 ) ;
assign n6043 =  ( n5388 ) ? ( VREG_20_7 ) : ( n6042 ) ;
assign n6044 =  ( n5387 ) ? ( VREG_20_8 ) : ( n6043 ) ;
assign n6045 =  ( n5386 ) ? ( VREG_20_9 ) : ( n6044 ) ;
assign n6046 =  ( n5385 ) ? ( VREG_20_10 ) : ( n6045 ) ;
assign n6047 =  ( n5384 ) ? ( VREG_20_11 ) : ( n6046 ) ;
assign n6048 =  ( n5383 ) ? ( VREG_20_12 ) : ( n6047 ) ;
assign n6049 =  ( n5382 ) ? ( VREG_20_13 ) : ( n6048 ) ;
assign n6050 =  ( n5381 ) ? ( VREG_20_14 ) : ( n6049 ) ;
assign n6051 =  ( n5380 ) ? ( VREG_20_15 ) : ( n6050 ) ;
assign n6052 =  ( n5379 ) ? ( VREG_21_0 ) : ( n6051 ) ;
assign n6053 =  ( n5378 ) ? ( VREG_21_1 ) : ( n6052 ) ;
assign n6054 =  ( n5377 ) ? ( VREG_21_2 ) : ( n6053 ) ;
assign n6055 =  ( n5376 ) ? ( VREG_21_3 ) : ( n6054 ) ;
assign n6056 =  ( n5375 ) ? ( VREG_21_4 ) : ( n6055 ) ;
assign n6057 =  ( n5374 ) ? ( VREG_21_5 ) : ( n6056 ) ;
assign n6058 =  ( n5373 ) ? ( VREG_21_6 ) : ( n6057 ) ;
assign n6059 =  ( n5372 ) ? ( VREG_21_7 ) : ( n6058 ) ;
assign n6060 =  ( n5371 ) ? ( VREG_21_8 ) : ( n6059 ) ;
assign n6061 =  ( n5370 ) ? ( VREG_21_9 ) : ( n6060 ) ;
assign n6062 =  ( n5369 ) ? ( VREG_21_10 ) : ( n6061 ) ;
assign n6063 =  ( n5368 ) ? ( VREG_21_11 ) : ( n6062 ) ;
assign n6064 =  ( n5367 ) ? ( VREG_21_12 ) : ( n6063 ) ;
assign n6065 =  ( n5366 ) ? ( VREG_21_13 ) : ( n6064 ) ;
assign n6066 =  ( n5365 ) ? ( VREG_21_14 ) : ( n6065 ) ;
assign n6067 =  ( n5364 ) ? ( VREG_21_15 ) : ( n6066 ) ;
assign n6068 =  ( n5363 ) ? ( VREG_22_0 ) : ( n6067 ) ;
assign n6069 =  ( n5362 ) ? ( VREG_22_1 ) : ( n6068 ) ;
assign n6070 =  ( n5361 ) ? ( VREG_22_2 ) : ( n6069 ) ;
assign n6071 =  ( n5360 ) ? ( VREG_22_3 ) : ( n6070 ) ;
assign n6072 =  ( n5359 ) ? ( VREG_22_4 ) : ( n6071 ) ;
assign n6073 =  ( n5358 ) ? ( VREG_22_5 ) : ( n6072 ) ;
assign n6074 =  ( n5357 ) ? ( VREG_22_6 ) : ( n6073 ) ;
assign n6075 =  ( n5356 ) ? ( VREG_22_7 ) : ( n6074 ) ;
assign n6076 =  ( n5355 ) ? ( VREG_22_8 ) : ( n6075 ) ;
assign n6077 =  ( n5354 ) ? ( VREG_22_9 ) : ( n6076 ) ;
assign n6078 =  ( n5353 ) ? ( VREG_22_10 ) : ( n6077 ) ;
assign n6079 =  ( n5352 ) ? ( VREG_22_11 ) : ( n6078 ) ;
assign n6080 =  ( n5351 ) ? ( VREG_22_12 ) : ( n6079 ) ;
assign n6081 =  ( n5350 ) ? ( VREG_22_13 ) : ( n6080 ) ;
assign n6082 =  ( n5349 ) ? ( VREG_22_14 ) : ( n6081 ) ;
assign n6083 =  ( n5348 ) ? ( VREG_22_15 ) : ( n6082 ) ;
assign n6084 =  ( n5347 ) ? ( VREG_23_0 ) : ( n6083 ) ;
assign n6085 =  ( n5346 ) ? ( VREG_23_1 ) : ( n6084 ) ;
assign n6086 =  ( n5345 ) ? ( VREG_23_2 ) : ( n6085 ) ;
assign n6087 =  ( n5344 ) ? ( VREG_23_3 ) : ( n6086 ) ;
assign n6088 =  ( n5343 ) ? ( VREG_23_4 ) : ( n6087 ) ;
assign n6089 =  ( n5342 ) ? ( VREG_23_5 ) : ( n6088 ) ;
assign n6090 =  ( n5341 ) ? ( VREG_23_6 ) : ( n6089 ) ;
assign n6091 =  ( n5340 ) ? ( VREG_23_7 ) : ( n6090 ) ;
assign n6092 =  ( n5339 ) ? ( VREG_23_8 ) : ( n6091 ) ;
assign n6093 =  ( n5338 ) ? ( VREG_23_9 ) : ( n6092 ) ;
assign n6094 =  ( n5337 ) ? ( VREG_23_10 ) : ( n6093 ) ;
assign n6095 =  ( n5336 ) ? ( VREG_23_11 ) : ( n6094 ) ;
assign n6096 =  ( n5335 ) ? ( VREG_23_12 ) : ( n6095 ) ;
assign n6097 =  ( n5334 ) ? ( VREG_23_13 ) : ( n6096 ) ;
assign n6098 =  ( n5333 ) ? ( VREG_23_14 ) : ( n6097 ) ;
assign n6099 =  ( n5332 ) ? ( VREG_23_15 ) : ( n6098 ) ;
assign n6100 =  ( n5331 ) ? ( VREG_24_0 ) : ( n6099 ) ;
assign n6101 =  ( n5330 ) ? ( VREG_24_1 ) : ( n6100 ) ;
assign n6102 =  ( n5329 ) ? ( VREG_24_2 ) : ( n6101 ) ;
assign n6103 =  ( n5328 ) ? ( VREG_24_3 ) : ( n6102 ) ;
assign n6104 =  ( n5327 ) ? ( VREG_24_4 ) : ( n6103 ) ;
assign n6105 =  ( n5326 ) ? ( VREG_24_5 ) : ( n6104 ) ;
assign n6106 =  ( n5325 ) ? ( VREG_24_6 ) : ( n6105 ) ;
assign n6107 =  ( n5324 ) ? ( VREG_24_7 ) : ( n6106 ) ;
assign n6108 =  ( n5323 ) ? ( VREG_24_8 ) : ( n6107 ) ;
assign n6109 =  ( n5322 ) ? ( VREG_24_9 ) : ( n6108 ) ;
assign n6110 =  ( n5321 ) ? ( VREG_24_10 ) : ( n6109 ) ;
assign n6111 =  ( n5320 ) ? ( VREG_24_11 ) : ( n6110 ) ;
assign n6112 =  ( n5319 ) ? ( VREG_24_12 ) : ( n6111 ) ;
assign n6113 =  ( n5318 ) ? ( VREG_24_13 ) : ( n6112 ) ;
assign n6114 =  ( n5317 ) ? ( VREG_24_14 ) : ( n6113 ) ;
assign n6115 =  ( n5316 ) ? ( VREG_24_15 ) : ( n6114 ) ;
assign n6116 =  ( n5315 ) ? ( VREG_25_0 ) : ( n6115 ) ;
assign n6117 =  ( n5314 ) ? ( VREG_25_1 ) : ( n6116 ) ;
assign n6118 =  ( n5313 ) ? ( VREG_25_2 ) : ( n6117 ) ;
assign n6119 =  ( n5312 ) ? ( VREG_25_3 ) : ( n6118 ) ;
assign n6120 =  ( n5311 ) ? ( VREG_25_4 ) : ( n6119 ) ;
assign n6121 =  ( n5310 ) ? ( VREG_25_5 ) : ( n6120 ) ;
assign n6122 =  ( n5309 ) ? ( VREG_25_6 ) : ( n6121 ) ;
assign n6123 =  ( n5308 ) ? ( VREG_25_7 ) : ( n6122 ) ;
assign n6124 =  ( n5307 ) ? ( VREG_25_8 ) : ( n6123 ) ;
assign n6125 =  ( n5306 ) ? ( VREG_25_9 ) : ( n6124 ) ;
assign n6126 =  ( n5305 ) ? ( VREG_25_10 ) : ( n6125 ) ;
assign n6127 =  ( n5304 ) ? ( VREG_25_11 ) : ( n6126 ) ;
assign n6128 =  ( n5303 ) ? ( VREG_25_12 ) : ( n6127 ) ;
assign n6129 =  ( n5302 ) ? ( VREG_25_13 ) : ( n6128 ) ;
assign n6130 =  ( n5301 ) ? ( VREG_25_14 ) : ( n6129 ) ;
assign n6131 =  ( n5300 ) ? ( VREG_25_15 ) : ( n6130 ) ;
assign n6132 =  ( n5299 ) ? ( VREG_26_0 ) : ( n6131 ) ;
assign n6133 =  ( n5298 ) ? ( VREG_26_1 ) : ( n6132 ) ;
assign n6134 =  ( n5297 ) ? ( VREG_26_2 ) : ( n6133 ) ;
assign n6135 =  ( n5296 ) ? ( VREG_26_3 ) : ( n6134 ) ;
assign n6136 =  ( n5295 ) ? ( VREG_26_4 ) : ( n6135 ) ;
assign n6137 =  ( n5294 ) ? ( VREG_26_5 ) : ( n6136 ) ;
assign n6138 =  ( n5293 ) ? ( VREG_26_6 ) : ( n6137 ) ;
assign n6139 =  ( n5292 ) ? ( VREG_26_7 ) : ( n6138 ) ;
assign n6140 =  ( n5291 ) ? ( VREG_26_8 ) : ( n6139 ) ;
assign n6141 =  ( n5290 ) ? ( VREG_26_9 ) : ( n6140 ) ;
assign n6142 =  ( n5289 ) ? ( VREG_26_10 ) : ( n6141 ) ;
assign n6143 =  ( n5288 ) ? ( VREG_26_11 ) : ( n6142 ) ;
assign n6144 =  ( n5287 ) ? ( VREG_26_12 ) : ( n6143 ) ;
assign n6145 =  ( n5286 ) ? ( VREG_26_13 ) : ( n6144 ) ;
assign n6146 =  ( n5285 ) ? ( VREG_26_14 ) : ( n6145 ) ;
assign n6147 =  ( n5284 ) ? ( VREG_26_15 ) : ( n6146 ) ;
assign n6148 =  ( n5283 ) ? ( VREG_27_0 ) : ( n6147 ) ;
assign n6149 =  ( n5282 ) ? ( VREG_27_1 ) : ( n6148 ) ;
assign n6150 =  ( n5281 ) ? ( VREG_27_2 ) : ( n6149 ) ;
assign n6151 =  ( n5280 ) ? ( VREG_27_3 ) : ( n6150 ) ;
assign n6152 =  ( n5279 ) ? ( VREG_27_4 ) : ( n6151 ) ;
assign n6153 =  ( n5278 ) ? ( VREG_27_5 ) : ( n6152 ) ;
assign n6154 =  ( n5277 ) ? ( VREG_27_6 ) : ( n6153 ) ;
assign n6155 =  ( n5276 ) ? ( VREG_27_7 ) : ( n6154 ) ;
assign n6156 =  ( n5275 ) ? ( VREG_27_8 ) : ( n6155 ) ;
assign n6157 =  ( n5274 ) ? ( VREG_27_9 ) : ( n6156 ) ;
assign n6158 =  ( n5273 ) ? ( VREG_27_10 ) : ( n6157 ) ;
assign n6159 =  ( n5272 ) ? ( VREG_27_11 ) : ( n6158 ) ;
assign n6160 =  ( n5271 ) ? ( VREG_27_12 ) : ( n6159 ) ;
assign n6161 =  ( n5270 ) ? ( VREG_27_13 ) : ( n6160 ) ;
assign n6162 =  ( n5269 ) ? ( VREG_27_14 ) : ( n6161 ) ;
assign n6163 =  ( n5268 ) ? ( VREG_27_15 ) : ( n6162 ) ;
assign n6164 =  ( n5267 ) ? ( VREG_28_0 ) : ( n6163 ) ;
assign n6165 =  ( n5266 ) ? ( VREG_28_1 ) : ( n6164 ) ;
assign n6166 =  ( n5265 ) ? ( VREG_28_2 ) : ( n6165 ) ;
assign n6167 =  ( n5264 ) ? ( VREG_28_3 ) : ( n6166 ) ;
assign n6168 =  ( n5263 ) ? ( VREG_28_4 ) : ( n6167 ) ;
assign n6169 =  ( n5262 ) ? ( VREG_28_5 ) : ( n6168 ) ;
assign n6170 =  ( n5261 ) ? ( VREG_28_6 ) : ( n6169 ) ;
assign n6171 =  ( n5260 ) ? ( VREG_28_7 ) : ( n6170 ) ;
assign n6172 =  ( n5259 ) ? ( VREG_28_8 ) : ( n6171 ) ;
assign n6173 =  ( n5258 ) ? ( VREG_28_9 ) : ( n6172 ) ;
assign n6174 =  ( n5257 ) ? ( VREG_28_10 ) : ( n6173 ) ;
assign n6175 =  ( n5256 ) ? ( VREG_28_11 ) : ( n6174 ) ;
assign n6176 =  ( n5255 ) ? ( VREG_28_12 ) : ( n6175 ) ;
assign n6177 =  ( n5254 ) ? ( VREG_28_13 ) : ( n6176 ) ;
assign n6178 =  ( n5253 ) ? ( VREG_28_14 ) : ( n6177 ) ;
assign n6179 =  ( n5252 ) ? ( VREG_28_15 ) : ( n6178 ) ;
assign n6180 =  ( n5251 ) ? ( VREG_29_0 ) : ( n6179 ) ;
assign n6181 =  ( n5250 ) ? ( VREG_29_1 ) : ( n6180 ) ;
assign n6182 =  ( n5249 ) ? ( VREG_29_2 ) : ( n6181 ) ;
assign n6183 =  ( n5248 ) ? ( VREG_29_3 ) : ( n6182 ) ;
assign n6184 =  ( n5247 ) ? ( VREG_29_4 ) : ( n6183 ) ;
assign n6185 =  ( n5246 ) ? ( VREG_29_5 ) : ( n6184 ) ;
assign n6186 =  ( n5245 ) ? ( VREG_29_6 ) : ( n6185 ) ;
assign n6187 =  ( n5244 ) ? ( VREG_29_7 ) : ( n6186 ) ;
assign n6188 =  ( n5243 ) ? ( VREG_29_8 ) : ( n6187 ) ;
assign n6189 =  ( n5242 ) ? ( VREG_29_9 ) : ( n6188 ) ;
assign n6190 =  ( n5241 ) ? ( VREG_29_10 ) : ( n6189 ) ;
assign n6191 =  ( n5240 ) ? ( VREG_29_11 ) : ( n6190 ) ;
assign n6192 =  ( n5239 ) ? ( VREG_29_12 ) : ( n6191 ) ;
assign n6193 =  ( n5238 ) ? ( VREG_29_13 ) : ( n6192 ) ;
assign n6194 =  ( n5237 ) ? ( VREG_29_14 ) : ( n6193 ) ;
assign n6195 =  ( n5236 ) ? ( VREG_29_15 ) : ( n6194 ) ;
assign n6196 =  ( n5235 ) ? ( VREG_30_0 ) : ( n6195 ) ;
assign n6197 =  ( n5234 ) ? ( VREG_30_1 ) : ( n6196 ) ;
assign n6198 =  ( n5233 ) ? ( VREG_30_2 ) : ( n6197 ) ;
assign n6199 =  ( n5232 ) ? ( VREG_30_3 ) : ( n6198 ) ;
assign n6200 =  ( n5231 ) ? ( VREG_30_4 ) : ( n6199 ) ;
assign n6201 =  ( n5230 ) ? ( VREG_30_5 ) : ( n6200 ) ;
assign n6202 =  ( n5229 ) ? ( VREG_30_6 ) : ( n6201 ) ;
assign n6203 =  ( n5228 ) ? ( VREG_30_7 ) : ( n6202 ) ;
assign n6204 =  ( n5227 ) ? ( VREG_30_8 ) : ( n6203 ) ;
assign n6205 =  ( n5226 ) ? ( VREG_30_9 ) : ( n6204 ) ;
assign n6206 =  ( n5225 ) ? ( VREG_30_10 ) : ( n6205 ) ;
assign n6207 =  ( n5224 ) ? ( VREG_30_11 ) : ( n6206 ) ;
assign n6208 =  ( n5223 ) ? ( VREG_30_12 ) : ( n6207 ) ;
assign n6209 =  ( n5222 ) ? ( VREG_30_13 ) : ( n6208 ) ;
assign n6210 =  ( n5221 ) ? ( VREG_30_14 ) : ( n6209 ) ;
assign n6211 =  ( n5220 ) ? ( VREG_30_15 ) : ( n6210 ) ;
assign n6212 =  ( n5219 ) ? ( VREG_31_0 ) : ( n6211 ) ;
assign n6213 =  ( n5217 ) ? ( VREG_31_1 ) : ( n6212 ) ;
assign n6214 =  ( n5215 ) ? ( VREG_31_2 ) : ( n6213 ) ;
assign n6215 =  ( n5213 ) ? ( VREG_31_3 ) : ( n6214 ) ;
assign n6216 =  ( n5211 ) ? ( VREG_31_4 ) : ( n6215 ) ;
assign n6217 =  ( n5209 ) ? ( VREG_31_5 ) : ( n6216 ) ;
assign n6218 =  ( n5207 ) ? ( VREG_31_6 ) : ( n6217 ) ;
assign n6219 =  ( n5205 ) ? ( VREG_31_7 ) : ( n6218 ) ;
assign n6220 =  ( n5203 ) ? ( VREG_31_8 ) : ( n6219 ) ;
assign n6221 =  ( n5201 ) ? ( VREG_31_9 ) : ( n6220 ) ;
assign n6222 =  ( n5199 ) ? ( VREG_31_10 ) : ( n6221 ) ;
assign n6223 =  ( n5197 ) ? ( VREG_31_11 ) : ( n6222 ) ;
assign n6224 =  ( n5195 ) ? ( VREG_31_12 ) : ( n6223 ) ;
assign n6225 =  ( n5193 ) ? ( VREG_31_13 ) : ( n6224 ) ;
assign n6226 =  ( n5191 ) ? ( VREG_31_14 ) : ( n6225 ) ;
assign n6227 =  ( n5189 ) ? ( VREG_31_15 ) : ( n6226 ) ;
assign n6228 =  ( n6227 ) + ( n140 )  ;
assign n6229 =  ( n6227 ) - ( n140 )  ;
assign n6230 =  ( n6227 ) & ( n140 )  ;
assign n6231 =  ( n6227 ) | ( n140 )  ;
assign n6232 =  ( ( n6227 ) * ( n140 ))  ;
assign n6233 =  ( n148 ) ? ( n6232 ) : ( VREG_0_10 ) ;
assign n6234 =  ( n146 ) ? ( n6231 ) : ( n6233 ) ;
assign n6235 =  ( n144 ) ? ( n6230 ) : ( n6234 ) ;
assign n6236 =  ( n142 ) ? ( n6229 ) : ( n6235 ) ;
assign n6237 =  ( n10 ) ? ( n6228 ) : ( n6236 ) ;
assign n6238 =  ( n77 ) & ( n5188 )  ;
assign n6239 =  ( n77 ) & ( n5190 )  ;
assign n6240 =  ( n77 ) & ( n5192 )  ;
assign n6241 =  ( n77 ) & ( n5194 )  ;
assign n6242 =  ( n77 ) & ( n5196 )  ;
assign n6243 =  ( n77 ) & ( n5198 )  ;
assign n6244 =  ( n77 ) & ( n5200 )  ;
assign n6245 =  ( n77 ) & ( n5202 )  ;
assign n6246 =  ( n77 ) & ( n5204 )  ;
assign n6247 =  ( n77 ) & ( n5206 )  ;
assign n6248 =  ( n77 ) & ( n5208 )  ;
assign n6249 =  ( n77 ) & ( n5210 )  ;
assign n6250 =  ( n77 ) & ( n5212 )  ;
assign n6251 =  ( n77 ) & ( n5214 )  ;
assign n6252 =  ( n77 ) & ( n5216 )  ;
assign n6253 =  ( n77 ) & ( n5218 )  ;
assign n6254 =  ( n78 ) & ( n5188 )  ;
assign n6255 =  ( n78 ) & ( n5190 )  ;
assign n6256 =  ( n78 ) & ( n5192 )  ;
assign n6257 =  ( n78 ) & ( n5194 )  ;
assign n6258 =  ( n78 ) & ( n5196 )  ;
assign n6259 =  ( n78 ) & ( n5198 )  ;
assign n6260 =  ( n78 ) & ( n5200 )  ;
assign n6261 =  ( n78 ) & ( n5202 )  ;
assign n6262 =  ( n78 ) & ( n5204 )  ;
assign n6263 =  ( n78 ) & ( n5206 )  ;
assign n6264 =  ( n78 ) & ( n5208 )  ;
assign n6265 =  ( n78 ) & ( n5210 )  ;
assign n6266 =  ( n78 ) & ( n5212 )  ;
assign n6267 =  ( n78 ) & ( n5214 )  ;
assign n6268 =  ( n78 ) & ( n5216 )  ;
assign n6269 =  ( n78 ) & ( n5218 )  ;
assign n6270 =  ( n79 ) & ( n5188 )  ;
assign n6271 =  ( n79 ) & ( n5190 )  ;
assign n6272 =  ( n79 ) & ( n5192 )  ;
assign n6273 =  ( n79 ) & ( n5194 )  ;
assign n6274 =  ( n79 ) & ( n5196 )  ;
assign n6275 =  ( n79 ) & ( n5198 )  ;
assign n6276 =  ( n79 ) & ( n5200 )  ;
assign n6277 =  ( n79 ) & ( n5202 )  ;
assign n6278 =  ( n79 ) & ( n5204 )  ;
assign n6279 =  ( n79 ) & ( n5206 )  ;
assign n6280 =  ( n79 ) & ( n5208 )  ;
assign n6281 =  ( n79 ) & ( n5210 )  ;
assign n6282 =  ( n79 ) & ( n5212 )  ;
assign n6283 =  ( n79 ) & ( n5214 )  ;
assign n6284 =  ( n79 ) & ( n5216 )  ;
assign n6285 =  ( n79 ) & ( n5218 )  ;
assign n6286 =  ( n80 ) & ( n5188 )  ;
assign n6287 =  ( n80 ) & ( n5190 )  ;
assign n6288 =  ( n80 ) & ( n5192 )  ;
assign n6289 =  ( n80 ) & ( n5194 )  ;
assign n6290 =  ( n80 ) & ( n5196 )  ;
assign n6291 =  ( n80 ) & ( n5198 )  ;
assign n6292 =  ( n80 ) & ( n5200 )  ;
assign n6293 =  ( n80 ) & ( n5202 )  ;
assign n6294 =  ( n80 ) & ( n5204 )  ;
assign n6295 =  ( n80 ) & ( n5206 )  ;
assign n6296 =  ( n80 ) & ( n5208 )  ;
assign n6297 =  ( n80 ) & ( n5210 )  ;
assign n6298 =  ( n80 ) & ( n5212 )  ;
assign n6299 =  ( n80 ) & ( n5214 )  ;
assign n6300 =  ( n80 ) & ( n5216 )  ;
assign n6301 =  ( n80 ) & ( n5218 )  ;
assign n6302 =  ( n81 ) & ( n5188 )  ;
assign n6303 =  ( n81 ) & ( n5190 )  ;
assign n6304 =  ( n81 ) & ( n5192 )  ;
assign n6305 =  ( n81 ) & ( n5194 )  ;
assign n6306 =  ( n81 ) & ( n5196 )  ;
assign n6307 =  ( n81 ) & ( n5198 )  ;
assign n6308 =  ( n81 ) & ( n5200 )  ;
assign n6309 =  ( n81 ) & ( n5202 )  ;
assign n6310 =  ( n81 ) & ( n5204 )  ;
assign n6311 =  ( n81 ) & ( n5206 )  ;
assign n6312 =  ( n81 ) & ( n5208 )  ;
assign n6313 =  ( n81 ) & ( n5210 )  ;
assign n6314 =  ( n81 ) & ( n5212 )  ;
assign n6315 =  ( n81 ) & ( n5214 )  ;
assign n6316 =  ( n81 ) & ( n5216 )  ;
assign n6317 =  ( n81 ) & ( n5218 )  ;
assign n6318 =  ( n82 ) & ( n5188 )  ;
assign n6319 =  ( n82 ) & ( n5190 )  ;
assign n6320 =  ( n82 ) & ( n5192 )  ;
assign n6321 =  ( n82 ) & ( n5194 )  ;
assign n6322 =  ( n82 ) & ( n5196 )  ;
assign n6323 =  ( n82 ) & ( n5198 )  ;
assign n6324 =  ( n82 ) & ( n5200 )  ;
assign n6325 =  ( n82 ) & ( n5202 )  ;
assign n6326 =  ( n82 ) & ( n5204 )  ;
assign n6327 =  ( n82 ) & ( n5206 )  ;
assign n6328 =  ( n82 ) & ( n5208 )  ;
assign n6329 =  ( n82 ) & ( n5210 )  ;
assign n6330 =  ( n82 ) & ( n5212 )  ;
assign n6331 =  ( n82 ) & ( n5214 )  ;
assign n6332 =  ( n82 ) & ( n5216 )  ;
assign n6333 =  ( n82 ) & ( n5218 )  ;
assign n6334 =  ( n83 ) & ( n5188 )  ;
assign n6335 =  ( n83 ) & ( n5190 )  ;
assign n6336 =  ( n83 ) & ( n5192 )  ;
assign n6337 =  ( n83 ) & ( n5194 )  ;
assign n6338 =  ( n83 ) & ( n5196 )  ;
assign n6339 =  ( n83 ) & ( n5198 )  ;
assign n6340 =  ( n83 ) & ( n5200 )  ;
assign n6341 =  ( n83 ) & ( n5202 )  ;
assign n6342 =  ( n83 ) & ( n5204 )  ;
assign n6343 =  ( n83 ) & ( n5206 )  ;
assign n6344 =  ( n83 ) & ( n5208 )  ;
assign n6345 =  ( n83 ) & ( n5210 )  ;
assign n6346 =  ( n83 ) & ( n5212 )  ;
assign n6347 =  ( n83 ) & ( n5214 )  ;
assign n6348 =  ( n83 ) & ( n5216 )  ;
assign n6349 =  ( n83 ) & ( n5218 )  ;
assign n6350 =  ( n84 ) & ( n5188 )  ;
assign n6351 =  ( n84 ) & ( n5190 )  ;
assign n6352 =  ( n84 ) & ( n5192 )  ;
assign n6353 =  ( n84 ) & ( n5194 )  ;
assign n6354 =  ( n84 ) & ( n5196 )  ;
assign n6355 =  ( n84 ) & ( n5198 )  ;
assign n6356 =  ( n84 ) & ( n5200 )  ;
assign n6357 =  ( n84 ) & ( n5202 )  ;
assign n6358 =  ( n84 ) & ( n5204 )  ;
assign n6359 =  ( n84 ) & ( n5206 )  ;
assign n6360 =  ( n84 ) & ( n5208 )  ;
assign n6361 =  ( n84 ) & ( n5210 )  ;
assign n6362 =  ( n84 ) & ( n5212 )  ;
assign n6363 =  ( n84 ) & ( n5214 )  ;
assign n6364 =  ( n84 ) & ( n5216 )  ;
assign n6365 =  ( n84 ) & ( n5218 )  ;
assign n6366 =  ( n85 ) & ( n5188 )  ;
assign n6367 =  ( n85 ) & ( n5190 )  ;
assign n6368 =  ( n85 ) & ( n5192 )  ;
assign n6369 =  ( n85 ) & ( n5194 )  ;
assign n6370 =  ( n85 ) & ( n5196 )  ;
assign n6371 =  ( n85 ) & ( n5198 )  ;
assign n6372 =  ( n85 ) & ( n5200 )  ;
assign n6373 =  ( n85 ) & ( n5202 )  ;
assign n6374 =  ( n85 ) & ( n5204 )  ;
assign n6375 =  ( n85 ) & ( n5206 )  ;
assign n6376 =  ( n85 ) & ( n5208 )  ;
assign n6377 =  ( n85 ) & ( n5210 )  ;
assign n6378 =  ( n85 ) & ( n5212 )  ;
assign n6379 =  ( n85 ) & ( n5214 )  ;
assign n6380 =  ( n85 ) & ( n5216 )  ;
assign n6381 =  ( n85 ) & ( n5218 )  ;
assign n6382 =  ( n86 ) & ( n5188 )  ;
assign n6383 =  ( n86 ) & ( n5190 )  ;
assign n6384 =  ( n86 ) & ( n5192 )  ;
assign n6385 =  ( n86 ) & ( n5194 )  ;
assign n6386 =  ( n86 ) & ( n5196 )  ;
assign n6387 =  ( n86 ) & ( n5198 )  ;
assign n6388 =  ( n86 ) & ( n5200 )  ;
assign n6389 =  ( n86 ) & ( n5202 )  ;
assign n6390 =  ( n86 ) & ( n5204 )  ;
assign n6391 =  ( n86 ) & ( n5206 )  ;
assign n6392 =  ( n86 ) & ( n5208 )  ;
assign n6393 =  ( n86 ) & ( n5210 )  ;
assign n6394 =  ( n86 ) & ( n5212 )  ;
assign n6395 =  ( n86 ) & ( n5214 )  ;
assign n6396 =  ( n86 ) & ( n5216 )  ;
assign n6397 =  ( n86 ) & ( n5218 )  ;
assign n6398 =  ( n87 ) & ( n5188 )  ;
assign n6399 =  ( n87 ) & ( n5190 )  ;
assign n6400 =  ( n87 ) & ( n5192 )  ;
assign n6401 =  ( n87 ) & ( n5194 )  ;
assign n6402 =  ( n87 ) & ( n5196 )  ;
assign n6403 =  ( n87 ) & ( n5198 )  ;
assign n6404 =  ( n87 ) & ( n5200 )  ;
assign n6405 =  ( n87 ) & ( n5202 )  ;
assign n6406 =  ( n87 ) & ( n5204 )  ;
assign n6407 =  ( n87 ) & ( n5206 )  ;
assign n6408 =  ( n87 ) & ( n5208 )  ;
assign n6409 =  ( n87 ) & ( n5210 )  ;
assign n6410 =  ( n87 ) & ( n5212 )  ;
assign n6411 =  ( n87 ) & ( n5214 )  ;
assign n6412 =  ( n87 ) & ( n5216 )  ;
assign n6413 =  ( n87 ) & ( n5218 )  ;
assign n6414 =  ( n88 ) & ( n5188 )  ;
assign n6415 =  ( n88 ) & ( n5190 )  ;
assign n6416 =  ( n88 ) & ( n5192 )  ;
assign n6417 =  ( n88 ) & ( n5194 )  ;
assign n6418 =  ( n88 ) & ( n5196 )  ;
assign n6419 =  ( n88 ) & ( n5198 )  ;
assign n6420 =  ( n88 ) & ( n5200 )  ;
assign n6421 =  ( n88 ) & ( n5202 )  ;
assign n6422 =  ( n88 ) & ( n5204 )  ;
assign n6423 =  ( n88 ) & ( n5206 )  ;
assign n6424 =  ( n88 ) & ( n5208 )  ;
assign n6425 =  ( n88 ) & ( n5210 )  ;
assign n6426 =  ( n88 ) & ( n5212 )  ;
assign n6427 =  ( n88 ) & ( n5214 )  ;
assign n6428 =  ( n88 ) & ( n5216 )  ;
assign n6429 =  ( n88 ) & ( n5218 )  ;
assign n6430 =  ( n89 ) & ( n5188 )  ;
assign n6431 =  ( n89 ) & ( n5190 )  ;
assign n6432 =  ( n89 ) & ( n5192 )  ;
assign n6433 =  ( n89 ) & ( n5194 )  ;
assign n6434 =  ( n89 ) & ( n5196 )  ;
assign n6435 =  ( n89 ) & ( n5198 )  ;
assign n6436 =  ( n89 ) & ( n5200 )  ;
assign n6437 =  ( n89 ) & ( n5202 )  ;
assign n6438 =  ( n89 ) & ( n5204 )  ;
assign n6439 =  ( n89 ) & ( n5206 )  ;
assign n6440 =  ( n89 ) & ( n5208 )  ;
assign n6441 =  ( n89 ) & ( n5210 )  ;
assign n6442 =  ( n89 ) & ( n5212 )  ;
assign n6443 =  ( n89 ) & ( n5214 )  ;
assign n6444 =  ( n89 ) & ( n5216 )  ;
assign n6445 =  ( n89 ) & ( n5218 )  ;
assign n6446 =  ( n90 ) & ( n5188 )  ;
assign n6447 =  ( n90 ) & ( n5190 )  ;
assign n6448 =  ( n90 ) & ( n5192 )  ;
assign n6449 =  ( n90 ) & ( n5194 )  ;
assign n6450 =  ( n90 ) & ( n5196 )  ;
assign n6451 =  ( n90 ) & ( n5198 )  ;
assign n6452 =  ( n90 ) & ( n5200 )  ;
assign n6453 =  ( n90 ) & ( n5202 )  ;
assign n6454 =  ( n90 ) & ( n5204 )  ;
assign n6455 =  ( n90 ) & ( n5206 )  ;
assign n6456 =  ( n90 ) & ( n5208 )  ;
assign n6457 =  ( n90 ) & ( n5210 )  ;
assign n6458 =  ( n90 ) & ( n5212 )  ;
assign n6459 =  ( n90 ) & ( n5214 )  ;
assign n6460 =  ( n90 ) & ( n5216 )  ;
assign n6461 =  ( n90 ) & ( n5218 )  ;
assign n6462 =  ( n91 ) & ( n5188 )  ;
assign n6463 =  ( n91 ) & ( n5190 )  ;
assign n6464 =  ( n91 ) & ( n5192 )  ;
assign n6465 =  ( n91 ) & ( n5194 )  ;
assign n6466 =  ( n91 ) & ( n5196 )  ;
assign n6467 =  ( n91 ) & ( n5198 )  ;
assign n6468 =  ( n91 ) & ( n5200 )  ;
assign n6469 =  ( n91 ) & ( n5202 )  ;
assign n6470 =  ( n91 ) & ( n5204 )  ;
assign n6471 =  ( n91 ) & ( n5206 )  ;
assign n6472 =  ( n91 ) & ( n5208 )  ;
assign n6473 =  ( n91 ) & ( n5210 )  ;
assign n6474 =  ( n91 ) & ( n5212 )  ;
assign n6475 =  ( n91 ) & ( n5214 )  ;
assign n6476 =  ( n91 ) & ( n5216 )  ;
assign n6477 =  ( n91 ) & ( n5218 )  ;
assign n6478 =  ( n92 ) & ( n5188 )  ;
assign n6479 =  ( n92 ) & ( n5190 )  ;
assign n6480 =  ( n92 ) & ( n5192 )  ;
assign n6481 =  ( n92 ) & ( n5194 )  ;
assign n6482 =  ( n92 ) & ( n5196 )  ;
assign n6483 =  ( n92 ) & ( n5198 )  ;
assign n6484 =  ( n92 ) & ( n5200 )  ;
assign n6485 =  ( n92 ) & ( n5202 )  ;
assign n6486 =  ( n92 ) & ( n5204 )  ;
assign n6487 =  ( n92 ) & ( n5206 )  ;
assign n6488 =  ( n92 ) & ( n5208 )  ;
assign n6489 =  ( n92 ) & ( n5210 )  ;
assign n6490 =  ( n92 ) & ( n5212 )  ;
assign n6491 =  ( n92 ) & ( n5214 )  ;
assign n6492 =  ( n92 ) & ( n5216 )  ;
assign n6493 =  ( n92 ) & ( n5218 )  ;
assign n6494 =  ( n93 ) & ( n5188 )  ;
assign n6495 =  ( n93 ) & ( n5190 )  ;
assign n6496 =  ( n93 ) & ( n5192 )  ;
assign n6497 =  ( n93 ) & ( n5194 )  ;
assign n6498 =  ( n93 ) & ( n5196 )  ;
assign n6499 =  ( n93 ) & ( n5198 )  ;
assign n6500 =  ( n93 ) & ( n5200 )  ;
assign n6501 =  ( n93 ) & ( n5202 )  ;
assign n6502 =  ( n93 ) & ( n5204 )  ;
assign n6503 =  ( n93 ) & ( n5206 )  ;
assign n6504 =  ( n93 ) & ( n5208 )  ;
assign n6505 =  ( n93 ) & ( n5210 )  ;
assign n6506 =  ( n93 ) & ( n5212 )  ;
assign n6507 =  ( n93 ) & ( n5214 )  ;
assign n6508 =  ( n93 ) & ( n5216 )  ;
assign n6509 =  ( n93 ) & ( n5218 )  ;
assign n6510 =  ( n94 ) & ( n5188 )  ;
assign n6511 =  ( n94 ) & ( n5190 )  ;
assign n6512 =  ( n94 ) & ( n5192 )  ;
assign n6513 =  ( n94 ) & ( n5194 )  ;
assign n6514 =  ( n94 ) & ( n5196 )  ;
assign n6515 =  ( n94 ) & ( n5198 )  ;
assign n6516 =  ( n94 ) & ( n5200 )  ;
assign n6517 =  ( n94 ) & ( n5202 )  ;
assign n6518 =  ( n94 ) & ( n5204 )  ;
assign n6519 =  ( n94 ) & ( n5206 )  ;
assign n6520 =  ( n94 ) & ( n5208 )  ;
assign n6521 =  ( n94 ) & ( n5210 )  ;
assign n6522 =  ( n94 ) & ( n5212 )  ;
assign n6523 =  ( n94 ) & ( n5214 )  ;
assign n6524 =  ( n94 ) & ( n5216 )  ;
assign n6525 =  ( n94 ) & ( n5218 )  ;
assign n6526 =  ( n95 ) & ( n5188 )  ;
assign n6527 =  ( n95 ) & ( n5190 )  ;
assign n6528 =  ( n95 ) & ( n5192 )  ;
assign n6529 =  ( n95 ) & ( n5194 )  ;
assign n6530 =  ( n95 ) & ( n5196 )  ;
assign n6531 =  ( n95 ) & ( n5198 )  ;
assign n6532 =  ( n95 ) & ( n5200 )  ;
assign n6533 =  ( n95 ) & ( n5202 )  ;
assign n6534 =  ( n95 ) & ( n5204 )  ;
assign n6535 =  ( n95 ) & ( n5206 )  ;
assign n6536 =  ( n95 ) & ( n5208 )  ;
assign n6537 =  ( n95 ) & ( n5210 )  ;
assign n6538 =  ( n95 ) & ( n5212 )  ;
assign n6539 =  ( n95 ) & ( n5214 )  ;
assign n6540 =  ( n95 ) & ( n5216 )  ;
assign n6541 =  ( n95 ) & ( n5218 )  ;
assign n6542 =  ( n96 ) & ( n5188 )  ;
assign n6543 =  ( n96 ) & ( n5190 )  ;
assign n6544 =  ( n96 ) & ( n5192 )  ;
assign n6545 =  ( n96 ) & ( n5194 )  ;
assign n6546 =  ( n96 ) & ( n5196 )  ;
assign n6547 =  ( n96 ) & ( n5198 )  ;
assign n6548 =  ( n96 ) & ( n5200 )  ;
assign n6549 =  ( n96 ) & ( n5202 )  ;
assign n6550 =  ( n96 ) & ( n5204 )  ;
assign n6551 =  ( n96 ) & ( n5206 )  ;
assign n6552 =  ( n96 ) & ( n5208 )  ;
assign n6553 =  ( n96 ) & ( n5210 )  ;
assign n6554 =  ( n96 ) & ( n5212 )  ;
assign n6555 =  ( n96 ) & ( n5214 )  ;
assign n6556 =  ( n96 ) & ( n5216 )  ;
assign n6557 =  ( n96 ) & ( n5218 )  ;
assign n6558 =  ( n97 ) & ( n5188 )  ;
assign n6559 =  ( n97 ) & ( n5190 )  ;
assign n6560 =  ( n97 ) & ( n5192 )  ;
assign n6561 =  ( n97 ) & ( n5194 )  ;
assign n6562 =  ( n97 ) & ( n5196 )  ;
assign n6563 =  ( n97 ) & ( n5198 )  ;
assign n6564 =  ( n97 ) & ( n5200 )  ;
assign n6565 =  ( n97 ) & ( n5202 )  ;
assign n6566 =  ( n97 ) & ( n5204 )  ;
assign n6567 =  ( n97 ) & ( n5206 )  ;
assign n6568 =  ( n97 ) & ( n5208 )  ;
assign n6569 =  ( n97 ) & ( n5210 )  ;
assign n6570 =  ( n97 ) & ( n5212 )  ;
assign n6571 =  ( n97 ) & ( n5214 )  ;
assign n6572 =  ( n97 ) & ( n5216 )  ;
assign n6573 =  ( n97 ) & ( n5218 )  ;
assign n6574 =  ( n98 ) & ( n5188 )  ;
assign n6575 =  ( n98 ) & ( n5190 )  ;
assign n6576 =  ( n98 ) & ( n5192 )  ;
assign n6577 =  ( n98 ) & ( n5194 )  ;
assign n6578 =  ( n98 ) & ( n5196 )  ;
assign n6579 =  ( n98 ) & ( n5198 )  ;
assign n6580 =  ( n98 ) & ( n5200 )  ;
assign n6581 =  ( n98 ) & ( n5202 )  ;
assign n6582 =  ( n98 ) & ( n5204 )  ;
assign n6583 =  ( n98 ) & ( n5206 )  ;
assign n6584 =  ( n98 ) & ( n5208 )  ;
assign n6585 =  ( n98 ) & ( n5210 )  ;
assign n6586 =  ( n98 ) & ( n5212 )  ;
assign n6587 =  ( n98 ) & ( n5214 )  ;
assign n6588 =  ( n98 ) & ( n5216 )  ;
assign n6589 =  ( n98 ) & ( n5218 )  ;
assign n6590 =  ( n99 ) & ( n5188 )  ;
assign n6591 =  ( n99 ) & ( n5190 )  ;
assign n6592 =  ( n99 ) & ( n5192 )  ;
assign n6593 =  ( n99 ) & ( n5194 )  ;
assign n6594 =  ( n99 ) & ( n5196 )  ;
assign n6595 =  ( n99 ) & ( n5198 )  ;
assign n6596 =  ( n99 ) & ( n5200 )  ;
assign n6597 =  ( n99 ) & ( n5202 )  ;
assign n6598 =  ( n99 ) & ( n5204 )  ;
assign n6599 =  ( n99 ) & ( n5206 )  ;
assign n6600 =  ( n99 ) & ( n5208 )  ;
assign n6601 =  ( n99 ) & ( n5210 )  ;
assign n6602 =  ( n99 ) & ( n5212 )  ;
assign n6603 =  ( n99 ) & ( n5214 )  ;
assign n6604 =  ( n99 ) & ( n5216 )  ;
assign n6605 =  ( n99 ) & ( n5218 )  ;
assign n6606 =  ( n100 ) & ( n5188 )  ;
assign n6607 =  ( n100 ) & ( n5190 )  ;
assign n6608 =  ( n100 ) & ( n5192 )  ;
assign n6609 =  ( n100 ) & ( n5194 )  ;
assign n6610 =  ( n100 ) & ( n5196 )  ;
assign n6611 =  ( n100 ) & ( n5198 )  ;
assign n6612 =  ( n100 ) & ( n5200 )  ;
assign n6613 =  ( n100 ) & ( n5202 )  ;
assign n6614 =  ( n100 ) & ( n5204 )  ;
assign n6615 =  ( n100 ) & ( n5206 )  ;
assign n6616 =  ( n100 ) & ( n5208 )  ;
assign n6617 =  ( n100 ) & ( n5210 )  ;
assign n6618 =  ( n100 ) & ( n5212 )  ;
assign n6619 =  ( n100 ) & ( n5214 )  ;
assign n6620 =  ( n100 ) & ( n5216 )  ;
assign n6621 =  ( n100 ) & ( n5218 )  ;
assign n6622 =  ( n101 ) & ( n5188 )  ;
assign n6623 =  ( n101 ) & ( n5190 )  ;
assign n6624 =  ( n101 ) & ( n5192 )  ;
assign n6625 =  ( n101 ) & ( n5194 )  ;
assign n6626 =  ( n101 ) & ( n5196 )  ;
assign n6627 =  ( n101 ) & ( n5198 )  ;
assign n6628 =  ( n101 ) & ( n5200 )  ;
assign n6629 =  ( n101 ) & ( n5202 )  ;
assign n6630 =  ( n101 ) & ( n5204 )  ;
assign n6631 =  ( n101 ) & ( n5206 )  ;
assign n6632 =  ( n101 ) & ( n5208 )  ;
assign n6633 =  ( n101 ) & ( n5210 )  ;
assign n6634 =  ( n101 ) & ( n5212 )  ;
assign n6635 =  ( n101 ) & ( n5214 )  ;
assign n6636 =  ( n101 ) & ( n5216 )  ;
assign n6637 =  ( n101 ) & ( n5218 )  ;
assign n6638 =  ( n102 ) & ( n5188 )  ;
assign n6639 =  ( n102 ) & ( n5190 )  ;
assign n6640 =  ( n102 ) & ( n5192 )  ;
assign n6641 =  ( n102 ) & ( n5194 )  ;
assign n6642 =  ( n102 ) & ( n5196 )  ;
assign n6643 =  ( n102 ) & ( n5198 )  ;
assign n6644 =  ( n102 ) & ( n5200 )  ;
assign n6645 =  ( n102 ) & ( n5202 )  ;
assign n6646 =  ( n102 ) & ( n5204 )  ;
assign n6647 =  ( n102 ) & ( n5206 )  ;
assign n6648 =  ( n102 ) & ( n5208 )  ;
assign n6649 =  ( n102 ) & ( n5210 )  ;
assign n6650 =  ( n102 ) & ( n5212 )  ;
assign n6651 =  ( n102 ) & ( n5214 )  ;
assign n6652 =  ( n102 ) & ( n5216 )  ;
assign n6653 =  ( n102 ) & ( n5218 )  ;
assign n6654 =  ( n103 ) & ( n5188 )  ;
assign n6655 =  ( n103 ) & ( n5190 )  ;
assign n6656 =  ( n103 ) & ( n5192 )  ;
assign n6657 =  ( n103 ) & ( n5194 )  ;
assign n6658 =  ( n103 ) & ( n5196 )  ;
assign n6659 =  ( n103 ) & ( n5198 )  ;
assign n6660 =  ( n103 ) & ( n5200 )  ;
assign n6661 =  ( n103 ) & ( n5202 )  ;
assign n6662 =  ( n103 ) & ( n5204 )  ;
assign n6663 =  ( n103 ) & ( n5206 )  ;
assign n6664 =  ( n103 ) & ( n5208 )  ;
assign n6665 =  ( n103 ) & ( n5210 )  ;
assign n6666 =  ( n103 ) & ( n5212 )  ;
assign n6667 =  ( n103 ) & ( n5214 )  ;
assign n6668 =  ( n103 ) & ( n5216 )  ;
assign n6669 =  ( n103 ) & ( n5218 )  ;
assign n6670 =  ( n104 ) & ( n5188 )  ;
assign n6671 =  ( n104 ) & ( n5190 )  ;
assign n6672 =  ( n104 ) & ( n5192 )  ;
assign n6673 =  ( n104 ) & ( n5194 )  ;
assign n6674 =  ( n104 ) & ( n5196 )  ;
assign n6675 =  ( n104 ) & ( n5198 )  ;
assign n6676 =  ( n104 ) & ( n5200 )  ;
assign n6677 =  ( n104 ) & ( n5202 )  ;
assign n6678 =  ( n104 ) & ( n5204 )  ;
assign n6679 =  ( n104 ) & ( n5206 )  ;
assign n6680 =  ( n104 ) & ( n5208 )  ;
assign n6681 =  ( n104 ) & ( n5210 )  ;
assign n6682 =  ( n104 ) & ( n5212 )  ;
assign n6683 =  ( n104 ) & ( n5214 )  ;
assign n6684 =  ( n104 ) & ( n5216 )  ;
assign n6685 =  ( n104 ) & ( n5218 )  ;
assign n6686 =  ( n105 ) & ( n5188 )  ;
assign n6687 =  ( n105 ) & ( n5190 )  ;
assign n6688 =  ( n105 ) & ( n5192 )  ;
assign n6689 =  ( n105 ) & ( n5194 )  ;
assign n6690 =  ( n105 ) & ( n5196 )  ;
assign n6691 =  ( n105 ) & ( n5198 )  ;
assign n6692 =  ( n105 ) & ( n5200 )  ;
assign n6693 =  ( n105 ) & ( n5202 )  ;
assign n6694 =  ( n105 ) & ( n5204 )  ;
assign n6695 =  ( n105 ) & ( n5206 )  ;
assign n6696 =  ( n105 ) & ( n5208 )  ;
assign n6697 =  ( n105 ) & ( n5210 )  ;
assign n6698 =  ( n105 ) & ( n5212 )  ;
assign n6699 =  ( n105 ) & ( n5214 )  ;
assign n6700 =  ( n105 ) & ( n5216 )  ;
assign n6701 =  ( n105 ) & ( n5218 )  ;
assign n6702 =  ( n106 ) & ( n5188 )  ;
assign n6703 =  ( n106 ) & ( n5190 )  ;
assign n6704 =  ( n106 ) & ( n5192 )  ;
assign n6705 =  ( n106 ) & ( n5194 )  ;
assign n6706 =  ( n106 ) & ( n5196 )  ;
assign n6707 =  ( n106 ) & ( n5198 )  ;
assign n6708 =  ( n106 ) & ( n5200 )  ;
assign n6709 =  ( n106 ) & ( n5202 )  ;
assign n6710 =  ( n106 ) & ( n5204 )  ;
assign n6711 =  ( n106 ) & ( n5206 )  ;
assign n6712 =  ( n106 ) & ( n5208 )  ;
assign n6713 =  ( n106 ) & ( n5210 )  ;
assign n6714 =  ( n106 ) & ( n5212 )  ;
assign n6715 =  ( n106 ) & ( n5214 )  ;
assign n6716 =  ( n106 ) & ( n5216 )  ;
assign n6717 =  ( n106 ) & ( n5218 )  ;
assign n6718 =  ( n107 ) & ( n5188 )  ;
assign n6719 =  ( n107 ) & ( n5190 )  ;
assign n6720 =  ( n107 ) & ( n5192 )  ;
assign n6721 =  ( n107 ) & ( n5194 )  ;
assign n6722 =  ( n107 ) & ( n5196 )  ;
assign n6723 =  ( n107 ) & ( n5198 )  ;
assign n6724 =  ( n107 ) & ( n5200 )  ;
assign n6725 =  ( n107 ) & ( n5202 )  ;
assign n6726 =  ( n107 ) & ( n5204 )  ;
assign n6727 =  ( n107 ) & ( n5206 )  ;
assign n6728 =  ( n107 ) & ( n5208 )  ;
assign n6729 =  ( n107 ) & ( n5210 )  ;
assign n6730 =  ( n107 ) & ( n5212 )  ;
assign n6731 =  ( n107 ) & ( n5214 )  ;
assign n6732 =  ( n107 ) & ( n5216 )  ;
assign n6733 =  ( n107 ) & ( n5218 )  ;
assign n6734 =  ( n108 ) & ( n5188 )  ;
assign n6735 =  ( n108 ) & ( n5190 )  ;
assign n6736 =  ( n108 ) & ( n5192 )  ;
assign n6737 =  ( n108 ) & ( n5194 )  ;
assign n6738 =  ( n108 ) & ( n5196 )  ;
assign n6739 =  ( n108 ) & ( n5198 )  ;
assign n6740 =  ( n108 ) & ( n5200 )  ;
assign n6741 =  ( n108 ) & ( n5202 )  ;
assign n6742 =  ( n108 ) & ( n5204 )  ;
assign n6743 =  ( n108 ) & ( n5206 )  ;
assign n6744 =  ( n108 ) & ( n5208 )  ;
assign n6745 =  ( n108 ) & ( n5210 )  ;
assign n6746 =  ( n108 ) & ( n5212 )  ;
assign n6747 =  ( n108 ) & ( n5214 )  ;
assign n6748 =  ( n108 ) & ( n5216 )  ;
assign n6749 =  ( n108 ) & ( n5218 )  ;
assign n6750 =  ( n6749 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n6751 =  ( n6748 ) ? ( VREG_0_1 ) : ( n6750 ) ;
assign n6752 =  ( n6747 ) ? ( VREG_0_2 ) : ( n6751 ) ;
assign n6753 =  ( n6746 ) ? ( VREG_0_3 ) : ( n6752 ) ;
assign n6754 =  ( n6745 ) ? ( VREG_0_4 ) : ( n6753 ) ;
assign n6755 =  ( n6744 ) ? ( VREG_0_5 ) : ( n6754 ) ;
assign n6756 =  ( n6743 ) ? ( VREG_0_6 ) : ( n6755 ) ;
assign n6757 =  ( n6742 ) ? ( VREG_0_7 ) : ( n6756 ) ;
assign n6758 =  ( n6741 ) ? ( VREG_0_8 ) : ( n6757 ) ;
assign n6759 =  ( n6740 ) ? ( VREG_0_9 ) : ( n6758 ) ;
assign n6760 =  ( n6739 ) ? ( VREG_0_10 ) : ( n6759 ) ;
assign n6761 =  ( n6738 ) ? ( VREG_0_11 ) : ( n6760 ) ;
assign n6762 =  ( n6737 ) ? ( VREG_0_12 ) : ( n6761 ) ;
assign n6763 =  ( n6736 ) ? ( VREG_0_13 ) : ( n6762 ) ;
assign n6764 =  ( n6735 ) ? ( VREG_0_14 ) : ( n6763 ) ;
assign n6765 =  ( n6734 ) ? ( VREG_0_15 ) : ( n6764 ) ;
assign n6766 =  ( n6733 ) ? ( VREG_1_0 ) : ( n6765 ) ;
assign n6767 =  ( n6732 ) ? ( VREG_1_1 ) : ( n6766 ) ;
assign n6768 =  ( n6731 ) ? ( VREG_1_2 ) : ( n6767 ) ;
assign n6769 =  ( n6730 ) ? ( VREG_1_3 ) : ( n6768 ) ;
assign n6770 =  ( n6729 ) ? ( VREG_1_4 ) : ( n6769 ) ;
assign n6771 =  ( n6728 ) ? ( VREG_1_5 ) : ( n6770 ) ;
assign n6772 =  ( n6727 ) ? ( VREG_1_6 ) : ( n6771 ) ;
assign n6773 =  ( n6726 ) ? ( VREG_1_7 ) : ( n6772 ) ;
assign n6774 =  ( n6725 ) ? ( VREG_1_8 ) : ( n6773 ) ;
assign n6775 =  ( n6724 ) ? ( VREG_1_9 ) : ( n6774 ) ;
assign n6776 =  ( n6723 ) ? ( VREG_1_10 ) : ( n6775 ) ;
assign n6777 =  ( n6722 ) ? ( VREG_1_11 ) : ( n6776 ) ;
assign n6778 =  ( n6721 ) ? ( VREG_1_12 ) : ( n6777 ) ;
assign n6779 =  ( n6720 ) ? ( VREG_1_13 ) : ( n6778 ) ;
assign n6780 =  ( n6719 ) ? ( VREG_1_14 ) : ( n6779 ) ;
assign n6781 =  ( n6718 ) ? ( VREG_1_15 ) : ( n6780 ) ;
assign n6782 =  ( n6717 ) ? ( VREG_2_0 ) : ( n6781 ) ;
assign n6783 =  ( n6716 ) ? ( VREG_2_1 ) : ( n6782 ) ;
assign n6784 =  ( n6715 ) ? ( VREG_2_2 ) : ( n6783 ) ;
assign n6785 =  ( n6714 ) ? ( VREG_2_3 ) : ( n6784 ) ;
assign n6786 =  ( n6713 ) ? ( VREG_2_4 ) : ( n6785 ) ;
assign n6787 =  ( n6712 ) ? ( VREG_2_5 ) : ( n6786 ) ;
assign n6788 =  ( n6711 ) ? ( VREG_2_6 ) : ( n6787 ) ;
assign n6789 =  ( n6710 ) ? ( VREG_2_7 ) : ( n6788 ) ;
assign n6790 =  ( n6709 ) ? ( VREG_2_8 ) : ( n6789 ) ;
assign n6791 =  ( n6708 ) ? ( VREG_2_9 ) : ( n6790 ) ;
assign n6792 =  ( n6707 ) ? ( VREG_2_10 ) : ( n6791 ) ;
assign n6793 =  ( n6706 ) ? ( VREG_2_11 ) : ( n6792 ) ;
assign n6794 =  ( n6705 ) ? ( VREG_2_12 ) : ( n6793 ) ;
assign n6795 =  ( n6704 ) ? ( VREG_2_13 ) : ( n6794 ) ;
assign n6796 =  ( n6703 ) ? ( VREG_2_14 ) : ( n6795 ) ;
assign n6797 =  ( n6702 ) ? ( VREG_2_15 ) : ( n6796 ) ;
assign n6798 =  ( n6701 ) ? ( VREG_3_0 ) : ( n6797 ) ;
assign n6799 =  ( n6700 ) ? ( VREG_3_1 ) : ( n6798 ) ;
assign n6800 =  ( n6699 ) ? ( VREG_3_2 ) : ( n6799 ) ;
assign n6801 =  ( n6698 ) ? ( VREG_3_3 ) : ( n6800 ) ;
assign n6802 =  ( n6697 ) ? ( VREG_3_4 ) : ( n6801 ) ;
assign n6803 =  ( n6696 ) ? ( VREG_3_5 ) : ( n6802 ) ;
assign n6804 =  ( n6695 ) ? ( VREG_3_6 ) : ( n6803 ) ;
assign n6805 =  ( n6694 ) ? ( VREG_3_7 ) : ( n6804 ) ;
assign n6806 =  ( n6693 ) ? ( VREG_3_8 ) : ( n6805 ) ;
assign n6807 =  ( n6692 ) ? ( VREG_3_9 ) : ( n6806 ) ;
assign n6808 =  ( n6691 ) ? ( VREG_3_10 ) : ( n6807 ) ;
assign n6809 =  ( n6690 ) ? ( VREG_3_11 ) : ( n6808 ) ;
assign n6810 =  ( n6689 ) ? ( VREG_3_12 ) : ( n6809 ) ;
assign n6811 =  ( n6688 ) ? ( VREG_3_13 ) : ( n6810 ) ;
assign n6812 =  ( n6687 ) ? ( VREG_3_14 ) : ( n6811 ) ;
assign n6813 =  ( n6686 ) ? ( VREG_3_15 ) : ( n6812 ) ;
assign n6814 =  ( n6685 ) ? ( VREG_4_0 ) : ( n6813 ) ;
assign n6815 =  ( n6684 ) ? ( VREG_4_1 ) : ( n6814 ) ;
assign n6816 =  ( n6683 ) ? ( VREG_4_2 ) : ( n6815 ) ;
assign n6817 =  ( n6682 ) ? ( VREG_4_3 ) : ( n6816 ) ;
assign n6818 =  ( n6681 ) ? ( VREG_4_4 ) : ( n6817 ) ;
assign n6819 =  ( n6680 ) ? ( VREG_4_5 ) : ( n6818 ) ;
assign n6820 =  ( n6679 ) ? ( VREG_4_6 ) : ( n6819 ) ;
assign n6821 =  ( n6678 ) ? ( VREG_4_7 ) : ( n6820 ) ;
assign n6822 =  ( n6677 ) ? ( VREG_4_8 ) : ( n6821 ) ;
assign n6823 =  ( n6676 ) ? ( VREG_4_9 ) : ( n6822 ) ;
assign n6824 =  ( n6675 ) ? ( VREG_4_10 ) : ( n6823 ) ;
assign n6825 =  ( n6674 ) ? ( VREG_4_11 ) : ( n6824 ) ;
assign n6826 =  ( n6673 ) ? ( VREG_4_12 ) : ( n6825 ) ;
assign n6827 =  ( n6672 ) ? ( VREG_4_13 ) : ( n6826 ) ;
assign n6828 =  ( n6671 ) ? ( VREG_4_14 ) : ( n6827 ) ;
assign n6829 =  ( n6670 ) ? ( VREG_4_15 ) : ( n6828 ) ;
assign n6830 =  ( n6669 ) ? ( VREG_5_0 ) : ( n6829 ) ;
assign n6831 =  ( n6668 ) ? ( VREG_5_1 ) : ( n6830 ) ;
assign n6832 =  ( n6667 ) ? ( VREG_5_2 ) : ( n6831 ) ;
assign n6833 =  ( n6666 ) ? ( VREG_5_3 ) : ( n6832 ) ;
assign n6834 =  ( n6665 ) ? ( VREG_5_4 ) : ( n6833 ) ;
assign n6835 =  ( n6664 ) ? ( VREG_5_5 ) : ( n6834 ) ;
assign n6836 =  ( n6663 ) ? ( VREG_5_6 ) : ( n6835 ) ;
assign n6837 =  ( n6662 ) ? ( VREG_5_7 ) : ( n6836 ) ;
assign n6838 =  ( n6661 ) ? ( VREG_5_8 ) : ( n6837 ) ;
assign n6839 =  ( n6660 ) ? ( VREG_5_9 ) : ( n6838 ) ;
assign n6840 =  ( n6659 ) ? ( VREG_5_10 ) : ( n6839 ) ;
assign n6841 =  ( n6658 ) ? ( VREG_5_11 ) : ( n6840 ) ;
assign n6842 =  ( n6657 ) ? ( VREG_5_12 ) : ( n6841 ) ;
assign n6843 =  ( n6656 ) ? ( VREG_5_13 ) : ( n6842 ) ;
assign n6844 =  ( n6655 ) ? ( VREG_5_14 ) : ( n6843 ) ;
assign n6845 =  ( n6654 ) ? ( VREG_5_15 ) : ( n6844 ) ;
assign n6846 =  ( n6653 ) ? ( VREG_6_0 ) : ( n6845 ) ;
assign n6847 =  ( n6652 ) ? ( VREG_6_1 ) : ( n6846 ) ;
assign n6848 =  ( n6651 ) ? ( VREG_6_2 ) : ( n6847 ) ;
assign n6849 =  ( n6650 ) ? ( VREG_6_3 ) : ( n6848 ) ;
assign n6850 =  ( n6649 ) ? ( VREG_6_4 ) : ( n6849 ) ;
assign n6851 =  ( n6648 ) ? ( VREG_6_5 ) : ( n6850 ) ;
assign n6852 =  ( n6647 ) ? ( VREG_6_6 ) : ( n6851 ) ;
assign n6853 =  ( n6646 ) ? ( VREG_6_7 ) : ( n6852 ) ;
assign n6854 =  ( n6645 ) ? ( VREG_6_8 ) : ( n6853 ) ;
assign n6855 =  ( n6644 ) ? ( VREG_6_9 ) : ( n6854 ) ;
assign n6856 =  ( n6643 ) ? ( VREG_6_10 ) : ( n6855 ) ;
assign n6857 =  ( n6642 ) ? ( VREG_6_11 ) : ( n6856 ) ;
assign n6858 =  ( n6641 ) ? ( VREG_6_12 ) : ( n6857 ) ;
assign n6859 =  ( n6640 ) ? ( VREG_6_13 ) : ( n6858 ) ;
assign n6860 =  ( n6639 ) ? ( VREG_6_14 ) : ( n6859 ) ;
assign n6861 =  ( n6638 ) ? ( VREG_6_15 ) : ( n6860 ) ;
assign n6862 =  ( n6637 ) ? ( VREG_7_0 ) : ( n6861 ) ;
assign n6863 =  ( n6636 ) ? ( VREG_7_1 ) : ( n6862 ) ;
assign n6864 =  ( n6635 ) ? ( VREG_7_2 ) : ( n6863 ) ;
assign n6865 =  ( n6634 ) ? ( VREG_7_3 ) : ( n6864 ) ;
assign n6866 =  ( n6633 ) ? ( VREG_7_4 ) : ( n6865 ) ;
assign n6867 =  ( n6632 ) ? ( VREG_7_5 ) : ( n6866 ) ;
assign n6868 =  ( n6631 ) ? ( VREG_7_6 ) : ( n6867 ) ;
assign n6869 =  ( n6630 ) ? ( VREG_7_7 ) : ( n6868 ) ;
assign n6870 =  ( n6629 ) ? ( VREG_7_8 ) : ( n6869 ) ;
assign n6871 =  ( n6628 ) ? ( VREG_7_9 ) : ( n6870 ) ;
assign n6872 =  ( n6627 ) ? ( VREG_7_10 ) : ( n6871 ) ;
assign n6873 =  ( n6626 ) ? ( VREG_7_11 ) : ( n6872 ) ;
assign n6874 =  ( n6625 ) ? ( VREG_7_12 ) : ( n6873 ) ;
assign n6875 =  ( n6624 ) ? ( VREG_7_13 ) : ( n6874 ) ;
assign n6876 =  ( n6623 ) ? ( VREG_7_14 ) : ( n6875 ) ;
assign n6877 =  ( n6622 ) ? ( VREG_7_15 ) : ( n6876 ) ;
assign n6878 =  ( n6621 ) ? ( VREG_8_0 ) : ( n6877 ) ;
assign n6879 =  ( n6620 ) ? ( VREG_8_1 ) : ( n6878 ) ;
assign n6880 =  ( n6619 ) ? ( VREG_8_2 ) : ( n6879 ) ;
assign n6881 =  ( n6618 ) ? ( VREG_8_3 ) : ( n6880 ) ;
assign n6882 =  ( n6617 ) ? ( VREG_8_4 ) : ( n6881 ) ;
assign n6883 =  ( n6616 ) ? ( VREG_8_5 ) : ( n6882 ) ;
assign n6884 =  ( n6615 ) ? ( VREG_8_6 ) : ( n6883 ) ;
assign n6885 =  ( n6614 ) ? ( VREG_8_7 ) : ( n6884 ) ;
assign n6886 =  ( n6613 ) ? ( VREG_8_8 ) : ( n6885 ) ;
assign n6887 =  ( n6612 ) ? ( VREG_8_9 ) : ( n6886 ) ;
assign n6888 =  ( n6611 ) ? ( VREG_8_10 ) : ( n6887 ) ;
assign n6889 =  ( n6610 ) ? ( VREG_8_11 ) : ( n6888 ) ;
assign n6890 =  ( n6609 ) ? ( VREG_8_12 ) : ( n6889 ) ;
assign n6891 =  ( n6608 ) ? ( VREG_8_13 ) : ( n6890 ) ;
assign n6892 =  ( n6607 ) ? ( VREG_8_14 ) : ( n6891 ) ;
assign n6893 =  ( n6606 ) ? ( VREG_8_15 ) : ( n6892 ) ;
assign n6894 =  ( n6605 ) ? ( VREG_9_0 ) : ( n6893 ) ;
assign n6895 =  ( n6604 ) ? ( VREG_9_1 ) : ( n6894 ) ;
assign n6896 =  ( n6603 ) ? ( VREG_9_2 ) : ( n6895 ) ;
assign n6897 =  ( n6602 ) ? ( VREG_9_3 ) : ( n6896 ) ;
assign n6898 =  ( n6601 ) ? ( VREG_9_4 ) : ( n6897 ) ;
assign n6899 =  ( n6600 ) ? ( VREG_9_5 ) : ( n6898 ) ;
assign n6900 =  ( n6599 ) ? ( VREG_9_6 ) : ( n6899 ) ;
assign n6901 =  ( n6598 ) ? ( VREG_9_7 ) : ( n6900 ) ;
assign n6902 =  ( n6597 ) ? ( VREG_9_8 ) : ( n6901 ) ;
assign n6903 =  ( n6596 ) ? ( VREG_9_9 ) : ( n6902 ) ;
assign n6904 =  ( n6595 ) ? ( VREG_9_10 ) : ( n6903 ) ;
assign n6905 =  ( n6594 ) ? ( VREG_9_11 ) : ( n6904 ) ;
assign n6906 =  ( n6593 ) ? ( VREG_9_12 ) : ( n6905 ) ;
assign n6907 =  ( n6592 ) ? ( VREG_9_13 ) : ( n6906 ) ;
assign n6908 =  ( n6591 ) ? ( VREG_9_14 ) : ( n6907 ) ;
assign n6909 =  ( n6590 ) ? ( VREG_9_15 ) : ( n6908 ) ;
assign n6910 =  ( n6589 ) ? ( VREG_10_0 ) : ( n6909 ) ;
assign n6911 =  ( n6588 ) ? ( VREG_10_1 ) : ( n6910 ) ;
assign n6912 =  ( n6587 ) ? ( VREG_10_2 ) : ( n6911 ) ;
assign n6913 =  ( n6586 ) ? ( VREG_10_3 ) : ( n6912 ) ;
assign n6914 =  ( n6585 ) ? ( VREG_10_4 ) : ( n6913 ) ;
assign n6915 =  ( n6584 ) ? ( VREG_10_5 ) : ( n6914 ) ;
assign n6916 =  ( n6583 ) ? ( VREG_10_6 ) : ( n6915 ) ;
assign n6917 =  ( n6582 ) ? ( VREG_10_7 ) : ( n6916 ) ;
assign n6918 =  ( n6581 ) ? ( VREG_10_8 ) : ( n6917 ) ;
assign n6919 =  ( n6580 ) ? ( VREG_10_9 ) : ( n6918 ) ;
assign n6920 =  ( n6579 ) ? ( VREG_10_10 ) : ( n6919 ) ;
assign n6921 =  ( n6578 ) ? ( VREG_10_11 ) : ( n6920 ) ;
assign n6922 =  ( n6577 ) ? ( VREG_10_12 ) : ( n6921 ) ;
assign n6923 =  ( n6576 ) ? ( VREG_10_13 ) : ( n6922 ) ;
assign n6924 =  ( n6575 ) ? ( VREG_10_14 ) : ( n6923 ) ;
assign n6925 =  ( n6574 ) ? ( VREG_10_15 ) : ( n6924 ) ;
assign n6926 =  ( n6573 ) ? ( VREG_11_0 ) : ( n6925 ) ;
assign n6927 =  ( n6572 ) ? ( VREG_11_1 ) : ( n6926 ) ;
assign n6928 =  ( n6571 ) ? ( VREG_11_2 ) : ( n6927 ) ;
assign n6929 =  ( n6570 ) ? ( VREG_11_3 ) : ( n6928 ) ;
assign n6930 =  ( n6569 ) ? ( VREG_11_4 ) : ( n6929 ) ;
assign n6931 =  ( n6568 ) ? ( VREG_11_5 ) : ( n6930 ) ;
assign n6932 =  ( n6567 ) ? ( VREG_11_6 ) : ( n6931 ) ;
assign n6933 =  ( n6566 ) ? ( VREG_11_7 ) : ( n6932 ) ;
assign n6934 =  ( n6565 ) ? ( VREG_11_8 ) : ( n6933 ) ;
assign n6935 =  ( n6564 ) ? ( VREG_11_9 ) : ( n6934 ) ;
assign n6936 =  ( n6563 ) ? ( VREG_11_10 ) : ( n6935 ) ;
assign n6937 =  ( n6562 ) ? ( VREG_11_11 ) : ( n6936 ) ;
assign n6938 =  ( n6561 ) ? ( VREG_11_12 ) : ( n6937 ) ;
assign n6939 =  ( n6560 ) ? ( VREG_11_13 ) : ( n6938 ) ;
assign n6940 =  ( n6559 ) ? ( VREG_11_14 ) : ( n6939 ) ;
assign n6941 =  ( n6558 ) ? ( VREG_11_15 ) : ( n6940 ) ;
assign n6942 =  ( n6557 ) ? ( VREG_12_0 ) : ( n6941 ) ;
assign n6943 =  ( n6556 ) ? ( VREG_12_1 ) : ( n6942 ) ;
assign n6944 =  ( n6555 ) ? ( VREG_12_2 ) : ( n6943 ) ;
assign n6945 =  ( n6554 ) ? ( VREG_12_3 ) : ( n6944 ) ;
assign n6946 =  ( n6553 ) ? ( VREG_12_4 ) : ( n6945 ) ;
assign n6947 =  ( n6552 ) ? ( VREG_12_5 ) : ( n6946 ) ;
assign n6948 =  ( n6551 ) ? ( VREG_12_6 ) : ( n6947 ) ;
assign n6949 =  ( n6550 ) ? ( VREG_12_7 ) : ( n6948 ) ;
assign n6950 =  ( n6549 ) ? ( VREG_12_8 ) : ( n6949 ) ;
assign n6951 =  ( n6548 ) ? ( VREG_12_9 ) : ( n6950 ) ;
assign n6952 =  ( n6547 ) ? ( VREG_12_10 ) : ( n6951 ) ;
assign n6953 =  ( n6546 ) ? ( VREG_12_11 ) : ( n6952 ) ;
assign n6954 =  ( n6545 ) ? ( VREG_12_12 ) : ( n6953 ) ;
assign n6955 =  ( n6544 ) ? ( VREG_12_13 ) : ( n6954 ) ;
assign n6956 =  ( n6543 ) ? ( VREG_12_14 ) : ( n6955 ) ;
assign n6957 =  ( n6542 ) ? ( VREG_12_15 ) : ( n6956 ) ;
assign n6958 =  ( n6541 ) ? ( VREG_13_0 ) : ( n6957 ) ;
assign n6959 =  ( n6540 ) ? ( VREG_13_1 ) : ( n6958 ) ;
assign n6960 =  ( n6539 ) ? ( VREG_13_2 ) : ( n6959 ) ;
assign n6961 =  ( n6538 ) ? ( VREG_13_3 ) : ( n6960 ) ;
assign n6962 =  ( n6537 ) ? ( VREG_13_4 ) : ( n6961 ) ;
assign n6963 =  ( n6536 ) ? ( VREG_13_5 ) : ( n6962 ) ;
assign n6964 =  ( n6535 ) ? ( VREG_13_6 ) : ( n6963 ) ;
assign n6965 =  ( n6534 ) ? ( VREG_13_7 ) : ( n6964 ) ;
assign n6966 =  ( n6533 ) ? ( VREG_13_8 ) : ( n6965 ) ;
assign n6967 =  ( n6532 ) ? ( VREG_13_9 ) : ( n6966 ) ;
assign n6968 =  ( n6531 ) ? ( VREG_13_10 ) : ( n6967 ) ;
assign n6969 =  ( n6530 ) ? ( VREG_13_11 ) : ( n6968 ) ;
assign n6970 =  ( n6529 ) ? ( VREG_13_12 ) : ( n6969 ) ;
assign n6971 =  ( n6528 ) ? ( VREG_13_13 ) : ( n6970 ) ;
assign n6972 =  ( n6527 ) ? ( VREG_13_14 ) : ( n6971 ) ;
assign n6973 =  ( n6526 ) ? ( VREG_13_15 ) : ( n6972 ) ;
assign n6974 =  ( n6525 ) ? ( VREG_14_0 ) : ( n6973 ) ;
assign n6975 =  ( n6524 ) ? ( VREG_14_1 ) : ( n6974 ) ;
assign n6976 =  ( n6523 ) ? ( VREG_14_2 ) : ( n6975 ) ;
assign n6977 =  ( n6522 ) ? ( VREG_14_3 ) : ( n6976 ) ;
assign n6978 =  ( n6521 ) ? ( VREG_14_4 ) : ( n6977 ) ;
assign n6979 =  ( n6520 ) ? ( VREG_14_5 ) : ( n6978 ) ;
assign n6980 =  ( n6519 ) ? ( VREG_14_6 ) : ( n6979 ) ;
assign n6981 =  ( n6518 ) ? ( VREG_14_7 ) : ( n6980 ) ;
assign n6982 =  ( n6517 ) ? ( VREG_14_8 ) : ( n6981 ) ;
assign n6983 =  ( n6516 ) ? ( VREG_14_9 ) : ( n6982 ) ;
assign n6984 =  ( n6515 ) ? ( VREG_14_10 ) : ( n6983 ) ;
assign n6985 =  ( n6514 ) ? ( VREG_14_11 ) : ( n6984 ) ;
assign n6986 =  ( n6513 ) ? ( VREG_14_12 ) : ( n6985 ) ;
assign n6987 =  ( n6512 ) ? ( VREG_14_13 ) : ( n6986 ) ;
assign n6988 =  ( n6511 ) ? ( VREG_14_14 ) : ( n6987 ) ;
assign n6989 =  ( n6510 ) ? ( VREG_14_15 ) : ( n6988 ) ;
assign n6990 =  ( n6509 ) ? ( VREG_15_0 ) : ( n6989 ) ;
assign n6991 =  ( n6508 ) ? ( VREG_15_1 ) : ( n6990 ) ;
assign n6992 =  ( n6507 ) ? ( VREG_15_2 ) : ( n6991 ) ;
assign n6993 =  ( n6506 ) ? ( VREG_15_3 ) : ( n6992 ) ;
assign n6994 =  ( n6505 ) ? ( VREG_15_4 ) : ( n6993 ) ;
assign n6995 =  ( n6504 ) ? ( VREG_15_5 ) : ( n6994 ) ;
assign n6996 =  ( n6503 ) ? ( VREG_15_6 ) : ( n6995 ) ;
assign n6997 =  ( n6502 ) ? ( VREG_15_7 ) : ( n6996 ) ;
assign n6998 =  ( n6501 ) ? ( VREG_15_8 ) : ( n6997 ) ;
assign n6999 =  ( n6500 ) ? ( VREG_15_9 ) : ( n6998 ) ;
assign n7000 =  ( n6499 ) ? ( VREG_15_10 ) : ( n6999 ) ;
assign n7001 =  ( n6498 ) ? ( VREG_15_11 ) : ( n7000 ) ;
assign n7002 =  ( n6497 ) ? ( VREG_15_12 ) : ( n7001 ) ;
assign n7003 =  ( n6496 ) ? ( VREG_15_13 ) : ( n7002 ) ;
assign n7004 =  ( n6495 ) ? ( VREG_15_14 ) : ( n7003 ) ;
assign n7005 =  ( n6494 ) ? ( VREG_15_15 ) : ( n7004 ) ;
assign n7006 =  ( n6493 ) ? ( VREG_16_0 ) : ( n7005 ) ;
assign n7007 =  ( n6492 ) ? ( VREG_16_1 ) : ( n7006 ) ;
assign n7008 =  ( n6491 ) ? ( VREG_16_2 ) : ( n7007 ) ;
assign n7009 =  ( n6490 ) ? ( VREG_16_3 ) : ( n7008 ) ;
assign n7010 =  ( n6489 ) ? ( VREG_16_4 ) : ( n7009 ) ;
assign n7011 =  ( n6488 ) ? ( VREG_16_5 ) : ( n7010 ) ;
assign n7012 =  ( n6487 ) ? ( VREG_16_6 ) : ( n7011 ) ;
assign n7013 =  ( n6486 ) ? ( VREG_16_7 ) : ( n7012 ) ;
assign n7014 =  ( n6485 ) ? ( VREG_16_8 ) : ( n7013 ) ;
assign n7015 =  ( n6484 ) ? ( VREG_16_9 ) : ( n7014 ) ;
assign n7016 =  ( n6483 ) ? ( VREG_16_10 ) : ( n7015 ) ;
assign n7017 =  ( n6482 ) ? ( VREG_16_11 ) : ( n7016 ) ;
assign n7018 =  ( n6481 ) ? ( VREG_16_12 ) : ( n7017 ) ;
assign n7019 =  ( n6480 ) ? ( VREG_16_13 ) : ( n7018 ) ;
assign n7020 =  ( n6479 ) ? ( VREG_16_14 ) : ( n7019 ) ;
assign n7021 =  ( n6478 ) ? ( VREG_16_15 ) : ( n7020 ) ;
assign n7022 =  ( n6477 ) ? ( VREG_17_0 ) : ( n7021 ) ;
assign n7023 =  ( n6476 ) ? ( VREG_17_1 ) : ( n7022 ) ;
assign n7024 =  ( n6475 ) ? ( VREG_17_2 ) : ( n7023 ) ;
assign n7025 =  ( n6474 ) ? ( VREG_17_3 ) : ( n7024 ) ;
assign n7026 =  ( n6473 ) ? ( VREG_17_4 ) : ( n7025 ) ;
assign n7027 =  ( n6472 ) ? ( VREG_17_5 ) : ( n7026 ) ;
assign n7028 =  ( n6471 ) ? ( VREG_17_6 ) : ( n7027 ) ;
assign n7029 =  ( n6470 ) ? ( VREG_17_7 ) : ( n7028 ) ;
assign n7030 =  ( n6469 ) ? ( VREG_17_8 ) : ( n7029 ) ;
assign n7031 =  ( n6468 ) ? ( VREG_17_9 ) : ( n7030 ) ;
assign n7032 =  ( n6467 ) ? ( VREG_17_10 ) : ( n7031 ) ;
assign n7033 =  ( n6466 ) ? ( VREG_17_11 ) : ( n7032 ) ;
assign n7034 =  ( n6465 ) ? ( VREG_17_12 ) : ( n7033 ) ;
assign n7035 =  ( n6464 ) ? ( VREG_17_13 ) : ( n7034 ) ;
assign n7036 =  ( n6463 ) ? ( VREG_17_14 ) : ( n7035 ) ;
assign n7037 =  ( n6462 ) ? ( VREG_17_15 ) : ( n7036 ) ;
assign n7038 =  ( n6461 ) ? ( VREG_18_0 ) : ( n7037 ) ;
assign n7039 =  ( n6460 ) ? ( VREG_18_1 ) : ( n7038 ) ;
assign n7040 =  ( n6459 ) ? ( VREG_18_2 ) : ( n7039 ) ;
assign n7041 =  ( n6458 ) ? ( VREG_18_3 ) : ( n7040 ) ;
assign n7042 =  ( n6457 ) ? ( VREG_18_4 ) : ( n7041 ) ;
assign n7043 =  ( n6456 ) ? ( VREG_18_5 ) : ( n7042 ) ;
assign n7044 =  ( n6455 ) ? ( VREG_18_6 ) : ( n7043 ) ;
assign n7045 =  ( n6454 ) ? ( VREG_18_7 ) : ( n7044 ) ;
assign n7046 =  ( n6453 ) ? ( VREG_18_8 ) : ( n7045 ) ;
assign n7047 =  ( n6452 ) ? ( VREG_18_9 ) : ( n7046 ) ;
assign n7048 =  ( n6451 ) ? ( VREG_18_10 ) : ( n7047 ) ;
assign n7049 =  ( n6450 ) ? ( VREG_18_11 ) : ( n7048 ) ;
assign n7050 =  ( n6449 ) ? ( VREG_18_12 ) : ( n7049 ) ;
assign n7051 =  ( n6448 ) ? ( VREG_18_13 ) : ( n7050 ) ;
assign n7052 =  ( n6447 ) ? ( VREG_18_14 ) : ( n7051 ) ;
assign n7053 =  ( n6446 ) ? ( VREG_18_15 ) : ( n7052 ) ;
assign n7054 =  ( n6445 ) ? ( VREG_19_0 ) : ( n7053 ) ;
assign n7055 =  ( n6444 ) ? ( VREG_19_1 ) : ( n7054 ) ;
assign n7056 =  ( n6443 ) ? ( VREG_19_2 ) : ( n7055 ) ;
assign n7057 =  ( n6442 ) ? ( VREG_19_3 ) : ( n7056 ) ;
assign n7058 =  ( n6441 ) ? ( VREG_19_4 ) : ( n7057 ) ;
assign n7059 =  ( n6440 ) ? ( VREG_19_5 ) : ( n7058 ) ;
assign n7060 =  ( n6439 ) ? ( VREG_19_6 ) : ( n7059 ) ;
assign n7061 =  ( n6438 ) ? ( VREG_19_7 ) : ( n7060 ) ;
assign n7062 =  ( n6437 ) ? ( VREG_19_8 ) : ( n7061 ) ;
assign n7063 =  ( n6436 ) ? ( VREG_19_9 ) : ( n7062 ) ;
assign n7064 =  ( n6435 ) ? ( VREG_19_10 ) : ( n7063 ) ;
assign n7065 =  ( n6434 ) ? ( VREG_19_11 ) : ( n7064 ) ;
assign n7066 =  ( n6433 ) ? ( VREG_19_12 ) : ( n7065 ) ;
assign n7067 =  ( n6432 ) ? ( VREG_19_13 ) : ( n7066 ) ;
assign n7068 =  ( n6431 ) ? ( VREG_19_14 ) : ( n7067 ) ;
assign n7069 =  ( n6430 ) ? ( VREG_19_15 ) : ( n7068 ) ;
assign n7070 =  ( n6429 ) ? ( VREG_20_0 ) : ( n7069 ) ;
assign n7071 =  ( n6428 ) ? ( VREG_20_1 ) : ( n7070 ) ;
assign n7072 =  ( n6427 ) ? ( VREG_20_2 ) : ( n7071 ) ;
assign n7073 =  ( n6426 ) ? ( VREG_20_3 ) : ( n7072 ) ;
assign n7074 =  ( n6425 ) ? ( VREG_20_4 ) : ( n7073 ) ;
assign n7075 =  ( n6424 ) ? ( VREG_20_5 ) : ( n7074 ) ;
assign n7076 =  ( n6423 ) ? ( VREG_20_6 ) : ( n7075 ) ;
assign n7077 =  ( n6422 ) ? ( VREG_20_7 ) : ( n7076 ) ;
assign n7078 =  ( n6421 ) ? ( VREG_20_8 ) : ( n7077 ) ;
assign n7079 =  ( n6420 ) ? ( VREG_20_9 ) : ( n7078 ) ;
assign n7080 =  ( n6419 ) ? ( VREG_20_10 ) : ( n7079 ) ;
assign n7081 =  ( n6418 ) ? ( VREG_20_11 ) : ( n7080 ) ;
assign n7082 =  ( n6417 ) ? ( VREG_20_12 ) : ( n7081 ) ;
assign n7083 =  ( n6416 ) ? ( VREG_20_13 ) : ( n7082 ) ;
assign n7084 =  ( n6415 ) ? ( VREG_20_14 ) : ( n7083 ) ;
assign n7085 =  ( n6414 ) ? ( VREG_20_15 ) : ( n7084 ) ;
assign n7086 =  ( n6413 ) ? ( VREG_21_0 ) : ( n7085 ) ;
assign n7087 =  ( n6412 ) ? ( VREG_21_1 ) : ( n7086 ) ;
assign n7088 =  ( n6411 ) ? ( VREG_21_2 ) : ( n7087 ) ;
assign n7089 =  ( n6410 ) ? ( VREG_21_3 ) : ( n7088 ) ;
assign n7090 =  ( n6409 ) ? ( VREG_21_4 ) : ( n7089 ) ;
assign n7091 =  ( n6408 ) ? ( VREG_21_5 ) : ( n7090 ) ;
assign n7092 =  ( n6407 ) ? ( VREG_21_6 ) : ( n7091 ) ;
assign n7093 =  ( n6406 ) ? ( VREG_21_7 ) : ( n7092 ) ;
assign n7094 =  ( n6405 ) ? ( VREG_21_8 ) : ( n7093 ) ;
assign n7095 =  ( n6404 ) ? ( VREG_21_9 ) : ( n7094 ) ;
assign n7096 =  ( n6403 ) ? ( VREG_21_10 ) : ( n7095 ) ;
assign n7097 =  ( n6402 ) ? ( VREG_21_11 ) : ( n7096 ) ;
assign n7098 =  ( n6401 ) ? ( VREG_21_12 ) : ( n7097 ) ;
assign n7099 =  ( n6400 ) ? ( VREG_21_13 ) : ( n7098 ) ;
assign n7100 =  ( n6399 ) ? ( VREG_21_14 ) : ( n7099 ) ;
assign n7101 =  ( n6398 ) ? ( VREG_21_15 ) : ( n7100 ) ;
assign n7102 =  ( n6397 ) ? ( VREG_22_0 ) : ( n7101 ) ;
assign n7103 =  ( n6396 ) ? ( VREG_22_1 ) : ( n7102 ) ;
assign n7104 =  ( n6395 ) ? ( VREG_22_2 ) : ( n7103 ) ;
assign n7105 =  ( n6394 ) ? ( VREG_22_3 ) : ( n7104 ) ;
assign n7106 =  ( n6393 ) ? ( VREG_22_4 ) : ( n7105 ) ;
assign n7107 =  ( n6392 ) ? ( VREG_22_5 ) : ( n7106 ) ;
assign n7108 =  ( n6391 ) ? ( VREG_22_6 ) : ( n7107 ) ;
assign n7109 =  ( n6390 ) ? ( VREG_22_7 ) : ( n7108 ) ;
assign n7110 =  ( n6389 ) ? ( VREG_22_8 ) : ( n7109 ) ;
assign n7111 =  ( n6388 ) ? ( VREG_22_9 ) : ( n7110 ) ;
assign n7112 =  ( n6387 ) ? ( VREG_22_10 ) : ( n7111 ) ;
assign n7113 =  ( n6386 ) ? ( VREG_22_11 ) : ( n7112 ) ;
assign n7114 =  ( n6385 ) ? ( VREG_22_12 ) : ( n7113 ) ;
assign n7115 =  ( n6384 ) ? ( VREG_22_13 ) : ( n7114 ) ;
assign n7116 =  ( n6383 ) ? ( VREG_22_14 ) : ( n7115 ) ;
assign n7117 =  ( n6382 ) ? ( VREG_22_15 ) : ( n7116 ) ;
assign n7118 =  ( n6381 ) ? ( VREG_23_0 ) : ( n7117 ) ;
assign n7119 =  ( n6380 ) ? ( VREG_23_1 ) : ( n7118 ) ;
assign n7120 =  ( n6379 ) ? ( VREG_23_2 ) : ( n7119 ) ;
assign n7121 =  ( n6378 ) ? ( VREG_23_3 ) : ( n7120 ) ;
assign n7122 =  ( n6377 ) ? ( VREG_23_4 ) : ( n7121 ) ;
assign n7123 =  ( n6376 ) ? ( VREG_23_5 ) : ( n7122 ) ;
assign n7124 =  ( n6375 ) ? ( VREG_23_6 ) : ( n7123 ) ;
assign n7125 =  ( n6374 ) ? ( VREG_23_7 ) : ( n7124 ) ;
assign n7126 =  ( n6373 ) ? ( VREG_23_8 ) : ( n7125 ) ;
assign n7127 =  ( n6372 ) ? ( VREG_23_9 ) : ( n7126 ) ;
assign n7128 =  ( n6371 ) ? ( VREG_23_10 ) : ( n7127 ) ;
assign n7129 =  ( n6370 ) ? ( VREG_23_11 ) : ( n7128 ) ;
assign n7130 =  ( n6369 ) ? ( VREG_23_12 ) : ( n7129 ) ;
assign n7131 =  ( n6368 ) ? ( VREG_23_13 ) : ( n7130 ) ;
assign n7132 =  ( n6367 ) ? ( VREG_23_14 ) : ( n7131 ) ;
assign n7133 =  ( n6366 ) ? ( VREG_23_15 ) : ( n7132 ) ;
assign n7134 =  ( n6365 ) ? ( VREG_24_0 ) : ( n7133 ) ;
assign n7135 =  ( n6364 ) ? ( VREG_24_1 ) : ( n7134 ) ;
assign n7136 =  ( n6363 ) ? ( VREG_24_2 ) : ( n7135 ) ;
assign n7137 =  ( n6362 ) ? ( VREG_24_3 ) : ( n7136 ) ;
assign n7138 =  ( n6361 ) ? ( VREG_24_4 ) : ( n7137 ) ;
assign n7139 =  ( n6360 ) ? ( VREG_24_5 ) : ( n7138 ) ;
assign n7140 =  ( n6359 ) ? ( VREG_24_6 ) : ( n7139 ) ;
assign n7141 =  ( n6358 ) ? ( VREG_24_7 ) : ( n7140 ) ;
assign n7142 =  ( n6357 ) ? ( VREG_24_8 ) : ( n7141 ) ;
assign n7143 =  ( n6356 ) ? ( VREG_24_9 ) : ( n7142 ) ;
assign n7144 =  ( n6355 ) ? ( VREG_24_10 ) : ( n7143 ) ;
assign n7145 =  ( n6354 ) ? ( VREG_24_11 ) : ( n7144 ) ;
assign n7146 =  ( n6353 ) ? ( VREG_24_12 ) : ( n7145 ) ;
assign n7147 =  ( n6352 ) ? ( VREG_24_13 ) : ( n7146 ) ;
assign n7148 =  ( n6351 ) ? ( VREG_24_14 ) : ( n7147 ) ;
assign n7149 =  ( n6350 ) ? ( VREG_24_15 ) : ( n7148 ) ;
assign n7150 =  ( n6349 ) ? ( VREG_25_0 ) : ( n7149 ) ;
assign n7151 =  ( n6348 ) ? ( VREG_25_1 ) : ( n7150 ) ;
assign n7152 =  ( n6347 ) ? ( VREG_25_2 ) : ( n7151 ) ;
assign n7153 =  ( n6346 ) ? ( VREG_25_3 ) : ( n7152 ) ;
assign n7154 =  ( n6345 ) ? ( VREG_25_4 ) : ( n7153 ) ;
assign n7155 =  ( n6344 ) ? ( VREG_25_5 ) : ( n7154 ) ;
assign n7156 =  ( n6343 ) ? ( VREG_25_6 ) : ( n7155 ) ;
assign n7157 =  ( n6342 ) ? ( VREG_25_7 ) : ( n7156 ) ;
assign n7158 =  ( n6341 ) ? ( VREG_25_8 ) : ( n7157 ) ;
assign n7159 =  ( n6340 ) ? ( VREG_25_9 ) : ( n7158 ) ;
assign n7160 =  ( n6339 ) ? ( VREG_25_10 ) : ( n7159 ) ;
assign n7161 =  ( n6338 ) ? ( VREG_25_11 ) : ( n7160 ) ;
assign n7162 =  ( n6337 ) ? ( VREG_25_12 ) : ( n7161 ) ;
assign n7163 =  ( n6336 ) ? ( VREG_25_13 ) : ( n7162 ) ;
assign n7164 =  ( n6335 ) ? ( VREG_25_14 ) : ( n7163 ) ;
assign n7165 =  ( n6334 ) ? ( VREG_25_15 ) : ( n7164 ) ;
assign n7166 =  ( n6333 ) ? ( VREG_26_0 ) : ( n7165 ) ;
assign n7167 =  ( n6332 ) ? ( VREG_26_1 ) : ( n7166 ) ;
assign n7168 =  ( n6331 ) ? ( VREG_26_2 ) : ( n7167 ) ;
assign n7169 =  ( n6330 ) ? ( VREG_26_3 ) : ( n7168 ) ;
assign n7170 =  ( n6329 ) ? ( VREG_26_4 ) : ( n7169 ) ;
assign n7171 =  ( n6328 ) ? ( VREG_26_5 ) : ( n7170 ) ;
assign n7172 =  ( n6327 ) ? ( VREG_26_6 ) : ( n7171 ) ;
assign n7173 =  ( n6326 ) ? ( VREG_26_7 ) : ( n7172 ) ;
assign n7174 =  ( n6325 ) ? ( VREG_26_8 ) : ( n7173 ) ;
assign n7175 =  ( n6324 ) ? ( VREG_26_9 ) : ( n7174 ) ;
assign n7176 =  ( n6323 ) ? ( VREG_26_10 ) : ( n7175 ) ;
assign n7177 =  ( n6322 ) ? ( VREG_26_11 ) : ( n7176 ) ;
assign n7178 =  ( n6321 ) ? ( VREG_26_12 ) : ( n7177 ) ;
assign n7179 =  ( n6320 ) ? ( VREG_26_13 ) : ( n7178 ) ;
assign n7180 =  ( n6319 ) ? ( VREG_26_14 ) : ( n7179 ) ;
assign n7181 =  ( n6318 ) ? ( VREG_26_15 ) : ( n7180 ) ;
assign n7182 =  ( n6317 ) ? ( VREG_27_0 ) : ( n7181 ) ;
assign n7183 =  ( n6316 ) ? ( VREG_27_1 ) : ( n7182 ) ;
assign n7184 =  ( n6315 ) ? ( VREG_27_2 ) : ( n7183 ) ;
assign n7185 =  ( n6314 ) ? ( VREG_27_3 ) : ( n7184 ) ;
assign n7186 =  ( n6313 ) ? ( VREG_27_4 ) : ( n7185 ) ;
assign n7187 =  ( n6312 ) ? ( VREG_27_5 ) : ( n7186 ) ;
assign n7188 =  ( n6311 ) ? ( VREG_27_6 ) : ( n7187 ) ;
assign n7189 =  ( n6310 ) ? ( VREG_27_7 ) : ( n7188 ) ;
assign n7190 =  ( n6309 ) ? ( VREG_27_8 ) : ( n7189 ) ;
assign n7191 =  ( n6308 ) ? ( VREG_27_9 ) : ( n7190 ) ;
assign n7192 =  ( n6307 ) ? ( VREG_27_10 ) : ( n7191 ) ;
assign n7193 =  ( n6306 ) ? ( VREG_27_11 ) : ( n7192 ) ;
assign n7194 =  ( n6305 ) ? ( VREG_27_12 ) : ( n7193 ) ;
assign n7195 =  ( n6304 ) ? ( VREG_27_13 ) : ( n7194 ) ;
assign n7196 =  ( n6303 ) ? ( VREG_27_14 ) : ( n7195 ) ;
assign n7197 =  ( n6302 ) ? ( VREG_27_15 ) : ( n7196 ) ;
assign n7198 =  ( n6301 ) ? ( VREG_28_0 ) : ( n7197 ) ;
assign n7199 =  ( n6300 ) ? ( VREG_28_1 ) : ( n7198 ) ;
assign n7200 =  ( n6299 ) ? ( VREG_28_2 ) : ( n7199 ) ;
assign n7201 =  ( n6298 ) ? ( VREG_28_3 ) : ( n7200 ) ;
assign n7202 =  ( n6297 ) ? ( VREG_28_4 ) : ( n7201 ) ;
assign n7203 =  ( n6296 ) ? ( VREG_28_5 ) : ( n7202 ) ;
assign n7204 =  ( n6295 ) ? ( VREG_28_6 ) : ( n7203 ) ;
assign n7205 =  ( n6294 ) ? ( VREG_28_7 ) : ( n7204 ) ;
assign n7206 =  ( n6293 ) ? ( VREG_28_8 ) : ( n7205 ) ;
assign n7207 =  ( n6292 ) ? ( VREG_28_9 ) : ( n7206 ) ;
assign n7208 =  ( n6291 ) ? ( VREG_28_10 ) : ( n7207 ) ;
assign n7209 =  ( n6290 ) ? ( VREG_28_11 ) : ( n7208 ) ;
assign n7210 =  ( n6289 ) ? ( VREG_28_12 ) : ( n7209 ) ;
assign n7211 =  ( n6288 ) ? ( VREG_28_13 ) : ( n7210 ) ;
assign n7212 =  ( n6287 ) ? ( VREG_28_14 ) : ( n7211 ) ;
assign n7213 =  ( n6286 ) ? ( VREG_28_15 ) : ( n7212 ) ;
assign n7214 =  ( n6285 ) ? ( VREG_29_0 ) : ( n7213 ) ;
assign n7215 =  ( n6284 ) ? ( VREG_29_1 ) : ( n7214 ) ;
assign n7216 =  ( n6283 ) ? ( VREG_29_2 ) : ( n7215 ) ;
assign n7217 =  ( n6282 ) ? ( VREG_29_3 ) : ( n7216 ) ;
assign n7218 =  ( n6281 ) ? ( VREG_29_4 ) : ( n7217 ) ;
assign n7219 =  ( n6280 ) ? ( VREG_29_5 ) : ( n7218 ) ;
assign n7220 =  ( n6279 ) ? ( VREG_29_6 ) : ( n7219 ) ;
assign n7221 =  ( n6278 ) ? ( VREG_29_7 ) : ( n7220 ) ;
assign n7222 =  ( n6277 ) ? ( VREG_29_8 ) : ( n7221 ) ;
assign n7223 =  ( n6276 ) ? ( VREG_29_9 ) : ( n7222 ) ;
assign n7224 =  ( n6275 ) ? ( VREG_29_10 ) : ( n7223 ) ;
assign n7225 =  ( n6274 ) ? ( VREG_29_11 ) : ( n7224 ) ;
assign n7226 =  ( n6273 ) ? ( VREG_29_12 ) : ( n7225 ) ;
assign n7227 =  ( n6272 ) ? ( VREG_29_13 ) : ( n7226 ) ;
assign n7228 =  ( n6271 ) ? ( VREG_29_14 ) : ( n7227 ) ;
assign n7229 =  ( n6270 ) ? ( VREG_29_15 ) : ( n7228 ) ;
assign n7230 =  ( n6269 ) ? ( VREG_30_0 ) : ( n7229 ) ;
assign n7231 =  ( n6268 ) ? ( VREG_30_1 ) : ( n7230 ) ;
assign n7232 =  ( n6267 ) ? ( VREG_30_2 ) : ( n7231 ) ;
assign n7233 =  ( n6266 ) ? ( VREG_30_3 ) : ( n7232 ) ;
assign n7234 =  ( n6265 ) ? ( VREG_30_4 ) : ( n7233 ) ;
assign n7235 =  ( n6264 ) ? ( VREG_30_5 ) : ( n7234 ) ;
assign n7236 =  ( n6263 ) ? ( VREG_30_6 ) : ( n7235 ) ;
assign n7237 =  ( n6262 ) ? ( VREG_30_7 ) : ( n7236 ) ;
assign n7238 =  ( n6261 ) ? ( VREG_30_8 ) : ( n7237 ) ;
assign n7239 =  ( n6260 ) ? ( VREG_30_9 ) : ( n7238 ) ;
assign n7240 =  ( n6259 ) ? ( VREG_30_10 ) : ( n7239 ) ;
assign n7241 =  ( n6258 ) ? ( VREG_30_11 ) : ( n7240 ) ;
assign n7242 =  ( n6257 ) ? ( VREG_30_12 ) : ( n7241 ) ;
assign n7243 =  ( n6256 ) ? ( VREG_30_13 ) : ( n7242 ) ;
assign n7244 =  ( n6255 ) ? ( VREG_30_14 ) : ( n7243 ) ;
assign n7245 =  ( n6254 ) ? ( VREG_30_15 ) : ( n7244 ) ;
assign n7246 =  ( n6253 ) ? ( VREG_31_0 ) : ( n7245 ) ;
assign n7247 =  ( n6252 ) ? ( VREG_31_1 ) : ( n7246 ) ;
assign n7248 =  ( n6251 ) ? ( VREG_31_2 ) : ( n7247 ) ;
assign n7249 =  ( n6250 ) ? ( VREG_31_3 ) : ( n7248 ) ;
assign n7250 =  ( n6249 ) ? ( VREG_31_4 ) : ( n7249 ) ;
assign n7251 =  ( n6248 ) ? ( VREG_31_5 ) : ( n7250 ) ;
assign n7252 =  ( n6247 ) ? ( VREG_31_6 ) : ( n7251 ) ;
assign n7253 =  ( n6246 ) ? ( VREG_31_7 ) : ( n7252 ) ;
assign n7254 =  ( n6245 ) ? ( VREG_31_8 ) : ( n7253 ) ;
assign n7255 =  ( n6244 ) ? ( VREG_31_9 ) : ( n7254 ) ;
assign n7256 =  ( n6243 ) ? ( VREG_31_10 ) : ( n7255 ) ;
assign n7257 =  ( n6242 ) ? ( VREG_31_11 ) : ( n7256 ) ;
assign n7258 =  ( n6241 ) ? ( VREG_31_12 ) : ( n7257 ) ;
assign n7259 =  ( n6240 ) ? ( VREG_31_13 ) : ( n7258 ) ;
assign n7260 =  ( n6239 ) ? ( VREG_31_14 ) : ( n7259 ) ;
assign n7261 =  ( n6238 ) ? ( VREG_31_15 ) : ( n7260 ) ;
assign n7262 =  ( n6227 ) + ( n7261 )  ;
assign n7263 =  ( n6227 ) - ( n7261 )  ;
assign n7264 =  ( n6227 ) & ( n7261 )  ;
assign n7265 =  ( n6227 ) | ( n7261 )  ;
assign n7266 =  ( ( n6227 ) * ( n7261 ))  ;
assign n7267 =  ( n148 ) ? ( n7266 ) : ( VREG_0_10 ) ;
assign n7268 =  ( n146 ) ? ( n7265 ) : ( n7267 ) ;
assign n7269 =  ( n144 ) ? ( n7264 ) : ( n7268 ) ;
assign n7270 =  ( n142 ) ? ( n7263 ) : ( n7269 ) ;
assign n7271 =  ( n10 ) ? ( n7262 ) : ( n7270 ) ;
assign n7272 = n3030[10:10] ;
assign n7273 =  ( n7272 ) == ( 1'd0 )  ;
assign n7274 =  ( n7273 ) ? ( VREG_0_10 ) : ( n6237 ) ;
assign n7275 =  ( n7273 ) ? ( VREG_0_10 ) : ( n7271 ) ;
assign n7276 =  ( n3034 ) ? ( n7275 ) : ( VREG_0_10 ) ;
assign n7277 =  ( n2965 ) ? ( n7274 ) : ( n7276 ) ;
assign n7278 =  ( n1930 ) ? ( n7271 ) : ( n7277 ) ;
assign n7279 =  ( n879 ) ? ( n6237 ) : ( n7278 ) ;
assign n7280 =  ( n6227 ) + ( n164 )  ;
assign n7281 =  ( n6227 ) - ( n164 )  ;
assign n7282 =  ( n6227 ) & ( n164 )  ;
assign n7283 =  ( n6227 ) | ( n164 )  ;
assign n7284 =  ( ( n6227 ) * ( n164 ))  ;
assign n7285 =  ( n172 ) ? ( n7284 ) : ( VREG_0_10 ) ;
assign n7286 =  ( n170 ) ? ( n7283 ) : ( n7285 ) ;
assign n7287 =  ( n168 ) ? ( n7282 ) : ( n7286 ) ;
assign n7288 =  ( n166 ) ? ( n7281 ) : ( n7287 ) ;
assign n7289 =  ( n162 ) ? ( n7280 ) : ( n7288 ) ;
assign n7290 =  ( n6227 ) + ( n180 )  ;
assign n7291 =  ( n6227 ) - ( n180 )  ;
assign n7292 =  ( n6227 ) & ( n180 )  ;
assign n7293 =  ( n6227 ) | ( n180 )  ;
assign n7294 =  ( ( n6227 ) * ( n180 ))  ;
assign n7295 =  ( n172 ) ? ( n7294 ) : ( VREG_0_10 ) ;
assign n7296 =  ( n170 ) ? ( n7293 ) : ( n7295 ) ;
assign n7297 =  ( n168 ) ? ( n7292 ) : ( n7296 ) ;
assign n7298 =  ( n166 ) ? ( n7291 ) : ( n7297 ) ;
assign n7299 =  ( n162 ) ? ( n7290 ) : ( n7298 ) ;
assign n7300 =  ( n7273 ) ? ( VREG_0_10 ) : ( n7299 ) ;
assign n7301 =  ( n3051 ) ? ( n7300 ) : ( VREG_0_10 ) ;
assign n7302 =  ( n3040 ) ? ( n7289 ) : ( n7301 ) ;
assign n7303 =  ( n192 ) ? ( VREG_0_10 ) : ( VREG_0_10 ) ;
assign n7304 =  ( n157 ) ? ( n7302 ) : ( n7303 ) ;
assign n7305 =  ( n6 ) ? ( n7279 ) : ( n7304 ) ;
assign n7306 =  ( n4 ) ? ( n7305 ) : ( VREG_0_10 ) ;
assign n7307 =  ( 32'd11 ) == ( 32'd15 )  ;
assign n7308 =  ( n12 ) & ( n7307 )  ;
assign n7309 =  ( 32'd11 ) == ( 32'd14 )  ;
assign n7310 =  ( n12 ) & ( n7309 )  ;
assign n7311 =  ( 32'd11 ) == ( 32'd13 )  ;
assign n7312 =  ( n12 ) & ( n7311 )  ;
assign n7313 =  ( 32'd11 ) == ( 32'd12 )  ;
assign n7314 =  ( n12 ) & ( n7313 )  ;
assign n7315 =  ( 32'd11 ) == ( 32'd11 )  ;
assign n7316 =  ( n12 ) & ( n7315 )  ;
assign n7317 =  ( 32'd11 ) == ( 32'd10 )  ;
assign n7318 =  ( n12 ) & ( n7317 )  ;
assign n7319 =  ( 32'd11 ) == ( 32'd9 )  ;
assign n7320 =  ( n12 ) & ( n7319 )  ;
assign n7321 =  ( 32'd11 ) == ( 32'd8 )  ;
assign n7322 =  ( n12 ) & ( n7321 )  ;
assign n7323 =  ( 32'd11 ) == ( 32'd7 )  ;
assign n7324 =  ( n12 ) & ( n7323 )  ;
assign n7325 =  ( 32'd11 ) == ( 32'd6 )  ;
assign n7326 =  ( n12 ) & ( n7325 )  ;
assign n7327 =  ( 32'd11 ) == ( 32'd5 )  ;
assign n7328 =  ( n12 ) & ( n7327 )  ;
assign n7329 =  ( 32'd11 ) == ( 32'd4 )  ;
assign n7330 =  ( n12 ) & ( n7329 )  ;
assign n7331 =  ( 32'd11 ) == ( 32'd3 )  ;
assign n7332 =  ( n12 ) & ( n7331 )  ;
assign n7333 =  ( 32'd11 ) == ( 32'd2 )  ;
assign n7334 =  ( n12 ) & ( n7333 )  ;
assign n7335 =  ( 32'd11 ) == ( 32'd1 )  ;
assign n7336 =  ( n12 ) & ( n7335 )  ;
assign n7337 =  ( 32'd11 ) == ( 32'd0 )  ;
assign n7338 =  ( n12 ) & ( n7337 )  ;
assign n7339 =  ( n13 ) & ( n7307 )  ;
assign n7340 =  ( n13 ) & ( n7309 )  ;
assign n7341 =  ( n13 ) & ( n7311 )  ;
assign n7342 =  ( n13 ) & ( n7313 )  ;
assign n7343 =  ( n13 ) & ( n7315 )  ;
assign n7344 =  ( n13 ) & ( n7317 )  ;
assign n7345 =  ( n13 ) & ( n7319 )  ;
assign n7346 =  ( n13 ) & ( n7321 )  ;
assign n7347 =  ( n13 ) & ( n7323 )  ;
assign n7348 =  ( n13 ) & ( n7325 )  ;
assign n7349 =  ( n13 ) & ( n7327 )  ;
assign n7350 =  ( n13 ) & ( n7329 )  ;
assign n7351 =  ( n13 ) & ( n7331 )  ;
assign n7352 =  ( n13 ) & ( n7333 )  ;
assign n7353 =  ( n13 ) & ( n7335 )  ;
assign n7354 =  ( n13 ) & ( n7337 )  ;
assign n7355 =  ( n14 ) & ( n7307 )  ;
assign n7356 =  ( n14 ) & ( n7309 )  ;
assign n7357 =  ( n14 ) & ( n7311 )  ;
assign n7358 =  ( n14 ) & ( n7313 )  ;
assign n7359 =  ( n14 ) & ( n7315 )  ;
assign n7360 =  ( n14 ) & ( n7317 )  ;
assign n7361 =  ( n14 ) & ( n7319 )  ;
assign n7362 =  ( n14 ) & ( n7321 )  ;
assign n7363 =  ( n14 ) & ( n7323 )  ;
assign n7364 =  ( n14 ) & ( n7325 )  ;
assign n7365 =  ( n14 ) & ( n7327 )  ;
assign n7366 =  ( n14 ) & ( n7329 )  ;
assign n7367 =  ( n14 ) & ( n7331 )  ;
assign n7368 =  ( n14 ) & ( n7333 )  ;
assign n7369 =  ( n14 ) & ( n7335 )  ;
assign n7370 =  ( n14 ) & ( n7337 )  ;
assign n7371 =  ( n15 ) & ( n7307 )  ;
assign n7372 =  ( n15 ) & ( n7309 )  ;
assign n7373 =  ( n15 ) & ( n7311 )  ;
assign n7374 =  ( n15 ) & ( n7313 )  ;
assign n7375 =  ( n15 ) & ( n7315 )  ;
assign n7376 =  ( n15 ) & ( n7317 )  ;
assign n7377 =  ( n15 ) & ( n7319 )  ;
assign n7378 =  ( n15 ) & ( n7321 )  ;
assign n7379 =  ( n15 ) & ( n7323 )  ;
assign n7380 =  ( n15 ) & ( n7325 )  ;
assign n7381 =  ( n15 ) & ( n7327 )  ;
assign n7382 =  ( n15 ) & ( n7329 )  ;
assign n7383 =  ( n15 ) & ( n7331 )  ;
assign n7384 =  ( n15 ) & ( n7333 )  ;
assign n7385 =  ( n15 ) & ( n7335 )  ;
assign n7386 =  ( n15 ) & ( n7337 )  ;
assign n7387 =  ( n16 ) & ( n7307 )  ;
assign n7388 =  ( n16 ) & ( n7309 )  ;
assign n7389 =  ( n16 ) & ( n7311 )  ;
assign n7390 =  ( n16 ) & ( n7313 )  ;
assign n7391 =  ( n16 ) & ( n7315 )  ;
assign n7392 =  ( n16 ) & ( n7317 )  ;
assign n7393 =  ( n16 ) & ( n7319 )  ;
assign n7394 =  ( n16 ) & ( n7321 )  ;
assign n7395 =  ( n16 ) & ( n7323 )  ;
assign n7396 =  ( n16 ) & ( n7325 )  ;
assign n7397 =  ( n16 ) & ( n7327 )  ;
assign n7398 =  ( n16 ) & ( n7329 )  ;
assign n7399 =  ( n16 ) & ( n7331 )  ;
assign n7400 =  ( n16 ) & ( n7333 )  ;
assign n7401 =  ( n16 ) & ( n7335 )  ;
assign n7402 =  ( n16 ) & ( n7337 )  ;
assign n7403 =  ( n17 ) & ( n7307 )  ;
assign n7404 =  ( n17 ) & ( n7309 )  ;
assign n7405 =  ( n17 ) & ( n7311 )  ;
assign n7406 =  ( n17 ) & ( n7313 )  ;
assign n7407 =  ( n17 ) & ( n7315 )  ;
assign n7408 =  ( n17 ) & ( n7317 )  ;
assign n7409 =  ( n17 ) & ( n7319 )  ;
assign n7410 =  ( n17 ) & ( n7321 )  ;
assign n7411 =  ( n17 ) & ( n7323 )  ;
assign n7412 =  ( n17 ) & ( n7325 )  ;
assign n7413 =  ( n17 ) & ( n7327 )  ;
assign n7414 =  ( n17 ) & ( n7329 )  ;
assign n7415 =  ( n17 ) & ( n7331 )  ;
assign n7416 =  ( n17 ) & ( n7333 )  ;
assign n7417 =  ( n17 ) & ( n7335 )  ;
assign n7418 =  ( n17 ) & ( n7337 )  ;
assign n7419 =  ( n18 ) & ( n7307 )  ;
assign n7420 =  ( n18 ) & ( n7309 )  ;
assign n7421 =  ( n18 ) & ( n7311 )  ;
assign n7422 =  ( n18 ) & ( n7313 )  ;
assign n7423 =  ( n18 ) & ( n7315 )  ;
assign n7424 =  ( n18 ) & ( n7317 )  ;
assign n7425 =  ( n18 ) & ( n7319 )  ;
assign n7426 =  ( n18 ) & ( n7321 )  ;
assign n7427 =  ( n18 ) & ( n7323 )  ;
assign n7428 =  ( n18 ) & ( n7325 )  ;
assign n7429 =  ( n18 ) & ( n7327 )  ;
assign n7430 =  ( n18 ) & ( n7329 )  ;
assign n7431 =  ( n18 ) & ( n7331 )  ;
assign n7432 =  ( n18 ) & ( n7333 )  ;
assign n7433 =  ( n18 ) & ( n7335 )  ;
assign n7434 =  ( n18 ) & ( n7337 )  ;
assign n7435 =  ( n19 ) & ( n7307 )  ;
assign n7436 =  ( n19 ) & ( n7309 )  ;
assign n7437 =  ( n19 ) & ( n7311 )  ;
assign n7438 =  ( n19 ) & ( n7313 )  ;
assign n7439 =  ( n19 ) & ( n7315 )  ;
assign n7440 =  ( n19 ) & ( n7317 )  ;
assign n7441 =  ( n19 ) & ( n7319 )  ;
assign n7442 =  ( n19 ) & ( n7321 )  ;
assign n7443 =  ( n19 ) & ( n7323 )  ;
assign n7444 =  ( n19 ) & ( n7325 )  ;
assign n7445 =  ( n19 ) & ( n7327 )  ;
assign n7446 =  ( n19 ) & ( n7329 )  ;
assign n7447 =  ( n19 ) & ( n7331 )  ;
assign n7448 =  ( n19 ) & ( n7333 )  ;
assign n7449 =  ( n19 ) & ( n7335 )  ;
assign n7450 =  ( n19 ) & ( n7337 )  ;
assign n7451 =  ( n20 ) & ( n7307 )  ;
assign n7452 =  ( n20 ) & ( n7309 )  ;
assign n7453 =  ( n20 ) & ( n7311 )  ;
assign n7454 =  ( n20 ) & ( n7313 )  ;
assign n7455 =  ( n20 ) & ( n7315 )  ;
assign n7456 =  ( n20 ) & ( n7317 )  ;
assign n7457 =  ( n20 ) & ( n7319 )  ;
assign n7458 =  ( n20 ) & ( n7321 )  ;
assign n7459 =  ( n20 ) & ( n7323 )  ;
assign n7460 =  ( n20 ) & ( n7325 )  ;
assign n7461 =  ( n20 ) & ( n7327 )  ;
assign n7462 =  ( n20 ) & ( n7329 )  ;
assign n7463 =  ( n20 ) & ( n7331 )  ;
assign n7464 =  ( n20 ) & ( n7333 )  ;
assign n7465 =  ( n20 ) & ( n7335 )  ;
assign n7466 =  ( n20 ) & ( n7337 )  ;
assign n7467 =  ( n21 ) & ( n7307 )  ;
assign n7468 =  ( n21 ) & ( n7309 )  ;
assign n7469 =  ( n21 ) & ( n7311 )  ;
assign n7470 =  ( n21 ) & ( n7313 )  ;
assign n7471 =  ( n21 ) & ( n7315 )  ;
assign n7472 =  ( n21 ) & ( n7317 )  ;
assign n7473 =  ( n21 ) & ( n7319 )  ;
assign n7474 =  ( n21 ) & ( n7321 )  ;
assign n7475 =  ( n21 ) & ( n7323 )  ;
assign n7476 =  ( n21 ) & ( n7325 )  ;
assign n7477 =  ( n21 ) & ( n7327 )  ;
assign n7478 =  ( n21 ) & ( n7329 )  ;
assign n7479 =  ( n21 ) & ( n7331 )  ;
assign n7480 =  ( n21 ) & ( n7333 )  ;
assign n7481 =  ( n21 ) & ( n7335 )  ;
assign n7482 =  ( n21 ) & ( n7337 )  ;
assign n7483 =  ( n22 ) & ( n7307 )  ;
assign n7484 =  ( n22 ) & ( n7309 )  ;
assign n7485 =  ( n22 ) & ( n7311 )  ;
assign n7486 =  ( n22 ) & ( n7313 )  ;
assign n7487 =  ( n22 ) & ( n7315 )  ;
assign n7488 =  ( n22 ) & ( n7317 )  ;
assign n7489 =  ( n22 ) & ( n7319 )  ;
assign n7490 =  ( n22 ) & ( n7321 )  ;
assign n7491 =  ( n22 ) & ( n7323 )  ;
assign n7492 =  ( n22 ) & ( n7325 )  ;
assign n7493 =  ( n22 ) & ( n7327 )  ;
assign n7494 =  ( n22 ) & ( n7329 )  ;
assign n7495 =  ( n22 ) & ( n7331 )  ;
assign n7496 =  ( n22 ) & ( n7333 )  ;
assign n7497 =  ( n22 ) & ( n7335 )  ;
assign n7498 =  ( n22 ) & ( n7337 )  ;
assign n7499 =  ( n23 ) & ( n7307 )  ;
assign n7500 =  ( n23 ) & ( n7309 )  ;
assign n7501 =  ( n23 ) & ( n7311 )  ;
assign n7502 =  ( n23 ) & ( n7313 )  ;
assign n7503 =  ( n23 ) & ( n7315 )  ;
assign n7504 =  ( n23 ) & ( n7317 )  ;
assign n7505 =  ( n23 ) & ( n7319 )  ;
assign n7506 =  ( n23 ) & ( n7321 )  ;
assign n7507 =  ( n23 ) & ( n7323 )  ;
assign n7508 =  ( n23 ) & ( n7325 )  ;
assign n7509 =  ( n23 ) & ( n7327 )  ;
assign n7510 =  ( n23 ) & ( n7329 )  ;
assign n7511 =  ( n23 ) & ( n7331 )  ;
assign n7512 =  ( n23 ) & ( n7333 )  ;
assign n7513 =  ( n23 ) & ( n7335 )  ;
assign n7514 =  ( n23 ) & ( n7337 )  ;
assign n7515 =  ( n24 ) & ( n7307 )  ;
assign n7516 =  ( n24 ) & ( n7309 )  ;
assign n7517 =  ( n24 ) & ( n7311 )  ;
assign n7518 =  ( n24 ) & ( n7313 )  ;
assign n7519 =  ( n24 ) & ( n7315 )  ;
assign n7520 =  ( n24 ) & ( n7317 )  ;
assign n7521 =  ( n24 ) & ( n7319 )  ;
assign n7522 =  ( n24 ) & ( n7321 )  ;
assign n7523 =  ( n24 ) & ( n7323 )  ;
assign n7524 =  ( n24 ) & ( n7325 )  ;
assign n7525 =  ( n24 ) & ( n7327 )  ;
assign n7526 =  ( n24 ) & ( n7329 )  ;
assign n7527 =  ( n24 ) & ( n7331 )  ;
assign n7528 =  ( n24 ) & ( n7333 )  ;
assign n7529 =  ( n24 ) & ( n7335 )  ;
assign n7530 =  ( n24 ) & ( n7337 )  ;
assign n7531 =  ( n25 ) & ( n7307 )  ;
assign n7532 =  ( n25 ) & ( n7309 )  ;
assign n7533 =  ( n25 ) & ( n7311 )  ;
assign n7534 =  ( n25 ) & ( n7313 )  ;
assign n7535 =  ( n25 ) & ( n7315 )  ;
assign n7536 =  ( n25 ) & ( n7317 )  ;
assign n7537 =  ( n25 ) & ( n7319 )  ;
assign n7538 =  ( n25 ) & ( n7321 )  ;
assign n7539 =  ( n25 ) & ( n7323 )  ;
assign n7540 =  ( n25 ) & ( n7325 )  ;
assign n7541 =  ( n25 ) & ( n7327 )  ;
assign n7542 =  ( n25 ) & ( n7329 )  ;
assign n7543 =  ( n25 ) & ( n7331 )  ;
assign n7544 =  ( n25 ) & ( n7333 )  ;
assign n7545 =  ( n25 ) & ( n7335 )  ;
assign n7546 =  ( n25 ) & ( n7337 )  ;
assign n7547 =  ( n26 ) & ( n7307 )  ;
assign n7548 =  ( n26 ) & ( n7309 )  ;
assign n7549 =  ( n26 ) & ( n7311 )  ;
assign n7550 =  ( n26 ) & ( n7313 )  ;
assign n7551 =  ( n26 ) & ( n7315 )  ;
assign n7552 =  ( n26 ) & ( n7317 )  ;
assign n7553 =  ( n26 ) & ( n7319 )  ;
assign n7554 =  ( n26 ) & ( n7321 )  ;
assign n7555 =  ( n26 ) & ( n7323 )  ;
assign n7556 =  ( n26 ) & ( n7325 )  ;
assign n7557 =  ( n26 ) & ( n7327 )  ;
assign n7558 =  ( n26 ) & ( n7329 )  ;
assign n7559 =  ( n26 ) & ( n7331 )  ;
assign n7560 =  ( n26 ) & ( n7333 )  ;
assign n7561 =  ( n26 ) & ( n7335 )  ;
assign n7562 =  ( n26 ) & ( n7337 )  ;
assign n7563 =  ( n27 ) & ( n7307 )  ;
assign n7564 =  ( n27 ) & ( n7309 )  ;
assign n7565 =  ( n27 ) & ( n7311 )  ;
assign n7566 =  ( n27 ) & ( n7313 )  ;
assign n7567 =  ( n27 ) & ( n7315 )  ;
assign n7568 =  ( n27 ) & ( n7317 )  ;
assign n7569 =  ( n27 ) & ( n7319 )  ;
assign n7570 =  ( n27 ) & ( n7321 )  ;
assign n7571 =  ( n27 ) & ( n7323 )  ;
assign n7572 =  ( n27 ) & ( n7325 )  ;
assign n7573 =  ( n27 ) & ( n7327 )  ;
assign n7574 =  ( n27 ) & ( n7329 )  ;
assign n7575 =  ( n27 ) & ( n7331 )  ;
assign n7576 =  ( n27 ) & ( n7333 )  ;
assign n7577 =  ( n27 ) & ( n7335 )  ;
assign n7578 =  ( n27 ) & ( n7337 )  ;
assign n7579 =  ( n28 ) & ( n7307 )  ;
assign n7580 =  ( n28 ) & ( n7309 )  ;
assign n7581 =  ( n28 ) & ( n7311 )  ;
assign n7582 =  ( n28 ) & ( n7313 )  ;
assign n7583 =  ( n28 ) & ( n7315 )  ;
assign n7584 =  ( n28 ) & ( n7317 )  ;
assign n7585 =  ( n28 ) & ( n7319 )  ;
assign n7586 =  ( n28 ) & ( n7321 )  ;
assign n7587 =  ( n28 ) & ( n7323 )  ;
assign n7588 =  ( n28 ) & ( n7325 )  ;
assign n7589 =  ( n28 ) & ( n7327 )  ;
assign n7590 =  ( n28 ) & ( n7329 )  ;
assign n7591 =  ( n28 ) & ( n7331 )  ;
assign n7592 =  ( n28 ) & ( n7333 )  ;
assign n7593 =  ( n28 ) & ( n7335 )  ;
assign n7594 =  ( n28 ) & ( n7337 )  ;
assign n7595 =  ( n29 ) & ( n7307 )  ;
assign n7596 =  ( n29 ) & ( n7309 )  ;
assign n7597 =  ( n29 ) & ( n7311 )  ;
assign n7598 =  ( n29 ) & ( n7313 )  ;
assign n7599 =  ( n29 ) & ( n7315 )  ;
assign n7600 =  ( n29 ) & ( n7317 )  ;
assign n7601 =  ( n29 ) & ( n7319 )  ;
assign n7602 =  ( n29 ) & ( n7321 )  ;
assign n7603 =  ( n29 ) & ( n7323 )  ;
assign n7604 =  ( n29 ) & ( n7325 )  ;
assign n7605 =  ( n29 ) & ( n7327 )  ;
assign n7606 =  ( n29 ) & ( n7329 )  ;
assign n7607 =  ( n29 ) & ( n7331 )  ;
assign n7608 =  ( n29 ) & ( n7333 )  ;
assign n7609 =  ( n29 ) & ( n7335 )  ;
assign n7610 =  ( n29 ) & ( n7337 )  ;
assign n7611 =  ( n30 ) & ( n7307 )  ;
assign n7612 =  ( n30 ) & ( n7309 )  ;
assign n7613 =  ( n30 ) & ( n7311 )  ;
assign n7614 =  ( n30 ) & ( n7313 )  ;
assign n7615 =  ( n30 ) & ( n7315 )  ;
assign n7616 =  ( n30 ) & ( n7317 )  ;
assign n7617 =  ( n30 ) & ( n7319 )  ;
assign n7618 =  ( n30 ) & ( n7321 )  ;
assign n7619 =  ( n30 ) & ( n7323 )  ;
assign n7620 =  ( n30 ) & ( n7325 )  ;
assign n7621 =  ( n30 ) & ( n7327 )  ;
assign n7622 =  ( n30 ) & ( n7329 )  ;
assign n7623 =  ( n30 ) & ( n7331 )  ;
assign n7624 =  ( n30 ) & ( n7333 )  ;
assign n7625 =  ( n30 ) & ( n7335 )  ;
assign n7626 =  ( n30 ) & ( n7337 )  ;
assign n7627 =  ( n31 ) & ( n7307 )  ;
assign n7628 =  ( n31 ) & ( n7309 )  ;
assign n7629 =  ( n31 ) & ( n7311 )  ;
assign n7630 =  ( n31 ) & ( n7313 )  ;
assign n7631 =  ( n31 ) & ( n7315 )  ;
assign n7632 =  ( n31 ) & ( n7317 )  ;
assign n7633 =  ( n31 ) & ( n7319 )  ;
assign n7634 =  ( n31 ) & ( n7321 )  ;
assign n7635 =  ( n31 ) & ( n7323 )  ;
assign n7636 =  ( n31 ) & ( n7325 )  ;
assign n7637 =  ( n31 ) & ( n7327 )  ;
assign n7638 =  ( n31 ) & ( n7329 )  ;
assign n7639 =  ( n31 ) & ( n7331 )  ;
assign n7640 =  ( n31 ) & ( n7333 )  ;
assign n7641 =  ( n31 ) & ( n7335 )  ;
assign n7642 =  ( n31 ) & ( n7337 )  ;
assign n7643 =  ( n32 ) & ( n7307 )  ;
assign n7644 =  ( n32 ) & ( n7309 )  ;
assign n7645 =  ( n32 ) & ( n7311 )  ;
assign n7646 =  ( n32 ) & ( n7313 )  ;
assign n7647 =  ( n32 ) & ( n7315 )  ;
assign n7648 =  ( n32 ) & ( n7317 )  ;
assign n7649 =  ( n32 ) & ( n7319 )  ;
assign n7650 =  ( n32 ) & ( n7321 )  ;
assign n7651 =  ( n32 ) & ( n7323 )  ;
assign n7652 =  ( n32 ) & ( n7325 )  ;
assign n7653 =  ( n32 ) & ( n7327 )  ;
assign n7654 =  ( n32 ) & ( n7329 )  ;
assign n7655 =  ( n32 ) & ( n7331 )  ;
assign n7656 =  ( n32 ) & ( n7333 )  ;
assign n7657 =  ( n32 ) & ( n7335 )  ;
assign n7658 =  ( n32 ) & ( n7337 )  ;
assign n7659 =  ( n33 ) & ( n7307 )  ;
assign n7660 =  ( n33 ) & ( n7309 )  ;
assign n7661 =  ( n33 ) & ( n7311 )  ;
assign n7662 =  ( n33 ) & ( n7313 )  ;
assign n7663 =  ( n33 ) & ( n7315 )  ;
assign n7664 =  ( n33 ) & ( n7317 )  ;
assign n7665 =  ( n33 ) & ( n7319 )  ;
assign n7666 =  ( n33 ) & ( n7321 )  ;
assign n7667 =  ( n33 ) & ( n7323 )  ;
assign n7668 =  ( n33 ) & ( n7325 )  ;
assign n7669 =  ( n33 ) & ( n7327 )  ;
assign n7670 =  ( n33 ) & ( n7329 )  ;
assign n7671 =  ( n33 ) & ( n7331 )  ;
assign n7672 =  ( n33 ) & ( n7333 )  ;
assign n7673 =  ( n33 ) & ( n7335 )  ;
assign n7674 =  ( n33 ) & ( n7337 )  ;
assign n7675 =  ( n34 ) & ( n7307 )  ;
assign n7676 =  ( n34 ) & ( n7309 )  ;
assign n7677 =  ( n34 ) & ( n7311 )  ;
assign n7678 =  ( n34 ) & ( n7313 )  ;
assign n7679 =  ( n34 ) & ( n7315 )  ;
assign n7680 =  ( n34 ) & ( n7317 )  ;
assign n7681 =  ( n34 ) & ( n7319 )  ;
assign n7682 =  ( n34 ) & ( n7321 )  ;
assign n7683 =  ( n34 ) & ( n7323 )  ;
assign n7684 =  ( n34 ) & ( n7325 )  ;
assign n7685 =  ( n34 ) & ( n7327 )  ;
assign n7686 =  ( n34 ) & ( n7329 )  ;
assign n7687 =  ( n34 ) & ( n7331 )  ;
assign n7688 =  ( n34 ) & ( n7333 )  ;
assign n7689 =  ( n34 ) & ( n7335 )  ;
assign n7690 =  ( n34 ) & ( n7337 )  ;
assign n7691 =  ( n35 ) & ( n7307 )  ;
assign n7692 =  ( n35 ) & ( n7309 )  ;
assign n7693 =  ( n35 ) & ( n7311 )  ;
assign n7694 =  ( n35 ) & ( n7313 )  ;
assign n7695 =  ( n35 ) & ( n7315 )  ;
assign n7696 =  ( n35 ) & ( n7317 )  ;
assign n7697 =  ( n35 ) & ( n7319 )  ;
assign n7698 =  ( n35 ) & ( n7321 )  ;
assign n7699 =  ( n35 ) & ( n7323 )  ;
assign n7700 =  ( n35 ) & ( n7325 )  ;
assign n7701 =  ( n35 ) & ( n7327 )  ;
assign n7702 =  ( n35 ) & ( n7329 )  ;
assign n7703 =  ( n35 ) & ( n7331 )  ;
assign n7704 =  ( n35 ) & ( n7333 )  ;
assign n7705 =  ( n35 ) & ( n7335 )  ;
assign n7706 =  ( n35 ) & ( n7337 )  ;
assign n7707 =  ( n36 ) & ( n7307 )  ;
assign n7708 =  ( n36 ) & ( n7309 )  ;
assign n7709 =  ( n36 ) & ( n7311 )  ;
assign n7710 =  ( n36 ) & ( n7313 )  ;
assign n7711 =  ( n36 ) & ( n7315 )  ;
assign n7712 =  ( n36 ) & ( n7317 )  ;
assign n7713 =  ( n36 ) & ( n7319 )  ;
assign n7714 =  ( n36 ) & ( n7321 )  ;
assign n7715 =  ( n36 ) & ( n7323 )  ;
assign n7716 =  ( n36 ) & ( n7325 )  ;
assign n7717 =  ( n36 ) & ( n7327 )  ;
assign n7718 =  ( n36 ) & ( n7329 )  ;
assign n7719 =  ( n36 ) & ( n7331 )  ;
assign n7720 =  ( n36 ) & ( n7333 )  ;
assign n7721 =  ( n36 ) & ( n7335 )  ;
assign n7722 =  ( n36 ) & ( n7337 )  ;
assign n7723 =  ( n37 ) & ( n7307 )  ;
assign n7724 =  ( n37 ) & ( n7309 )  ;
assign n7725 =  ( n37 ) & ( n7311 )  ;
assign n7726 =  ( n37 ) & ( n7313 )  ;
assign n7727 =  ( n37 ) & ( n7315 )  ;
assign n7728 =  ( n37 ) & ( n7317 )  ;
assign n7729 =  ( n37 ) & ( n7319 )  ;
assign n7730 =  ( n37 ) & ( n7321 )  ;
assign n7731 =  ( n37 ) & ( n7323 )  ;
assign n7732 =  ( n37 ) & ( n7325 )  ;
assign n7733 =  ( n37 ) & ( n7327 )  ;
assign n7734 =  ( n37 ) & ( n7329 )  ;
assign n7735 =  ( n37 ) & ( n7331 )  ;
assign n7736 =  ( n37 ) & ( n7333 )  ;
assign n7737 =  ( n37 ) & ( n7335 )  ;
assign n7738 =  ( n37 ) & ( n7337 )  ;
assign n7739 =  ( n38 ) & ( n7307 )  ;
assign n7740 =  ( n38 ) & ( n7309 )  ;
assign n7741 =  ( n38 ) & ( n7311 )  ;
assign n7742 =  ( n38 ) & ( n7313 )  ;
assign n7743 =  ( n38 ) & ( n7315 )  ;
assign n7744 =  ( n38 ) & ( n7317 )  ;
assign n7745 =  ( n38 ) & ( n7319 )  ;
assign n7746 =  ( n38 ) & ( n7321 )  ;
assign n7747 =  ( n38 ) & ( n7323 )  ;
assign n7748 =  ( n38 ) & ( n7325 )  ;
assign n7749 =  ( n38 ) & ( n7327 )  ;
assign n7750 =  ( n38 ) & ( n7329 )  ;
assign n7751 =  ( n38 ) & ( n7331 )  ;
assign n7752 =  ( n38 ) & ( n7333 )  ;
assign n7753 =  ( n38 ) & ( n7335 )  ;
assign n7754 =  ( n38 ) & ( n7337 )  ;
assign n7755 =  ( n39 ) & ( n7307 )  ;
assign n7756 =  ( n39 ) & ( n7309 )  ;
assign n7757 =  ( n39 ) & ( n7311 )  ;
assign n7758 =  ( n39 ) & ( n7313 )  ;
assign n7759 =  ( n39 ) & ( n7315 )  ;
assign n7760 =  ( n39 ) & ( n7317 )  ;
assign n7761 =  ( n39 ) & ( n7319 )  ;
assign n7762 =  ( n39 ) & ( n7321 )  ;
assign n7763 =  ( n39 ) & ( n7323 )  ;
assign n7764 =  ( n39 ) & ( n7325 )  ;
assign n7765 =  ( n39 ) & ( n7327 )  ;
assign n7766 =  ( n39 ) & ( n7329 )  ;
assign n7767 =  ( n39 ) & ( n7331 )  ;
assign n7768 =  ( n39 ) & ( n7333 )  ;
assign n7769 =  ( n39 ) & ( n7335 )  ;
assign n7770 =  ( n39 ) & ( n7337 )  ;
assign n7771 =  ( n40 ) & ( n7307 )  ;
assign n7772 =  ( n40 ) & ( n7309 )  ;
assign n7773 =  ( n40 ) & ( n7311 )  ;
assign n7774 =  ( n40 ) & ( n7313 )  ;
assign n7775 =  ( n40 ) & ( n7315 )  ;
assign n7776 =  ( n40 ) & ( n7317 )  ;
assign n7777 =  ( n40 ) & ( n7319 )  ;
assign n7778 =  ( n40 ) & ( n7321 )  ;
assign n7779 =  ( n40 ) & ( n7323 )  ;
assign n7780 =  ( n40 ) & ( n7325 )  ;
assign n7781 =  ( n40 ) & ( n7327 )  ;
assign n7782 =  ( n40 ) & ( n7329 )  ;
assign n7783 =  ( n40 ) & ( n7331 )  ;
assign n7784 =  ( n40 ) & ( n7333 )  ;
assign n7785 =  ( n40 ) & ( n7335 )  ;
assign n7786 =  ( n40 ) & ( n7337 )  ;
assign n7787 =  ( n41 ) & ( n7307 )  ;
assign n7788 =  ( n41 ) & ( n7309 )  ;
assign n7789 =  ( n41 ) & ( n7311 )  ;
assign n7790 =  ( n41 ) & ( n7313 )  ;
assign n7791 =  ( n41 ) & ( n7315 )  ;
assign n7792 =  ( n41 ) & ( n7317 )  ;
assign n7793 =  ( n41 ) & ( n7319 )  ;
assign n7794 =  ( n41 ) & ( n7321 )  ;
assign n7795 =  ( n41 ) & ( n7323 )  ;
assign n7796 =  ( n41 ) & ( n7325 )  ;
assign n7797 =  ( n41 ) & ( n7327 )  ;
assign n7798 =  ( n41 ) & ( n7329 )  ;
assign n7799 =  ( n41 ) & ( n7331 )  ;
assign n7800 =  ( n41 ) & ( n7333 )  ;
assign n7801 =  ( n41 ) & ( n7335 )  ;
assign n7802 =  ( n41 ) & ( n7337 )  ;
assign n7803 =  ( n42 ) & ( n7307 )  ;
assign n7804 =  ( n42 ) & ( n7309 )  ;
assign n7805 =  ( n42 ) & ( n7311 )  ;
assign n7806 =  ( n42 ) & ( n7313 )  ;
assign n7807 =  ( n42 ) & ( n7315 )  ;
assign n7808 =  ( n42 ) & ( n7317 )  ;
assign n7809 =  ( n42 ) & ( n7319 )  ;
assign n7810 =  ( n42 ) & ( n7321 )  ;
assign n7811 =  ( n42 ) & ( n7323 )  ;
assign n7812 =  ( n42 ) & ( n7325 )  ;
assign n7813 =  ( n42 ) & ( n7327 )  ;
assign n7814 =  ( n42 ) & ( n7329 )  ;
assign n7815 =  ( n42 ) & ( n7331 )  ;
assign n7816 =  ( n42 ) & ( n7333 )  ;
assign n7817 =  ( n42 ) & ( n7335 )  ;
assign n7818 =  ( n42 ) & ( n7337 )  ;
assign n7819 =  ( n43 ) & ( n7307 )  ;
assign n7820 =  ( n43 ) & ( n7309 )  ;
assign n7821 =  ( n43 ) & ( n7311 )  ;
assign n7822 =  ( n43 ) & ( n7313 )  ;
assign n7823 =  ( n43 ) & ( n7315 )  ;
assign n7824 =  ( n43 ) & ( n7317 )  ;
assign n7825 =  ( n43 ) & ( n7319 )  ;
assign n7826 =  ( n43 ) & ( n7321 )  ;
assign n7827 =  ( n43 ) & ( n7323 )  ;
assign n7828 =  ( n43 ) & ( n7325 )  ;
assign n7829 =  ( n43 ) & ( n7327 )  ;
assign n7830 =  ( n43 ) & ( n7329 )  ;
assign n7831 =  ( n43 ) & ( n7331 )  ;
assign n7832 =  ( n43 ) & ( n7333 )  ;
assign n7833 =  ( n43 ) & ( n7335 )  ;
assign n7834 =  ( n43 ) & ( n7337 )  ;
assign n7835 =  ( n7834 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n7836 =  ( n7833 ) ? ( VREG_0_1 ) : ( n7835 ) ;
assign n7837 =  ( n7832 ) ? ( VREG_0_2 ) : ( n7836 ) ;
assign n7838 =  ( n7831 ) ? ( VREG_0_3 ) : ( n7837 ) ;
assign n7839 =  ( n7830 ) ? ( VREG_0_4 ) : ( n7838 ) ;
assign n7840 =  ( n7829 ) ? ( VREG_0_5 ) : ( n7839 ) ;
assign n7841 =  ( n7828 ) ? ( VREG_0_6 ) : ( n7840 ) ;
assign n7842 =  ( n7827 ) ? ( VREG_0_7 ) : ( n7841 ) ;
assign n7843 =  ( n7826 ) ? ( VREG_0_8 ) : ( n7842 ) ;
assign n7844 =  ( n7825 ) ? ( VREG_0_9 ) : ( n7843 ) ;
assign n7845 =  ( n7824 ) ? ( VREG_0_10 ) : ( n7844 ) ;
assign n7846 =  ( n7823 ) ? ( VREG_0_11 ) : ( n7845 ) ;
assign n7847 =  ( n7822 ) ? ( VREG_0_12 ) : ( n7846 ) ;
assign n7848 =  ( n7821 ) ? ( VREG_0_13 ) : ( n7847 ) ;
assign n7849 =  ( n7820 ) ? ( VREG_0_14 ) : ( n7848 ) ;
assign n7850 =  ( n7819 ) ? ( VREG_0_15 ) : ( n7849 ) ;
assign n7851 =  ( n7818 ) ? ( VREG_1_0 ) : ( n7850 ) ;
assign n7852 =  ( n7817 ) ? ( VREG_1_1 ) : ( n7851 ) ;
assign n7853 =  ( n7816 ) ? ( VREG_1_2 ) : ( n7852 ) ;
assign n7854 =  ( n7815 ) ? ( VREG_1_3 ) : ( n7853 ) ;
assign n7855 =  ( n7814 ) ? ( VREG_1_4 ) : ( n7854 ) ;
assign n7856 =  ( n7813 ) ? ( VREG_1_5 ) : ( n7855 ) ;
assign n7857 =  ( n7812 ) ? ( VREG_1_6 ) : ( n7856 ) ;
assign n7858 =  ( n7811 ) ? ( VREG_1_7 ) : ( n7857 ) ;
assign n7859 =  ( n7810 ) ? ( VREG_1_8 ) : ( n7858 ) ;
assign n7860 =  ( n7809 ) ? ( VREG_1_9 ) : ( n7859 ) ;
assign n7861 =  ( n7808 ) ? ( VREG_1_10 ) : ( n7860 ) ;
assign n7862 =  ( n7807 ) ? ( VREG_1_11 ) : ( n7861 ) ;
assign n7863 =  ( n7806 ) ? ( VREG_1_12 ) : ( n7862 ) ;
assign n7864 =  ( n7805 ) ? ( VREG_1_13 ) : ( n7863 ) ;
assign n7865 =  ( n7804 ) ? ( VREG_1_14 ) : ( n7864 ) ;
assign n7866 =  ( n7803 ) ? ( VREG_1_15 ) : ( n7865 ) ;
assign n7867 =  ( n7802 ) ? ( VREG_2_0 ) : ( n7866 ) ;
assign n7868 =  ( n7801 ) ? ( VREG_2_1 ) : ( n7867 ) ;
assign n7869 =  ( n7800 ) ? ( VREG_2_2 ) : ( n7868 ) ;
assign n7870 =  ( n7799 ) ? ( VREG_2_3 ) : ( n7869 ) ;
assign n7871 =  ( n7798 ) ? ( VREG_2_4 ) : ( n7870 ) ;
assign n7872 =  ( n7797 ) ? ( VREG_2_5 ) : ( n7871 ) ;
assign n7873 =  ( n7796 ) ? ( VREG_2_6 ) : ( n7872 ) ;
assign n7874 =  ( n7795 ) ? ( VREG_2_7 ) : ( n7873 ) ;
assign n7875 =  ( n7794 ) ? ( VREG_2_8 ) : ( n7874 ) ;
assign n7876 =  ( n7793 ) ? ( VREG_2_9 ) : ( n7875 ) ;
assign n7877 =  ( n7792 ) ? ( VREG_2_10 ) : ( n7876 ) ;
assign n7878 =  ( n7791 ) ? ( VREG_2_11 ) : ( n7877 ) ;
assign n7879 =  ( n7790 ) ? ( VREG_2_12 ) : ( n7878 ) ;
assign n7880 =  ( n7789 ) ? ( VREG_2_13 ) : ( n7879 ) ;
assign n7881 =  ( n7788 ) ? ( VREG_2_14 ) : ( n7880 ) ;
assign n7882 =  ( n7787 ) ? ( VREG_2_15 ) : ( n7881 ) ;
assign n7883 =  ( n7786 ) ? ( VREG_3_0 ) : ( n7882 ) ;
assign n7884 =  ( n7785 ) ? ( VREG_3_1 ) : ( n7883 ) ;
assign n7885 =  ( n7784 ) ? ( VREG_3_2 ) : ( n7884 ) ;
assign n7886 =  ( n7783 ) ? ( VREG_3_3 ) : ( n7885 ) ;
assign n7887 =  ( n7782 ) ? ( VREG_3_4 ) : ( n7886 ) ;
assign n7888 =  ( n7781 ) ? ( VREG_3_5 ) : ( n7887 ) ;
assign n7889 =  ( n7780 ) ? ( VREG_3_6 ) : ( n7888 ) ;
assign n7890 =  ( n7779 ) ? ( VREG_3_7 ) : ( n7889 ) ;
assign n7891 =  ( n7778 ) ? ( VREG_3_8 ) : ( n7890 ) ;
assign n7892 =  ( n7777 ) ? ( VREG_3_9 ) : ( n7891 ) ;
assign n7893 =  ( n7776 ) ? ( VREG_3_10 ) : ( n7892 ) ;
assign n7894 =  ( n7775 ) ? ( VREG_3_11 ) : ( n7893 ) ;
assign n7895 =  ( n7774 ) ? ( VREG_3_12 ) : ( n7894 ) ;
assign n7896 =  ( n7773 ) ? ( VREG_3_13 ) : ( n7895 ) ;
assign n7897 =  ( n7772 ) ? ( VREG_3_14 ) : ( n7896 ) ;
assign n7898 =  ( n7771 ) ? ( VREG_3_15 ) : ( n7897 ) ;
assign n7899 =  ( n7770 ) ? ( VREG_4_0 ) : ( n7898 ) ;
assign n7900 =  ( n7769 ) ? ( VREG_4_1 ) : ( n7899 ) ;
assign n7901 =  ( n7768 ) ? ( VREG_4_2 ) : ( n7900 ) ;
assign n7902 =  ( n7767 ) ? ( VREG_4_3 ) : ( n7901 ) ;
assign n7903 =  ( n7766 ) ? ( VREG_4_4 ) : ( n7902 ) ;
assign n7904 =  ( n7765 ) ? ( VREG_4_5 ) : ( n7903 ) ;
assign n7905 =  ( n7764 ) ? ( VREG_4_6 ) : ( n7904 ) ;
assign n7906 =  ( n7763 ) ? ( VREG_4_7 ) : ( n7905 ) ;
assign n7907 =  ( n7762 ) ? ( VREG_4_8 ) : ( n7906 ) ;
assign n7908 =  ( n7761 ) ? ( VREG_4_9 ) : ( n7907 ) ;
assign n7909 =  ( n7760 ) ? ( VREG_4_10 ) : ( n7908 ) ;
assign n7910 =  ( n7759 ) ? ( VREG_4_11 ) : ( n7909 ) ;
assign n7911 =  ( n7758 ) ? ( VREG_4_12 ) : ( n7910 ) ;
assign n7912 =  ( n7757 ) ? ( VREG_4_13 ) : ( n7911 ) ;
assign n7913 =  ( n7756 ) ? ( VREG_4_14 ) : ( n7912 ) ;
assign n7914 =  ( n7755 ) ? ( VREG_4_15 ) : ( n7913 ) ;
assign n7915 =  ( n7754 ) ? ( VREG_5_0 ) : ( n7914 ) ;
assign n7916 =  ( n7753 ) ? ( VREG_5_1 ) : ( n7915 ) ;
assign n7917 =  ( n7752 ) ? ( VREG_5_2 ) : ( n7916 ) ;
assign n7918 =  ( n7751 ) ? ( VREG_5_3 ) : ( n7917 ) ;
assign n7919 =  ( n7750 ) ? ( VREG_5_4 ) : ( n7918 ) ;
assign n7920 =  ( n7749 ) ? ( VREG_5_5 ) : ( n7919 ) ;
assign n7921 =  ( n7748 ) ? ( VREG_5_6 ) : ( n7920 ) ;
assign n7922 =  ( n7747 ) ? ( VREG_5_7 ) : ( n7921 ) ;
assign n7923 =  ( n7746 ) ? ( VREG_5_8 ) : ( n7922 ) ;
assign n7924 =  ( n7745 ) ? ( VREG_5_9 ) : ( n7923 ) ;
assign n7925 =  ( n7744 ) ? ( VREG_5_10 ) : ( n7924 ) ;
assign n7926 =  ( n7743 ) ? ( VREG_5_11 ) : ( n7925 ) ;
assign n7927 =  ( n7742 ) ? ( VREG_5_12 ) : ( n7926 ) ;
assign n7928 =  ( n7741 ) ? ( VREG_5_13 ) : ( n7927 ) ;
assign n7929 =  ( n7740 ) ? ( VREG_5_14 ) : ( n7928 ) ;
assign n7930 =  ( n7739 ) ? ( VREG_5_15 ) : ( n7929 ) ;
assign n7931 =  ( n7738 ) ? ( VREG_6_0 ) : ( n7930 ) ;
assign n7932 =  ( n7737 ) ? ( VREG_6_1 ) : ( n7931 ) ;
assign n7933 =  ( n7736 ) ? ( VREG_6_2 ) : ( n7932 ) ;
assign n7934 =  ( n7735 ) ? ( VREG_6_3 ) : ( n7933 ) ;
assign n7935 =  ( n7734 ) ? ( VREG_6_4 ) : ( n7934 ) ;
assign n7936 =  ( n7733 ) ? ( VREG_6_5 ) : ( n7935 ) ;
assign n7937 =  ( n7732 ) ? ( VREG_6_6 ) : ( n7936 ) ;
assign n7938 =  ( n7731 ) ? ( VREG_6_7 ) : ( n7937 ) ;
assign n7939 =  ( n7730 ) ? ( VREG_6_8 ) : ( n7938 ) ;
assign n7940 =  ( n7729 ) ? ( VREG_6_9 ) : ( n7939 ) ;
assign n7941 =  ( n7728 ) ? ( VREG_6_10 ) : ( n7940 ) ;
assign n7942 =  ( n7727 ) ? ( VREG_6_11 ) : ( n7941 ) ;
assign n7943 =  ( n7726 ) ? ( VREG_6_12 ) : ( n7942 ) ;
assign n7944 =  ( n7725 ) ? ( VREG_6_13 ) : ( n7943 ) ;
assign n7945 =  ( n7724 ) ? ( VREG_6_14 ) : ( n7944 ) ;
assign n7946 =  ( n7723 ) ? ( VREG_6_15 ) : ( n7945 ) ;
assign n7947 =  ( n7722 ) ? ( VREG_7_0 ) : ( n7946 ) ;
assign n7948 =  ( n7721 ) ? ( VREG_7_1 ) : ( n7947 ) ;
assign n7949 =  ( n7720 ) ? ( VREG_7_2 ) : ( n7948 ) ;
assign n7950 =  ( n7719 ) ? ( VREG_7_3 ) : ( n7949 ) ;
assign n7951 =  ( n7718 ) ? ( VREG_7_4 ) : ( n7950 ) ;
assign n7952 =  ( n7717 ) ? ( VREG_7_5 ) : ( n7951 ) ;
assign n7953 =  ( n7716 ) ? ( VREG_7_6 ) : ( n7952 ) ;
assign n7954 =  ( n7715 ) ? ( VREG_7_7 ) : ( n7953 ) ;
assign n7955 =  ( n7714 ) ? ( VREG_7_8 ) : ( n7954 ) ;
assign n7956 =  ( n7713 ) ? ( VREG_7_9 ) : ( n7955 ) ;
assign n7957 =  ( n7712 ) ? ( VREG_7_10 ) : ( n7956 ) ;
assign n7958 =  ( n7711 ) ? ( VREG_7_11 ) : ( n7957 ) ;
assign n7959 =  ( n7710 ) ? ( VREG_7_12 ) : ( n7958 ) ;
assign n7960 =  ( n7709 ) ? ( VREG_7_13 ) : ( n7959 ) ;
assign n7961 =  ( n7708 ) ? ( VREG_7_14 ) : ( n7960 ) ;
assign n7962 =  ( n7707 ) ? ( VREG_7_15 ) : ( n7961 ) ;
assign n7963 =  ( n7706 ) ? ( VREG_8_0 ) : ( n7962 ) ;
assign n7964 =  ( n7705 ) ? ( VREG_8_1 ) : ( n7963 ) ;
assign n7965 =  ( n7704 ) ? ( VREG_8_2 ) : ( n7964 ) ;
assign n7966 =  ( n7703 ) ? ( VREG_8_3 ) : ( n7965 ) ;
assign n7967 =  ( n7702 ) ? ( VREG_8_4 ) : ( n7966 ) ;
assign n7968 =  ( n7701 ) ? ( VREG_8_5 ) : ( n7967 ) ;
assign n7969 =  ( n7700 ) ? ( VREG_8_6 ) : ( n7968 ) ;
assign n7970 =  ( n7699 ) ? ( VREG_8_7 ) : ( n7969 ) ;
assign n7971 =  ( n7698 ) ? ( VREG_8_8 ) : ( n7970 ) ;
assign n7972 =  ( n7697 ) ? ( VREG_8_9 ) : ( n7971 ) ;
assign n7973 =  ( n7696 ) ? ( VREG_8_10 ) : ( n7972 ) ;
assign n7974 =  ( n7695 ) ? ( VREG_8_11 ) : ( n7973 ) ;
assign n7975 =  ( n7694 ) ? ( VREG_8_12 ) : ( n7974 ) ;
assign n7976 =  ( n7693 ) ? ( VREG_8_13 ) : ( n7975 ) ;
assign n7977 =  ( n7692 ) ? ( VREG_8_14 ) : ( n7976 ) ;
assign n7978 =  ( n7691 ) ? ( VREG_8_15 ) : ( n7977 ) ;
assign n7979 =  ( n7690 ) ? ( VREG_9_0 ) : ( n7978 ) ;
assign n7980 =  ( n7689 ) ? ( VREG_9_1 ) : ( n7979 ) ;
assign n7981 =  ( n7688 ) ? ( VREG_9_2 ) : ( n7980 ) ;
assign n7982 =  ( n7687 ) ? ( VREG_9_3 ) : ( n7981 ) ;
assign n7983 =  ( n7686 ) ? ( VREG_9_4 ) : ( n7982 ) ;
assign n7984 =  ( n7685 ) ? ( VREG_9_5 ) : ( n7983 ) ;
assign n7985 =  ( n7684 ) ? ( VREG_9_6 ) : ( n7984 ) ;
assign n7986 =  ( n7683 ) ? ( VREG_9_7 ) : ( n7985 ) ;
assign n7987 =  ( n7682 ) ? ( VREG_9_8 ) : ( n7986 ) ;
assign n7988 =  ( n7681 ) ? ( VREG_9_9 ) : ( n7987 ) ;
assign n7989 =  ( n7680 ) ? ( VREG_9_10 ) : ( n7988 ) ;
assign n7990 =  ( n7679 ) ? ( VREG_9_11 ) : ( n7989 ) ;
assign n7991 =  ( n7678 ) ? ( VREG_9_12 ) : ( n7990 ) ;
assign n7992 =  ( n7677 ) ? ( VREG_9_13 ) : ( n7991 ) ;
assign n7993 =  ( n7676 ) ? ( VREG_9_14 ) : ( n7992 ) ;
assign n7994 =  ( n7675 ) ? ( VREG_9_15 ) : ( n7993 ) ;
assign n7995 =  ( n7674 ) ? ( VREG_10_0 ) : ( n7994 ) ;
assign n7996 =  ( n7673 ) ? ( VREG_10_1 ) : ( n7995 ) ;
assign n7997 =  ( n7672 ) ? ( VREG_10_2 ) : ( n7996 ) ;
assign n7998 =  ( n7671 ) ? ( VREG_10_3 ) : ( n7997 ) ;
assign n7999 =  ( n7670 ) ? ( VREG_10_4 ) : ( n7998 ) ;
assign n8000 =  ( n7669 ) ? ( VREG_10_5 ) : ( n7999 ) ;
assign n8001 =  ( n7668 ) ? ( VREG_10_6 ) : ( n8000 ) ;
assign n8002 =  ( n7667 ) ? ( VREG_10_7 ) : ( n8001 ) ;
assign n8003 =  ( n7666 ) ? ( VREG_10_8 ) : ( n8002 ) ;
assign n8004 =  ( n7665 ) ? ( VREG_10_9 ) : ( n8003 ) ;
assign n8005 =  ( n7664 ) ? ( VREG_10_10 ) : ( n8004 ) ;
assign n8006 =  ( n7663 ) ? ( VREG_10_11 ) : ( n8005 ) ;
assign n8007 =  ( n7662 ) ? ( VREG_10_12 ) : ( n8006 ) ;
assign n8008 =  ( n7661 ) ? ( VREG_10_13 ) : ( n8007 ) ;
assign n8009 =  ( n7660 ) ? ( VREG_10_14 ) : ( n8008 ) ;
assign n8010 =  ( n7659 ) ? ( VREG_10_15 ) : ( n8009 ) ;
assign n8011 =  ( n7658 ) ? ( VREG_11_0 ) : ( n8010 ) ;
assign n8012 =  ( n7657 ) ? ( VREG_11_1 ) : ( n8011 ) ;
assign n8013 =  ( n7656 ) ? ( VREG_11_2 ) : ( n8012 ) ;
assign n8014 =  ( n7655 ) ? ( VREG_11_3 ) : ( n8013 ) ;
assign n8015 =  ( n7654 ) ? ( VREG_11_4 ) : ( n8014 ) ;
assign n8016 =  ( n7653 ) ? ( VREG_11_5 ) : ( n8015 ) ;
assign n8017 =  ( n7652 ) ? ( VREG_11_6 ) : ( n8016 ) ;
assign n8018 =  ( n7651 ) ? ( VREG_11_7 ) : ( n8017 ) ;
assign n8019 =  ( n7650 ) ? ( VREG_11_8 ) : ( n8018 ) ;
assign n8020 =  ( n7649 ) ? ( VREG_11_9 ) : ( n8019 ) ;
assign n8021 =  ( n7648 ) ? ( VREG_11_10 ) : ( n8020 ) ;
assign n8022 =  ( n7647 ) ? ( VREG_11_11 ) : ( n8021 ) ;
assign n8023 =  ( n7646 ) ? ( VREG_11_12 ) : ( n8022 ) ;
assign n8024 =  ( n7645 ) ? ( VREG_11_13 ) : ( n8023 ) ;
assign n8025 =  ( n7644 ) ? ( VREG_11_14 ) : ( n8024 ) ;
assign n8026 =  ( n7643 ) ? ( VREG_11_15 ) : ( n8025 ) ;
assign n8027 =  ( n7642 ) ? ( VREG_12_0 ) : ( n8026 ) ;
assign n8028 =  ( n7641 ) ? ( VREG_12_1 ) : ( n8027 ) ;
assign n8029 =  ( n7640 ) ? ( VREG_12_2 ) : ( n8028 ) ;
assign n8030 =  ( n7639 ) ? ( VREG_12_3 ) : ( n8029 ) ;
assign n8031 =  ( n7638 ) ? ( VREG_12_4 ) : ( n8030 ) ;
assign n8032 =  ( n7637 ) ? ( VREG_12_5 ) : ( n8031 ) ;
assign n8033 =  ( n7636 ) ? ( VREG_12_6 ) : ( n8032 ) ;
assign n8034 =  ( n7635 ) ? ( VREG_12_7 ) : ( n8033 ) ;
assign n8035 =  ( n7634 ) ? ( VREG_12_8 ) : ( n8034 ) ;
assign n8036 =  ( n7633 ) ? ( VREG_12_9 ) : ( n8035 ) ;
assign n8037 =  ( n7632 ) ? ( VREG_12_10 ) : ( n8036 ) ;
assign n8038 =  ( n7631 ) ? ( VREG_12_11 ) : ( n8037 ) ;
assign n8039 =  ( n7630 ) ? ( VREG_12_12 ) : ( n8038 ) ;
assign n8040 =  ( n7629 ) ? ( VREG_12_13 ) : ( n8039 ) ;
assign n8041 =  ( n7628 ) ? ( VREG_12_14 ) : ( n8040 ) ;
assign n8042 =  ( n7627 ) ? ( VREG_12_15 ) : ( n8041 ) ;
assign n8043 =  ( n7626 ) ? ( VREG_13_0 ) : ( n8042 ) ;
assign n8044 =  ( n7625 ) ? ( VREG_13_1 ) : ( n8043 ) ;
assign n8045 =  ( n7624 ) ? ( VREG_13_2 ) : ( n8044 ) ;
assign n8046 =  ( n7623 ) ? ( VREG_13_3 ) : ( n8045 ) ;
assign n8047 =  ( n7622 ) ? ( VREG_13_4 ) : ( n8046 ) ;
assign n8048 =  ( n7621 ) ? ( VREG_13_5 ) : ( n8047 ) ;
assign n8049 =  ( n7620 ) ? ( VREG_13_6 ) : ( n8048 ) ;
assign n8050 =  ( n7619 ) ? ( VREG_13_7 ) : ( n8049 ) ;
assign n8051 =  ( n7618 ) ? ( VREG_13_8 ) : ( n8050 ) ;
assign n8052 =  ( n7617 ) ? ( VREG_13_9 ) : ( n8051 ) ;
assign n8053 =  ( n7616 ) ? ( VREG_13_10 ) : ( n8052 ) ;
assign n8054 =  ( n7615 ) ? ( VREG_13_11 ) : ( n8053 ) ;
assign n8055 =  ( n7614 ) ? ( VREG_13_12 ) : ( n8054 ) ;
assign n8056 =  ( n7613 ) ? ( VREG_13_13 ) : ( n8055 ) ;
assign n8057 =  ( n7612 ) ? ( VREG_13_14 ) : ( n8056 ) ;
assign n8058 =  ( n7611 ) ? ( VREG_13_15 ) : ( n8057 ) ;
assign n8059 =  ( n7610 ) ? ( VREG_14_0 ) : ( n8058 ) ;
assign n8060 =  ( n7609 ) ? ( VREG_14_1 ) : ( n8059 ) ;
assign n8061 =  ( n7608 ) ? ( VREG_14_2 ) : ( n8060 ) ;
assign n8062 =  ( n7607 ) ? ( VREG_14_3 ) : ( n8061 ) ;
assign n8063 =  ( n7606 ) ? ( VREG_14_4 ) : ( n8062 ) ;
assign n8064 =  ( n7605 ) ? ( VREG_14_5 ) : ( n8063 ) ;
assign n8065 =  ( n7604 ) ? ( VREG_14_6 ) : ( n8064 ) ;
assign n8066 =  ( n7603 ) ? ( VREG_14_7 ) : ( n8065 ) ;
assign n8067 =  ( n7602 ) ? ( VREG_14_8 ) : ( n8066 ) ;
assign n8068 =  ( n7601 ) ? ( VREG_14_9 ) : ( n8067 ) ;
assign n8069 =  ( n7600 ) ? ( VREG_14_10 ) : ( n8068 ) ;
assign n8070 =  ( n7599 ) ? ( VREG_14_11 ) : ( n8069 ) ;
assign n8071 =  ( n7598 ) ? ( VREG_14_12 ) : ( n8070 ) ;
assign n8072 =  ( n7597 ) ? ( VREG_14_13 ) : ( n8071 ) ;
assign n8073 =  ( n7596 ) ? ( VREG_14_14 ) : ( n8072 ) ;
assign n8074 =  ( n7595 ) ? ( VREG_14_15 ) : ( n8073 ) ;
assign n8075 =  ( n7594 ) ? ( VREG_15_0 ) : ( n8074 ) ;
assign n8076 =  ( n7593 ) ? ( VREG_15_1 ) : ( n8075 ) ;
assign n8077 =  ( n7592 ) ? ( VREG_15_2 ) : ( n8076 ) ;
assign n8078 =  ( n7591 ) ? ( VREG_15_3 ) : ( n8077 ) ;
assign n8079 =  ( n7590 ) ? ( VREG_15_4 ) : ( n8078 ) ;
assign n8080 =  ( n7589 ) ? ( VREG_15_5 ) : ( n8079 ) ;
assign n8081 =  ( n7588 ) ? ( VREG_15_6 ) : ( n8080 ) ;
assign n8082 =  ( n7587 ) ? ( VREG_15_7 ) : ( n8081 ) ;
assign n8083 =  ( n7586 ) ? ( VREG_15_8 ) : ( n8082 ) ;
assign n8084 =  ( n7585 ) ? ( VREG_15_9 ) : ( n8083 ) ;
assign n8085 =  ( n7584 ) ? ( VREG_15_10 ) : ( n8084 ) ;
assign n8086 =  ( n7583 ) ? ( VREG_15_11 ) : ( n8085 ) ;
assign n8087 =  ( n7582 ) ? ( VREG_15_12 ) : ( n8086 ) ;
assign n8088 =  ( n7581 ) ? ( VREG_15_13 ) : ( n8087 ) ;
assign n8089 =  ( n7580 ) ? ( VREG_15_14 ) : ( n8088 ) ;
assign n8090 =  ( n7579 ) ? ( VREG_15_15 ) : ( n8089 ) ;
assign n8091 =  ( n7578 ) ? ( VREG_16_0 ) : ( n8090 ) ;
assign n8092 =  ( n7577 ) ? ( VREG_16_1 ) : ( n8091 ) ;
assign n8093 =  ( n7576 ) ? ( VREG_16_2 ) : ( n8092 ) ;
assign n8094 =  ( n7575 ) ? ( VREG_16_3 ) : ( n8093 ) ;
assign n8095 =  ( n7574 ) ? ( VREG_16_4 ) : ( n8094 ) ;
assign n8096 =  ( n7573 ) ? ( VREG_16_5 ) : ( n8095 ) ;
assign n8097 =  ( n7572 ) ? ( VREG_16_6 ) : ( n8096 ) ;
assign n8098 =  ( n7571 ) ? ( VREG_16_7 ) : ( n8097 ) ;
assign n8099 =  ( n7570 ) ? ( VREG_16_8 ) : ( n8098 ) ;
assign n8100 =  ( n7569 ) ? ( VREG_16_9 ) : ( n8099 ) ;
assign n8101 =  ( n7568 ) ? ( VREG_16_10 ) : ( n8100 ) ;
assign n8102 =  ( n7567 ) ? ( VREG_16_11 ) : ( n8101 ) ;
assign n8103 =  ( n7566 ) ? ( VREG_16_12 ) : ( n8102 ) ;
assign n8104 =  ( n7565 ) ? ( VREG_16_13 ) : ( n8103 ) ;
assign n8105 =  ( n7564 ) ? ( VREG_16_14 ) : ( n8104 ) ;
assign n8106 =  ( n7563 ) ? ( VREG_16_15 ) : ( n8105 ) ;
assign n8107 =  ( n7562 ) ? ( VREG_17_0 ) : ( n8106 ) ;
assign n8108 =  ( n7561 ) ? ( VREG_17_1 ) : ( n8107 ) ;
assign n8109 =  ( n7560 ) ? ( VREG_17_2 ) : ( n8108 ) ;
assign n8110 =  ( n7559 ) ? ( VREG_17_3 ) : ( n8109 ) ;
assign n8111 =  ( n7558 ) ? ( VREG_17_4 ) : ( n8110 ) ;
assign n8112 =  ( n7557 ) ? ( VREG_17_5 ) : ( n8111 ) ;
assign n8113 =  ( n7556 ) ? ( VREG_17_6 ) : ( n8112 ) ;
assign n8114 =  ( n7555 ) ? ( VREG_17_7 ) : ( n8113 ) ;
assign n8115 =  ( n7554 ) ? ( VREG_17_8 ) : ( n8114 ) ;
assign n8116 =  ( n7553 ) ? ( VREG_17_9 ) : ( n8115 ) ;
assign n8117 =  ( n7552 ) ? ( VREG_17_10 ) : ( n8116 ) ;
assign n8118 =  ( n7551 ) ? ( VREG_17_11 ) : ( n8117 ) ;
assign n8119 =  ( n7550 ) ? ( VREG_17_12 ) : ( n8118 ) ;
assign n8120 =  ( n7549 ) ? ( VREG_17_13 ) : ( n8119 ) ;
assign n8121 =  ( n7548 ) ? ( VREG_17_14 ) : ( n8120 ) ;
assign n8122 =  ( n7547 ) ? ( VREG_17_15 ) : ( n8121 ) ;
assign n8123 =  ( n7546 ) ? ( VREG_18_0 ) : ( n8122 ) ;
assign n8124 =  ( n7545 ) ? ( VREG_18_1 ) : ( n8123 ) ;
assign n8125 =  ( n7544 ) ? ( VREG_18_2 ) : ( n8124 ) ;
assign n8126 =  ( n7543 ) ? ( VREG_18_3 ) : ( n8125 ) ;
assign n8127 =  ( n7542 ) ? ( VREG_18_4 ) : ( n8126 ) ;
assign n8128 =  ( n7541 ) ? ( VREG_18_5 ) : ( n8127 ) ;
assign n8129 =  ( n7540 ) ? ( VREG_18_6 ) : ( n8128 ) ;
assign n8130 =  ( n7539 ) ? ( VREG_18_7 ) : ( n8129 ) ;
assign n8131 =  ( n7538 ) ? ( VREG_18_8 ) : ( n8130 ) ;
assign n8132 =  ( n7537 ) ? ( VREG_18_9 ) : ( n8131 ) ;
assign n8133 =  ( n7536 ) ? ( VREG_18_10 ) : ( n8132 ) ;
assign n8134 =  ( n7535 ) ? ( VREG_18_11 ) : ( n8133 ) ;
assign n8135 =  ( n7534 ) ? ( VREG_18_12 ) : ( n8134 ) ;
assign n8136 =  ( n7533 ) ? ( VREG_18_13 ) : ( n8135 ) ;
assign n8137 =  ( n7532 ) ? ( VREG_18_14 ) : ( n8136 ) ;
assign n8138 =  ( n7531 ) ? ( VREG_18_15 ) : ( n8137 ) ;
assign n8139 =  ( n7530 ) ? ( VREG_19_0 ) : ( n8138 ) ;
assign n8140 =  ( n7529 ) ? ( VREG_19_1 ) : ( n8139 ) ;
assign n8141 =  ( n7528 ) ? ( VREG_19_2 ) : ( n8140 ) ;
assign n8142 =  ( n7527 ) ? ( VREG_19_3 ) : ( n8141 ) ;
assign n8143 =  ( n7526 ) ? ( VREG_19_4 ) : ( n8142 ) ;
assign n8144 =  ( n7525 ) ? ( VREG_19_5 ) : ( n8143 ) ;
assign n8145 =  ( n7524 ) ? ( VREG_19_6 ) : ( n8144 ) ;
assign n8146 =  ( n7523 ) ? ( VREG_19_7 ) : ( n8145 ) ;
assign n8147 =  ( n7522 ) ? ( VREG_19_8 ) : ( n8146 ) ;
assign n8148 =  ( n7521 ) ? ( VREG_19_9 ) : ( n8147 ) ;
assign n8149 =  ( n7520 ) ? ( VREG_19_10 ) : ( n8148 ) ;
assign n8150 =  ( n7519 ) ? ( VREG_19_11 ) : ( n8149 ) ;
assign n8151 =  ( n7518 ) ? ( VREG_19_12 ) : ( n8150 ) ;
assign n8152 =  ( n7517 ) ? ( VREG_19_13 ) : ( n8151 ) ;
assign n8153 =  ( n7516 ) ? ( VREG_19_14 ) : ( n8152 ) ;
assign n8154 =  ( n7515 ) ? ( VREG_19_15 ) : ( n8153 ) ;
assign n8155 =  ( n7514 ) ? ( VREG_20_0 ) : ( n8154 ) ;
assign n8156 =  ( n7513 ) ? ( VREG_20_1 ) : ( n8155 ) ;
assign n8157 =  ( n7512 ) ? ( VREG_20_2 ) : ( n8156 ) ;
assign n8158 =  ( n7511 ) ? ( VREG_20_3 ) : ( n8157 ) ;
assign n8159 =  ( n7510 ) ? ( VREG_20_4 ) : ( n8158 ) ;
assign n8160 =  ( n7509 ) ? ( VREG_20_5 ) : ( n8159 ) ;
assign n8161 =  ( n7508 ) ? ( VREG_20_6 ) : ( n8160 ) ;
assign n8162 =  ( n7507 ) ? ( VREG_20_7 ) : ( n8161 ) ;
assign n8163 =  ( n7506 ) ? ( VREG_20_8 ) : ( n8162 ) ;
assign n8164 =  ( n7505 ) ? ( VREG_20_9 ) : ( n8163 ) ;
assign n8165 =  ( n7504 ) ? ( VREG_20_10 ) : ( n8164 ) ;
assign n8166 =  ( n7503 ) ? ( VREG_20_11 ) : ( n8165 ) ;
assign n8167 =  ( n7502 ) ? ( VREG_20_12 ) : ( n8166 ) ;
assign n8168 =  ( n7501 ) ? ( VREG_20_13 ) : ( n8167 ) ;
assign n8169 =  ( n7500 ) ? ( VREG_20_14 ) : ( n8168 ) ;
assign n8170 =  ( n7499 ) ? ( VREG_20_15 ) : ( n8169 ) ;
assign n8171 =  ( n7498 ) ? ( VREG_21_0 ) : ( n8170 ) ;
assign n8172 =  ( n7497 ) ? ( VREG_21_1 ) : ( n8171 ) ;
assign n8173 =  ( n7496 ) ? ( VREG_21_2 ) : ( n8172 ) ;
assign n8174 =  ( n7495 ) ? ( VREG_21_3 ) : ( n8173 ) ;
assign n8175 =  ( n7494 ) ? ( VREG_21_4 ) : ( n8174 ) ;
assign n8176 =  ( n7493 ) ? ( VREG_21_5 ) : ( n8175 ) ;
assign n8177 =  ( n7492 ) ? ( VREG_21_6 ) : ( n8176 ) ;
assign n8178 =  ( n7491 ) ? ( VREG_21_7 ) : ( n8177 ) ;
assign n8179 =  ( n7490 ) ? ( VREG_21_8 ) : ( n8178 ) ;
assign n8180 =  ( n7489 ) ? ( VREG_21_9 ) : ( n8179 ) ;
assign n8181 =  ( n7488 ) ? ( VREG_21_10 ) : ( n8180 ) ;
assign n8182 =  ( n7487 ) ? ( VREG_21_11 ) : ( n8181 ) ;
assign n8183 =  ( n7486 ) ? ( VREG_21_12 ) : ( n8182 ) ;
assign n8184 =  ( n7485 ) ? ( VREG_21_13 ) : ( n8183 ) ;
assign n8185 =  ( n7484 ) ? ( VREG_21_14 ) : ( n8184 ) ;
assign n8186 =  ( n7483 ) ? ( VREG_21_15 ) : ( n8185 ) ;
assign n8187 =  ( n7482 ) ? ( VREG_22_0 ) : ( n8186 ) ;
assign n8188 =  ( n7481 ) ? ( VREG_22_1 ) : ( n8187 ) ;
assign n8189 =  ( n7480 ) ? ( VREG_22_2 ) : ( n8188 ) ;
assign n8190 =  ( n7479 ) ? ( VREG_22_3 ) : ( n8189 ) ;
assign n8191 =  ( n7478 ) ? ( VREG_22_4 ) : ( n8190 ) ;
assign n8192 =  ( n7477 ) ? ( VREG_22_5 ) : ( n8191 ) ;
assign n8193 =  ( n7476 ) ? ( VREG_22_6 ) : ( n8192 ) ;
assign n8194 =  ( n7475 ) ? ( VREG_22_7 ) : ( n8193 ) ;
assign n8195 =  ( n7474 ) ? ( VREG_22_8 ) : ( n8194 ) ;
assign n8196 =  ( n7473 ) ? ( VREG_22_9 ) : ( n8195 ) ;
assign n8197 =  ( n7472 ) ? ( VREG_22_10 ) : ( n8196 ) ;
assign n8198 =  ( n7471 ) ? ( VREG_22_11 ) : ( n8197 ) ;
assign n8199 =  ( n7470 ) ? ( VREG_22_12 ) : ( n8198 ) ;
assign n8200 =  ( n7469 ) ? ( VREG_22_13 ) : ( n8199 ) ;
assign n8201 =  ( n7468 ) ? ( VREG_22_14 ) : ( n8200 ) ;
assign n8202 =  ( n7467 ) ? ( VREG_22_15 ) : ( n8201 ) ;
assign n8203 =  ( n7466 ) ? ( VREG_23_0 ) : ( n8202 ) ;
assign n8204 =  ( n7465 ) ? ( VREG_23_1 ) : ( n8203 ) ;
assign n8205 =  ( n7464 ) ? ( VREG_23_2 ) : ( n8204 ) ;
assign n8206 =  ( n7463 ) ? ( VREG_23_3 ) : ( n8205 ) ;
assign n8207 =  ( n7462 ) ? ( VREG_23_4 ) : ( n8206 ) ;
assign n8208 =  ( n7461 ) ? ( VREG_23_5 ) : ( n8207 ) ;
assign n8209 =  ( n7460 ) ? ( VREG_23_6 ) : ( n8208 ) ;
assign n8210 =  ( n7459 ) ? ( VREG_23_7 ) : ( n8209 ) ;
assign n8211 =  ( n7458 ) ? ( VREG_23_8 ) : ( n8210 ) ;
assign n8212 =  ( n7457 ) ? ( VREG_23_9 ) : ( n8211 ) ;
assign n8213 =  ( n7456 ) ? ( VREG_23_10 ) : ( n8212 ) ;
assign n8214 =  ( n7455 ) ? ( VREG_23_11 ) : ( n8213 ) ;
assign n8215 =  ( n7454 ) ? ( VREG_23_12 ) : ( n8214 ) ;
assign n8216 =  ( n7453 ) ? ( VREG_23_13 ) : ( n8215 ) ;
assign n8217 =  ( n7452 ) ? ( VREG_23_14 ) : ( n8216 ) ;
assign n8218 =  ( n7451 ) ? ( VREG_23_15 ) : ( n8217 ) ;
assign n8219 =  ( n7450 ) ? ( VREG_24_0 ) : ( n8218 ) ;
assign n8220 =  ( n7449 ) ? ( VREG_24_1 ) : ( n8219 ) ;
assign n8221 =  ( n7448 ) ? ( VREG_24_2 ) : ( n8220 ) ;
assign n8222 =  ( n7447 ) ? ( VREG_24_3 ) : ( n8221 ) ;
assign n8223 =  ( n7446 ) ? ( VREG_24_4 ) : ( n8222 ) ;
assign n8224 =  ( n7445 ) ? ( VREG_24_5 ) : ( n8223 ) ;
assign n8225 =  ( n7444 ) ? ( VREG_24_6 ) : ( n8224 ) ;
assign n8226 =  ( n7443 ) ? ( VREG_24_7 ) : ( n8225 ) ;
assign n8227 =  ( n7442 ) ? ( VREG_24_8 ) : ( n8226 ) ;
assign n8228 =  ( n7441 ) ? ( VREG_24_9 ) : ( n8227 ) ;
assign n8229 =  ( n7440 ) ? ( VREG_24_10 ) : ( n8228 ) ;
assign n8230 =  ( n7439 ) ? ( VREG_24_11 ) : ( n8229 ) ;
assign n8231 =  ( n7438 ) ? ( VREG_24_12 ) : ( n8230 ) ;
assign n8232 =  ( n7437 ) ? ( VREG_24_13 ) : ( n8231 ) ;
assign n8233 =  ( n7436 ) ? ( VREG_24_14 ) : ( n8232 ) ;
assign n8234 =  ( n7435 ) ? ( VREG_24_15 ) : ( n8233 ) ;
assign n8235 =  ( n7434 ) ? ( VREG_25_0 ) : ( n8234 ) ;
assign n8236 =  ( n7433 ) ? ( VREG_25_1 ) : ( n8235 ) ;
assign n8237 =  ( n7432 ) ? ( VREG_25_2 ) : ( n8236 ) ;
assign n8238 =  ( n7431 ) ? ( VREG_25_3 ) : ( n8237 ) ;
assign n8239 =  ( n7430 ) ? ( VREG_25_4 ) : ( n8238 ) ;
assign n8240 =  ( n7429 ) ? ( VREG_25_5 ) : ( n8239 ) ;
assign n8241 =  ( n7428 ) ? ( VREG_25_6 ) : ( n8240 ) ;
assign n8242 =  ( n7427 ) ? ( VREG_25_7 ) : ( n8241 ) ;
assign n8243 =  ( n7426 ) ? ( VREG_25_8 ) : ( n8242 ) ;
assign n8244 =  ( n7425 ) ? ( VREG_25_9 ) : ( n8243 ) ;
assign n8245 =  ( n7424 ) ? ( VREG_25_10 ) : ( n8244 ) ;
assign n8246 =  ( n7423 ) ? ( VREG_25_11 ) : ( n8245 ) ;
assign n8247 =  ( n7422 ) ? ( VREG_25_12 ) : ( n8246 ) ;
assign n8248 =  ( n7421 ) ? ( VREG_25_13 ) : ( n8247 ) ;
assign n8249 =  ( n7420 ) ? ( VREG_25_14 ) : ( n8248 ) ;
assign n8250 =  ( n7419 ) ? ( VREG_25_15 ) : ( n8249 ) ;
assign n8251 =  ( n7418 ) ? ( VREG_26_0 ) : ( n8250 ) ;
assign n8252 =  ( n7417 ) ? ( VREG_26_1 ) : ( n8251 ) ;
assign n8253 =  ( n7416 ) ? ( VREG_26_2 ) : ( n8252 ) ;
assign n8254 =  ( n7415 ) ? ( VREG_26_3 ) : ( n8253 ) ;
assign n8255 =  ( n7414 ) ? ( VREG_26_4 ) : ( n8254 ) ;
assign n8256 =  ( n7413 ) ? ( VREG_26_5 ) : ( n8255 ) ;
assign n8257 =  ( n7412 ) ? ( VREG_26_6 ) : ( n8256 ) ;
assign n8258 =  ( n7411 ) ? ( VREG_26_7 ) : ( n8257 ) ;
assign n8259 =  ( n7410 ) ? ( VREG_26_8 ) : ( n8258 ) ;
assign n8260 =  ( n7409 ) ? ( VREG_26_9 ) : ( n8259 ) ;
assign n8261 =  ( n7408 ) ? ( VREG_26_10 ) : ( n8260 ) ;
assign n8262 =  ( n7407 ) ? ( VREG_26_11 ) : ( n8261 ) ;
assign n8263 =  ( n7406 ) ? ( VREG_26_12 ) : ( n8262 ) ;
assign n8264 =  ( n7405 ) ? ( VREG_26_13 ) : ( n8263 ) ;
assign n8265 =  ( n7404 ) ? ( VREG_26_14 ) : ( n8264 ) ;
assign n8266 =  ( n7403 ) ? ( VREG_26_15 ) : ( n8265 ) ;
assign n8267 =  ( n7402 ) ? ( VREG_27_0 ) : ( n8266 ) ;
assign n8268 =  ( n7401 ) ? ( VREG_27_1 ) : ( n8267 ) ;
assign n8269 =  ( n7400 ) ? ( VREG_27_2 ) : ( n8268 ) ;
assign n8270 =  ( n7399 ) ? ( VREG_27_3 ) : ( n8269 ) ;
assign n8271 =  ( n7398 ) ? ( VREG_27_4 ) : ( n8270 ) ;
assign n8272 =  ( n7397 ) ? ( VREG_27_5 ) : ( n8271 ) ;
assign n8273 =  ( n7396 ) ? ( VREG_27_6 ) : ( n8272 ) ;
assign n8274 =  ( n7395 ) ? ( VREG_27_7 ) : ( n8273 ) ;
assign n8275 =  ( n7394 ) ? ( VREG_27_8 ) : ( n8274 ) ;
assign n8276 =  ( n7393 ) ? ( VREG_27_9 ) : ( n8275 ) ;
assign n8277 =  ( n7392 ) ? ( VREG_27_10 ) : ( n8276 ) ;
assign n8278 =  ( n7391 ) ? ( VREG_27_11 ) : ( n8277 ) ;
assign n8279 =  ( n7390 ) ? ( VREG_27_12 ) : ( n8278 ) ;
assign n8280 =  ( n7389 ) ? ( VREG_27_13 ) : ( n8279 ) ;
assign n8281 =  ( n7388 ) ? ( VREG_27_14 ) : ( n8280 ) ;
assign n8282 =  ( n7387 ) ? ( VREG_27_15 ) : ( n8281 ) ;
assign n8283 =  ( n7386 ) ? ( VREG_28_0 ) : ( n8282 ) ;
assign n8284 =  ( n7385 ) ? ( VREG_28_1 ) : ( n8283 ) ;
assign n8285 =  ( n7384 ) ? ( VREG_28_2 ) : ( n8284 ) ;
assign n8286 =  ( n7383 ) ? ( VREG_28_3 ) : ( n8285 ) ;
assign n8287 =  ( n7382 ) ? ( VREG_28_4 ) : ( n8286 ) ;
assign n8288 =  ( n7381 ) ? ( VREG_28_5 ) : ( n8287 ) ;
assign n8289 =  ( n7380 ) ? ( VREG_28_6 ) : ( n8288 ) ;
assign n8290 =  ( n7379 ) ? ( VREG_28_7 ) : ( n8289 ) ;
assign n8291 =  ( n7378 ) ? ( VREG_28_8 ) : ( n8290 ) ;
assign n8292 =  ( n7377 ) ? ( VREG_28_9 ) : ( n8291 ) ;
assign n8293 =  ( n7376 ) ? ( VREG_28_10 ) : ( n8292 ) ;
assign n8294 =  ( n7375 ) ? ( VREG_28_11 ) : ( n8293 ) ;
assign n8295 =  ( n7374 ) ? ( VREG_28_12 ) : ( n8294 ) ;
assign n8296 =  ( n7373 ) ? ( VREG_28_13 ) : ( n8295 ) ;
assign n8297 =  ( n7372 ) ? ( VREG_28_14 ) : ( n8296 ) ;
assign n8298 =  ( n7371 ) ? ( VREG_28_15 ) : ( n8297 ) ;
assign n8299 =  ( n7370 ) ? ( VREG_29_0 ) : ( n8298 ) ;
assign n8300 =  ( n7369 ) ? ( VREG_29_1 ) : ( n8299 ) ;
assign n8301 =  ( n7368 ) ? ( VREG_29_2 ) : ( n8300 ) ;
assign n8302 =  ( n7367 ) ? ( VREG_29_3 ) : ( n8301 ) ;
assign n8303 =  ( n7366 ) ? ( VREG_29_4 ) : ( n8302 ) ;
assign n8304 =  ( n7365 ) ? ( VREG_29_5 ) : ( n8303 ) ;
assign n8305 =  ( n7364 ) ? ( VREG_29_6 ) : ( n8304 ) ;
assign n8306 =  ( n7363 ) ? ( VREG_29_7 ) : ( n8305 ) ;
assign n8307 =  ( n7362 ) ? ( VREG_29_8 ) : ( n8306 ) ;
assign n8308 =  ( n7361 ) ? ( VREG_29_9 ) : ( n8307 ) ;
assign n8309 =  ( n7360 ) ? ( VREG_29_10 ) : ( n8308 ) ;
assign n8310 =  ( n7359 ) ? ( VREG_29_11 ) : ( n8309 ) ;
assign n8311 =  ( n7358 ) ? ( VREG_29_12 ) : ( n8310 ) ;
assign n8312 =  ( n7357 ) ? ( VREG_29_13 ) : ( n8311 ) ;
assign n8313 =  ( n7356 ) ? ( VREG_29_14 ) : ( n8312 ) ;
assign n8314 =  ( n7355 ) ? ( VREG_29_15 ) : ( n8313 ) ;
assign n8315 =  ( n7354 ) ? ( VREG_30_0 ) : ( n8314 ) ;
assign n8316 =  ( n7353 ) ? ( VREG_30_1 ) : ( n8315 ) ;
assign n8317 =  ( n7352 ) ? ( VREG_30_2 ) : ( n8316 ) ;
assign n8318 =  ( n7351 ) ? ( VREG_30_3 ) : ( n8317 ) ;
assign n8319 =  ( n7350 ) ? ( VREG_30_4 ) : ( n8318 ) ;
assign n8320 =  ( n7349 ) ? ( VREG_30_5 ) : ( n8319 ) ;
assign n8321 =  ( n7348 ) ? ( VREG_30_6 ) : ( n8320 ) ;
assign n8322 =  ( n7347 ) ? ( VREG_30_7 ) : ( n8321 ) ;
assign n8323 =  ( n7346 ) ? ( VREG_30_8 ) : ( n8322 ) ;
assign n8324 =  ( n7345 ) ? ( VREG_30_9 ) : ( n8323 ) ;
assign n8325 =  ( n7344 ) ? ( VREG_30_10 ) : ( n8324 ) ;
assign n8326 =  ( n7343 ) ? ( VREG_30_11 ) : ( n8325 ) ;
assign n8327 =  ( n7342 ) ? ( VREG_30_12 ) : ( n8326 ) ;
assign n8328 =  ( n7341 ) ? ( VREG_30_13 ) : ( n8327 ) ;
assign n8329 =  ( n7340 ) ? ( VREG_30_14 ) : ( n8328 ) ;
assign n8330 =  ( n7339 ) ? ( VREG_30_15 ) : ( n8329 ) ;
assign n8331 =  ( n7338 ) ? ( VREG_31_0 ) : ( n8330 ) ;
assign n8332 =  ( n7336 ) ? ( VREG_31_1 ) : ( n8331 ) ;
assign n8333 =  ( n7334 ) ? ( VREG_31_2 ) : ( n8332 ) ;
assign n8334 =  ( n7332 ) ? ( VREG_31_3 ) : ( n8333 ) ;
assign n8335 =  ( n7330 ) ? ( VREG_31_4 ) : ( n8334 ) ;
assign n8336 =  ( n7328 ) ? ( VREG_31_5 ) : ( n8335 ) ;
assign n8337 =  ( n7326 ) ? ( VREG_31_6 ) : ( n8336 ) ;
assign n8338 =  ( n7324 ) ? ( VREG_31_7 ) : ( n8337 ) ;
assign n8339 =  ( n7322 ) ? ( VREG_31_8 ) : ( n8338 ) ;
assign n8340 =  ( n7320 ) ? ( VREG_31_9 ) : ( n8339 ) ;
assign n8341 =  ( n7318 ) ? ( VREG_31_10 ) : ( n8340 ) ;
assign n8342 =  ( n7316 ) ? ( VREG_31_11 ) : ( n8341 ) ;
assign n8343 =  ( n7314 ) ? ( VREG_31_12 ) : ( n8342 ) ;
assign n8344 =  ( n7312 ) ? ( VREG_31_13 ) : ( n8343 ) ;
assign n8345 =  ( n7310 ) ? ( VREG_31_14 ) : ( n8344 ) ;
assign n8346 =  ( n7308 ) ? ( VREG_31_15 ) : ( n8345 ) ;
assign n8347 =  ( n8346 ) + ( n140 )  ;
assign n8348 =  ( n8346 ) - ( n140 )  ;
assign n8349 =  ( n8346 ) & ( n140 )  ;
assign n8350 =  ( n8346 ) | ( n140 )  ;
assign n8351 =  ( ( n8346 ) * ( n140 ))  ;
assign n8352 =  ( n148 ) ? ( n8351 ) : ( VREG_0_11 ) ;
assign n8353 =  ( n146 ) ? ( n8350 ) : ( n8352 ) ;
assign n8354 =  ( n144 ) ? ( n8349 ) : ( n8353 ) ;
assign n8355 =  ( n142 ) ? ( n8348 ) : ( n8354 ) ;
assign n8356 =  ( n10 ) ? ( n8347 ) : ( n8355 ) ;
assign n8357 =  ( n77 ) & ( n7307 )  ;
assign n8358 =  ( n77 ) & ( n7309 )  ;
assign n8359 =  ( n77 ) & ( n7311 )  ;
assign n8360 =  ( n77 ) & ( n7313 )  ;
assign n8361 =  ( n77 ) & ( n7315 )  ;
assign n8362 =  ( n77 ) & ( n7317 )  ;
assign n8363 =  ( n77 ) & ( n7319 )  ;
assign n8364 =  ( n77 ) & ( n7321 )  ;
assign n8365 =  ( n77 ) & ( n7323 )  ;
assign n8366 =  ( n77 ) & ( n7325 )  ;
assign n8367 =  ( n77 ) & ( n7327 )  ;
assign n8368 =  ( n77 ) & ( n7329 )  ;
assign n8369 =  ( n77 ) & ( n7331 )  ;
assign n8370 =  ( n77 ) & ( n7333 )  ;
assign n8371 =  ( n77 ) & ( n7335 )  ;
assign n8372 =  ( n77 ) & ( n7337 )  ;
assign n8373 =  ( n78 ) & ( n7307 )  ;
assign n8374 =  ( n78 ) & ( n7309 )  ;
assign n8375 =  ( n78 ) & ( n7311 )  ;
assign n8376 =  ( n78 ) & ( n7313 )  ;
assign n8377 =  ( n78 ) & ( n7315 )  ;
assign n8378 =  ( n78 ) & ( n7317 )  ;
assign n8379 =  ( n78 ) & ( n7319 )  ;
assign n8380 =  ( n78 ) & ( n7321 )  ;
assign n8381 =  ( n78 ) & ( n7323 )  ;
assign n8382 =  ( n78 ) & ( n7325 )  ;
assign n8383 =  ( n78 ) & ( n7327 )  ;
assign n8384 =  ( n78 ) & ( n7329 )  ;
assign n8385 =  ( n78 ) & ( n7331 )  ;
assign n8386 =  ( n78 ) & ( n7333 )  ;
assign n8387 =  ( n78 ) & ( n7335 )  ;
assign n8388 =  ( n78 ) & ( n7337 )  ;
assign n8389 =  ( n79 ) & ( n7307 )  ;
assign n8390 =  ( n79 ) & ( n7309 )  ;
assign n8391 =  ( n79 ) & ( n7311 )  ;
assign n8392 =  ( n79 ) & ( n7313 )  ;
assign n8393 =  ( n79 ) & ( n7315 )  ;
assign n8394 =  ( n79 ) & ( n7317 )  ;
assign n8395 =  ( n79 ) & ( n7319 )  ;
assign n8396 =  ( n79 ) & ( n7321 )  ;
assign n8397 =  ( n79 ) & ( n7323 )  ;
assign n8398 =  ( n79 ) & ( n7325 )  ;
assign n8399 =  ( n79 ) & ( n7327 )  ;
assign n8400 =  ( n79 ) & ( n7329 )  ;
assign n8401 =  ( n79 ) & ( n7331 )  ;
assign n8402 =  ( n79 ) & ( n7333 )  ;
assign n8403 =  ( n79 ) & ( n7335 )  ;
assign n8404 =  ( n79 ) & ( n7337 )  ;
assign n8405 =  ( n80 ) & ( n7307 )  ;
assign n8406 =  ( n80 ) & ( n7309 )  ;
assign n8407 =  ( n80 ) & ( n7311 )  ;
assign n8408 =  ( n80 ) & ( n7313 )  ;
assign n8409 =  ( n80 ) & ( n7315 )  ;
assign n8410 =  ( n80 ) & ( n7317 )  ;
assign n8411 =  ( n80 ) & ( n7319 )  ;
assign n8412 =  ( n80 ) & ( n7321 )  ;
assign n8413 =  ( n80 ) & ( n7323 )  ;
assign n8414 =  ( n80 ) & ( n7325 )  ;
assign n8415 =  ( n80 ) & ( n7327 )  ;
assign n8416 =  ( n80 ) & ( n7329 )  ;
assign n8417 =  ( n80 ) & ( n7331 )  ;
assign n8418 =  ( n80 ) & ( n7333 )  ;
assign n8419 =  ( n80 ) & ( n7335 )  ;
assign n8420 =  ( n80 ) & ( n7337 )  ;
assign n8421 =  ( n81 ) & ( n7307 )  ;
assign n8422 =  ( n81 ) & ( n7309 )  ;
assign n8423 =  ( n81 ) & ( n7311 )  ;
assign n8424 =  ( n81 ) & ( n7313 )  ;
assign n8425 =  ( n81 ) & ( n7315 )  ;
assign n8426 =  ( n81 ) & ( n7317 )  ;
assign n8427 =  ( n81 ) & ( n7319 )  ;
assign n8428 =  ( n81 ) & ( n7321 )  ;
assign n8429 =  ( n81 ) & ( n7323 )  ;
assign n8430 =  ( n81 ) & ( n7325 )  ;
assign n8431 =  ( n81 ) & ( n7327 )  ;
assign n8432 =  ( n81 ) & ( n7329 )  ;
assign n8433 =  ( n81 ) & ( n7331 )  ;
assign n8434 =  ( n81 ) & ( n7333 )  ;
assign n8435 =  ( n81 ) & ( n7335 )  ;
assign n8436 =  ( n81 ) & ( n7337 )  ;
assign n8437 =  ( n82 ) & ( n7307 )  ;
assign n8438 =  ( n82 ) & ( n7309 )  ;
assign n8439 =  ( n82 ) & ( n7311 )  ;
assign n8440 =  ( n82 ) & ( n7313 )  ;
assign n8441 =  ( n82 ) & ( n7315 )  ;
assign n8442 =  ( n82 ) & ( n7317 )  ;
assign n8443 =  ( n82 ) & ( n7319 )  ;
assign n8444 =  ( n82 ) & ( n7321 )  ;
assign n8445 =  ( n82 ) & ( n7323 )  ;
assign n8446 =  ( n82 ) & ( n7325 )  ;
assign n8447 =  ( n82 ) & ( n7327 )  ;
assign n8448 =  ( n82 ) & ( n7329 )  ;
assign n8449 =  ( n82 ) & ( n7331 )  ;
assign n8450 =  ( n82 ) & ( n7333 )  ;
assign n8451 =  ( n82 ) & ( n7335 )  ;
assign n8452 =  ( n82 ) & ( n7337 )  ;
assign n8453 =  ( n83 ) & ( n7307 )  ;
assign n8454 =  ( n83 ) & ( n7309 )  ;
assign n8455 =  ( n83 ) & ( n7311 )  ;
assign n8456 =  ( n83 ) & ( n7313 )  ;
assign n8457 =  ( n83 ) & ( n7315 )  ;
assign n8458 =  ( n83 ) & ( n7317 )  ;
assign n8459 =  ( n83 ) & ( n7319 )  ;
assign n8460 =  ( n83 ) & ( n7321 )  ;
assign n8461 =  ( n83 ) & ( n7323 )  ;
assign n8462 =  ( n83 ) & ( n7325 )  ;
assign n8463 =  ( n83 ) & ( n7327 )  ;
assign n8464 =  ( n83 ) & ( n7329 )  ;
assign n8465 =  ( n83 ) & ( n7331 )  ;
assign n8466 =  ( n83 ) & ( n7333 )  ;
assign n8467 =  ( n83 ) & ( n7335 )  ;
assign n8468 =  ( n83 ) & ( n7337 )  ;
assign n8469 =  ( n84 ) & ( n7307 )  ;
assign n8470 =  ( n84 ) & ( n7309 )  ;
assign n8471 =  ( n84 ) & ( n7311 )  ;
assign n8472 =  ( n84 ) & ( n7313 )  ;
assign n8473 =  ( n84 ) & ( n7315 )  ;
assign n8474 =  ( n84 ) & ( n7317 )  ;
assign n8475 =  ( n84 ) & ( n7319 )  ;
assign n8476 =  ( n84 ) & ( n7321 )  ;
assign n8477 =  ( n84 ) & ( n7323 )  ;
assign n8478 =  ( n84 ) & ( n7325 )  ;
assign n8479 =  ( n84 ) & ( n7327 )  ;
assign n8480 =  ( n84 ) & ( n7329 )  ;
assign n8481 =  ( n84 ) & ( n7331 )  ;
assign n8482 =  ( n84 ) & ( n7333 )  ;
assign n8483 =  ( n84 ) & ( n7335 )  ;
assign n8484 =  ( n84 ) & ( n7337 )  ;
assign n8485 =  ( n85 ) & ( n7307 )  ;
assign n8486 =  ( n85 ) & ( n7309 )  ;
assign n8487 =  ( n85 ) & ( n7311 )  ;
assign n8488 =  ( n85 ) & ( n7313 )  ;
assign n8489 =  ( n85 ) & ( n7315 )  ;
assign n8490 =  ( n85 ) & ( n7317 )  ;
assign n8491 =  ( n85 ) & ( n7319 )  ;
assign n8492 =  ( n85 ) & ( n7321 )  ;
assign n8493 =  ( n85 ) & ( n7323 )  ;
assign n8494 =  ( n85 ) & ( n7325 )  ;
assign n8495 =  ( n85 ) & ( n7327 )  ;
assign n8496 =  ( n85 ) & ( n7329 )  ;
assign n8497 =  ( n85 ) & ( n7331 )  ;
assign n8498 =  ( n85 ) & ( n7333 )  ;
assign n8499 =  ( n85 ) & ( n7335 )  ;
assign n8500 =  ( n85 ) & ( n7337 )  ;
assign n8501 =  ( n86 ) & ( n7307 )  ;
assign n8502 =  ( n86 ) & ( n7309 )  ;
assign n8503 =  ( n86 ) & ( n7311 )  ;
assign n8504 =  ( n86 ) & ( n7313 )  ;
assign n8505 =  ( n86 ) & ( n7315 )  ;
assign n8506 =  ( n86 ) & ( n7317 )  ;
assign n8507 =  ( n86 ) & ( n7319 )  ;
assign n8508 =  ( n86 ) & ( n7321 )  ;
assign n8509 =  ( n86 ) & ( n7323 )  ;
assign n8510 =  ( n86 ) & ( n7325 )  ;
assign n8511 =  ( n86 ) & ( n7327 )  ;
assign n8512 =  ( n86 ) & ( n7329 )  ;
assign n8513 =  ( n86 ) & ( n7331 )  ;
assign n8514 =  ( n86 ) & ( n7333 )  ;
assign n8515 =  ( n86 ) & ( n7335 )  ;
assign n8516 =  ( n86 ) & ( n7337 )  ;
assign n8517 =  ( n87 ) & ( n7307 )  ;
assign n8518 =  ( n87 ) & ( n7309 )  ;
assign n8519 =  ( n87 ) & ( n7311 )  ;
assign n8520 =  ( n87 ) & ( n7313 )  ;
assign n8521 =  ( n87 ) & ( n7315 )  ;
assign n8522 =  ( n87 ) & ( n7317 )  ;
assign n8523 =  ( n87 ) & ( n7319 )  ;
assign n8524 =  ( n87 ) & ( n7321 )  ;
assign n8525 =  ( n87 ) & ( n7323 )  ;
assign n8526 =  ( n87 ) & ( n7325 )  ;
assign n8527 =  ( n87 ) & ( n7327 )  ;
assign n8528 =  ( n87 ) & ( n7329 )  ;
assign n8529 =  ( n87 ) & ( n7331 )  ;
assign n8530 =  ( n87 ) & ( n7333 )  ;
assign n8531 =  ( n87 ) & ( n7335 )  ;
assign n8532 =  ( n87 ) & ( n7337 )  ;
assign n8533 =  ( n88 ) & ( n7307 )  ;
assign n8534 =  ( n88 ) & ( n7309 )  ;
assign n8535 =  ( n88 ) & ( n7311 )  ;
assign n8536 =  ( n88 ) & ( n7313 )  ;
assign n8537 =  ( n88 ) & ( n7315 )  ;
assign n8538 =  ( n88 ) & ( n7317 )  ;
assign n8539 =  ( n88 ) & ( n7319 )  ;
assign n8540 =  ( n88 ) & ( n7321 )  ;
assign n8541 =  ( n88 ) & ( n7323 )  ;
assign n8542 =  ( n88 ) & ( n7325 )  ;
assign n8543 =  ( n88 ) & ( n7327 )  ;
assign n8544 =  ( n88 ) & ( n7329 )  ;
assign n8545 =  ( n88 ) & ( n7331 )  ;
assign n8546 =  ( n88 ) & ( n7333 )  ;
assign n8547 =  ( n88 ) & ( n7335 )  ;
assign n8548 =  ( n88 ) & ( n7337 )  ;
assign n8549 =  ( n89 ) & ( n7307 )  ;
assign n8550 =  ( n89 ) & ( n7309 )  ;
assign n8551 =  ( n89 ) & ( n7311 )  ;
assign n8552 =  ( n89 ) & ( n7313 )  ;
assign n8553 =  ( n89 ) & ( n7315 )  ;
assign n8554 =  ( n89 ) & ( n7317 )  ;
assign n8555 =  ( n89 ) & ( n7319 )  ;
assign n8556 =  ( n89 ) & ( n7321 )  ;
assign n8557 =  ( n89 ) & ( n7323 )  ;
assign n8558 =  ( n89 ) & ( n7325 )  ;
assign n8559 =  ( n89 ) & ( n7327 )  ;
assign n8560 =  ( n89 ) & ( n7329 )  ;
assign n8561 =  ( n89 ) & ( n7331 )  ;
assign n8562 =  ( n89 ) & ( n7333 )  ;
assign n8563 =  ( n89 ) & ( n7335 )  ;
assign n8564 =  ( n89 ) & ( n7337 )  ;
assign n8565 =  ( n90 ) & ( n7307 )  ;
assign n8566 =  ( n90 ) & ( n7309 )  ;
assign n8567 =  ( n90 ) & ( n7311 )  ;
assign n8568 =  ( n90 ) & ( n7313 )  ;
assign n8569 =  ( n90 ) & ( n7315 )  ;
assign n8570 =  ( n90 ) & ( n7317 )  ;
assign n8571 =  ( n90 ) & ( n7319 )  ;
assign n8572 =  ( n90 ) & ( n7321 )  ;
assign n8573 =  ( n90 ) & ( n7323 )  ;
assign n8574 =  ( n90 ) & ( n7325 )  ;
assign n8575 =  ( n90 ) & ( n7327 )  ;
assign n8576 =  ( n90 ) & ( n7329 )  ;
assign n8577 =  ( n90 ) & ( n7331 )  ;
assign n8578 =  ( n90 ) & ( n7333 )  ;
assign n8579 =  ( n90 ) & ( n7335 )  ;
assign n8580 =  ( n90 ) & ( n7337 )  ;
assign n8581 =  ( n91 ) & ( n7307 )  ;
assign n8582 =  ( n91 ) & ( n7309 )  ;
assign n8583 =  ( n91 ) & ( n7311 )  ;
assign n8584 =  ( n91 ) & ( n7313 )  ;
assign n8585 =  ( n91 ) & ( n7315 )  ;
assign n8586 =  ( n91 ) & ( n7317 )  ;
assign n8587 =  ( n91 ) & ( n7319 )  ;
assign n8588 =  ( n91 ) & ( n7321 )  ;
assign n8589 =  ( n91 ) & ( n7323 )  ;
assign n8590 =  ( n91 ) & ( n7325 )  ;
assign n8591 =  ( n91 ) & ( n7327 )  ;
assign n8592 =  ( n91 ) & ( n7329 )  ;
assign n8593 =  ( n91 ) & ( n7331 )  ;
assign n8594 =  ( n91 ) & ( n7333 )  ;
assign n8595 =  ( n91 ) & ( n7335 )  ;
assign n8596 =  ( n91 ) & ( n7337 )  ;
assign n8597 =  ( n92 ) & ( n7307 )  ;
assign n8598 =  ( n92 ) & ( n7309 )  ;
assign n8599 =  ( n92 ) & ( n7311 )  ;
assign n8600 =  ( n92 ) & ( n7313 )  ;
assign n8601 =  ( n92 ) & ( n7315 )  ;
assign n8602 =  ( n92 ) & ( n7317 )  ;
assign n8603 =  ( n92 ) & ( n7319 )  ;
assign n8604 =  ( n92 ) & ( n7321 )  ;
assign n8605 =  ( n92 ) & ( n7323 )  ;
assign n8606 =  ( n92 ) & ( n7325 )  ;
assign n8607 =  ( n92 ) & ( n7327 )  ;
assign n8608 =  ( n92 ) & ( n7329 )  ;
assign n8609 =  ( n92 ) & ( n7331 )  ;
assign n8610 =  ( n92 ) & ( n7333 )  ;
assign n8611 =  ( n92 ) & ( n7335 )  ;
assign n8612 =  ( n92 ) & ( n7337 )  ;
assign n8613 =  ( n93 ) & ( n7307 )  ;
assign n8614 =  ( n93 ) & ( n7309 )  ;
assign n8615 =  ( n93 ) & ( n7311 )  ;
assign n8616 =  ( n93 ) & ( n7313 )  ;
assign n8617 =  ( n93 ) & ( n7315 )  ;
assign n8618 =  ( n93 ) & ( n7317 )  ;
assign n8619 =  ( n93 ) & ( n7319 )  ;
assign n8620 =  ( n93 ) & ( n7321 )  ;
assign n8621 =  ( n93 ) & ( n7323 )  ;
assign n8622 =  ( n93 ) & ( n7325 )  ;
assign n8623 =  ( n93 ) & ( n7327 )  ;
assign n8624 =  ( n93 ) & ( n7329 )  ;
assign n8625 =  ( n93 ) & ( n7331 )  ;
assign n8626 =  ( n93 ) & ( n7333 )  ;
assign n8627 =  ( n93 ) & ( n7335 )  ;
assign n8628 =  ( n93 ) & ( n7337 )  ;
assign n8629 =  ( n94 ) & ( n7307 )  ;
assign n8630 =  ( n94 ) & ( n7309 )  ;
assign n8631 =  ( n94 ) & ( n7311 )  ;
assign n8632 =  ( n94 ) & ( n7313 )  ;
assign n8633 =  ( n94 ) & ( n7315 )  ;
assign n8634 =  ( n94 ) & ( n7317 )  ;
assign n8635 =  ( n94 ) & ( n7319 )  ;
assign n8636 =  ( n94 ) & ( n7321 )  ;
assign n8637 =  ( n94 ) & ( n7323 )  ;
assign n8638 =  ( n94 ) & ( n7325 )  ;
assign n8639 =  ( n94 ) & ( n7327 )  ;
assign n8640 =  ( n94 ) & ( n7329 )  ;
assign n8641 =  ( n94 ) & ( n7331 )  ;
assign n8642 =  ( n94 ) & ( n7333 )  ;
assign n8643 =  ( n94 ) & ( n7335 )  ;
assign n8644 =  ( n94 ) & ( n7337 )  ;
assign n8645 =  ( n95 ) & ( n7307 )  ;
assign n8646 =  ( n95 ) & ( n7309 )  ;
assign n8647 =  ( n95 ) & ( n7311 )  ;
assign n8648 =  ( n95 ) & ( n7313 )  ;
assign n8649 =  ( n95 ) & ( n7315 )  ;
assign n8650 =  ( n95 ) & ( n7317 )  ;
assign n8651 =  ( n95 ) & ( n7319 )  ;
assign n8652 =  ( n95 ) & ( n7321 )  ;
assign n8653 =  ( n95 ) & ( n7323 )  ;
assign n8654 =  ( n95 ) & ( n7325 )  ;
assign n8655 =  ( n95 ) & ( n7327 )  ;
assign n8656 =  ( n95 ) & ( n7329 )  ;
assign n8657 =  ( n95 ) & ( n7331 )  ;
assign n8658 =  ( n95 ) & ( n7333 )  ;
assign n8659 =  ( n95 ) & ( n7335 )  ;
assign n8660 =  ( n95 ) & ( n7337 )  ;
assign n8661 =  ( n96 ) & ( n7307 )  ;
assign n8662 =  ( n96 ) & ( n7309 )  ;
assign n8663 =  ( n96 ) & ( n7311 )  ;
assign n8664 =  ( n96 ) & ( n7313 )  ;
assign n8665 =  ( n96 ) & ( n7315 )  ;
assign n8666 =  ( n96 ) & ( n7317 )  ;
assign n8667 =  ( n96 ) & ( n7319 )  ;
assign n8668 =  ( n96 ) & ( n7321 )  ;
assign n8669 =  ( n96 ) & ( n7323 )  ;
assign n8670 =  ( n96 ) & ( n7325 )  ;
assign n8671 =  ( n96 ) & ( n7327 )  ;
assign n8672 =  ( n96 ) & ( n7329 )  ;
assign n8673 =  ( n96 ) & ( n7331 )  ;
assign n8674 =  ( n96 ) & ( n7333 )  ;
assign n8675 =  ( n96 ) & ( n7335 )  ;
assign n8676 =  ( n96 ) & ( n7337 )  ;
assign n8677 =  ( n97 ) & ( n7307 )  ;
assign n8678 =  ( n97 ) & ( n7309 )  ;
assign n8679 =  ( n97 ) & ( n7311 )  ;
assign n8680 =  ( n97 ) & ( n7313 )  ;
assign n8681 =  ( n97 ) & ( n7315 )  ;
assign n8682 =  ( n97 ) & ( n7317 )  ;
assign n8683 =  ( n97 ) & ( n7319 )  ;
assign n8684 =  ( n97 ) & ( n7321 )  ;
assign n8685 =  ( n97 ) & ( n7323 )  ;
assign n8686 =  ( n97 ) & ( n7325 )  ;
assign n8687 =  ( n97 ) & ( n7327 )  ;
assign n8688 =  ( n97 ) & ( n7329 )  ;
assign n8689 =  ( n97 ) & ( n7331 )  ;
assign n8690 =  ( n97 ) & ( n7333 )  ;
assign n8691 =  ( n97 ) & ( n7335 )  ;
assign n8692 =  ( n97 ) & ( n7337 )  ;
assign n8693 =  ( n98 ) & ( n7307 )  ;
assign n8694 =  ( n98 ) & ( n7309 )  ;
assign n8695 =  ( n98 ) & ( n7311 )  ;
assign n8696 =  ( n98 ) & ( n7313 )  ;
assign n8697 =  ( n98 ) & ( n7315 )  ;
assign n8698 =  ( n98 ) & ( n7317 )  ;
assign n8699 =  ( n98 ) & ( n7319 )  ;
assign n8700 =  ( n98 ) & ( n7321 )  ;
assign n8701 =  ( n98 ) & ( n7323 )  ;
assign n8702 =  ( n98 ) & ( n7325 )  ;
assign n8703 =  ( n98 ) & ( n7327 )  ;
assign n8704 =  ( n98 ) & ( n7329 )  ;
assign n8705 =  ( n98 ) & ( n7331 )  ;
assign n8706 =  ( n98 ) & ( n7333 )  ;
assign n8707 =  ( n98 ) & ( n7335 )  ;
assign n8708 =  ( n98 ) & ( n7337 )  ;
assign n8709 =  ( n99 ) & ( n7307 )  ;
assign n8710 =  ( n99 ) & ( n7309 )  ;
assign n8711 =  ( n99 ) & ( n7311 )  ;
assign n8712 =  ( n99 ) & ( n7313 )  ;
assign n8713 =  ( n99 ) & ( n7315 )  ;
assign n8714 =  ( n99 ) & ( n7317 )  ;
assign n8715 =  ( n99 ) & ( n7319 )  ;
assign n8716 =  ( n99 ) & ( n7321 )  ;
assign n8717 =  ( n99 ) & ( n7323 )  ;
assign n8718 =  ( n99 ) & ( n7325 )  ;
assign n8719 =  ( n99 ) & ( n7327 )  ;
assign n8720 =  ( n99 ) & ( n7329 )  ;
assign n8721 =  ( n99 ) & ( n7331 )  ;
assign n8722 =  ( n99 ) & ( n7333 )  ;
assign n8723 =  ( n99 ) & ( n7335 )  ;
assign n8724 =  ( n99 ) & ( n7337 )  ;
assign n8725 =  ( n100 ) & ( n7307 )  ;
assign n8726 =  ( n100 ) & ( n7309 )  ;
assign n8727 =  ( n100 ) & ( n7311 )  ;
assign n8728 =  ( n100 ) & ( n7313 )  ;
assign n8729 =  ( n100 ) & ( n7315 )  ;
assign n8730 =  ( n100 ) & ( n7317 )  ;
assign n8731 =  ( n100 ) & ( n7319 )  ;
assign n8732 =  ( n100 ) & ( n7321 )  ;
assign n8733 =  ( n100 ) & ( n7323 )  ;
assign n8734 =  ( n100 ) & ( n7325 )  ;
assign n8735 =  ( n100 ) & ( n7327 )  ;
assign n8736 =  ( n100 ) & ( n7329 )  ;
assign n8737 =  ( n100 ) & ( n7331 )  ;
assign n8738 =  ( n100 ) & ( n7333 )  ;
assign n8739 =  ( n100 ) & ( n7335 )  ;
assign n8740 =  ( n100 ) & ( n7337 )  ;
assign n8741 =  ( n101 ) & ( n7307 )  ;
assign n8742 =  ( n101 ) & ( n7309 )  ;
assign n8743 =  ( n101 ) & ( n7311 )  ;
assign n8744 =  ( n101 ) & ( n7313 )  ;
assign n8745 =  ( n101 ) & ( n7315 )  ;
assign n8746 =  ( n101 ) & ( n7317 )  ;
assign n8747 =  ( n101 ) & ( n7319 )  ;
assign n8748 =  ( n101 ) & ( n7321 )  ;
assign n8749 =  ( n101 ) & ( n7323 )  ;
assign n8750 =  ( n101 ) & ( n7325 )  ;
assign n8751 =  ( n101 ) & ( n7327 )  ;
assign n8752 =  ( n101 ) & ( n7329 )  ;
assign n8753 =  ( n101 ) & ( n7331 )  ;
assign n8754 =  ( n101 ) & ( n7333 )  ;
assign n8755 =  ( n101 ) & ( n7335 )  ;
assign n8756 =  ( n101 ) & ( n7337 )  ;
assign n8757 =  ( n102 ) & ( n7307 )  ;
assign n8758 =  ( n102 ) & ( n7309 )  ;
assign n8759 =  ( n102 ) & ( n7311 )  ;
assign n8760 =  ( n102 ) & ( n7313 )  ;
assign n8761 =  ( n102 ) & ( n7315 )  ;
assign n8762 =  ( n102 ) & ( n7317 )  ;
assign n8763 =  ( n102 ) & ( n7319 )  ;
assign n8764 =  ( n102 ) & ( n7321 )  ;
assign n8765 =  ( n102 ) & ( n7323 )  ;
assign n8766 =  ( n102 ) & ( n7325 )  ;
assign n8767 =  ( n102 ) & ( n7327 )  ;
assign n8768 =  ( n102 ) & ( n7329 )  ;
assign n8769 =  ( n102 ) & ( n7331 )  ;
assign n8770 =  ( n102 ) & ( n7333 )  ;
assign n8771 =  ( n102 ) & ( n7335 )  ;
assign n8772 =  ( n102 ) & ( n7337 )  ;
assign n8773 =  ( n103 ) & ( n7307 )  ;
assign n8774 =  ( n103 ) & ( n7309 )  ;
assign n8775 =  ( n103 ) & ( n7311 )  ;
assign n8776 =  ( n103 ) & ( n7313 )  ;
assign n8777 =  ( n103 ) & ( n7315 )  ;
assign n8778 =  ( n103 ) & ( n7317 )  ;
assign n8779 =  ( n103 ) & ( n7319 )  ;
assign n8780 =  ( n103 ) & ( n7321 )  ;
assign n8781 =  ( n103 ) & ( n7323 )  ;
assign n8782 =  ( n103 ) & ( n7325 )  ;
assign n8783 =  ( n103 ) & ( n7327 )  ;
assign n8784 =  ( n103 ) & ( n7329 )  ;
assign n8785 =  ( n103 ) & ( n7331 )  ;
assign n8786 =  ( n103 ) & ( n7333 )  ;
assign n8787 =  ( n103 ) & ( n7335 )  ;
assign n8788 =  ( n103 ) & ( n7337 )  ;
assign n8789 =  ( n104 ) & ( n7307 )  ;
assign n8790 =  ( n104 ) & ( n7309 )  ;
assign n8791 =  ( n104 ) & ( n7311 )  ;
assign n8792 =  ( n104 ) & ( n7313 )  ;
assign n8793 =  ( n104 ) & ( n7315 )  ;
assign n8794 =  ( n104 ) & ( n7317 )  ;
assign n8795 =  ( n104 ) & ( n7319 )  ;
assign n8796 =  ( n104 ) & ( n7321 )  ;
assign n8797 =  ( n104 ) & ( n7323 )  ;
assign n8798 =  ( n104 ) & ( n7325 )  ;
assign n8799 =  ( n104 ) & ( n7327 )  ;
assign n8800 =  ( n104 ) & ( n7329 )  ;
assign n8801 =  ( n104 ) & ( n7331 )  ;
assign n8802 =  ( n104 ) & ( n7333 )  ;
assign n8803 =  ( n104 ) & ( n7335 )  ;
assign n8804 =  ( n104 ) & ( n7337 )  ;
assign n8805 =  ( n105 ) & ( n7307 )  ;
assign n8806 =  ( n105 ) & ( n7309 )  ;
assign n8807 =  ( n105 ) & ( n7311 )  ;
assign n8808 =  ( n105 ) & ( n7313 )  ;
assign n8809 =  ( n105 ) & ( n7315 )  ;
assign n8810 =  ( n105 ) & ( n7317 )  ;
assign n8811 =  ( n105 ) & ( n7319 )  ;
assign n8812 =  ( n105 ) & ( n7321 )  ;
assign n8813 =  ( n105 ) & ( n7323 )  ;
assign n8814 =  ( n105 ) & ( n7325 )  ;
assign n8815 =  ( n105 ) & ( n7327 )  ;
assign n8816 =  ( n105 ) & ( n7329 )  ;
assign n8817 =  ( n105 ) & ( n7331 )  ;
assign n8818 =  ( n105 ) & ( n7333 )  ;
assign n8819 =  ( n105 ) & ( n7335 )  ;
assign n8820 =  ( n105 ) & ( n7337 )  ;
assign n8821 =  ( n106 ) & ( n7307 )  ;
assign n8822 =  ( n106 ) & ( n7309 )  ;
assign n8823 =  ( n106 ) & ( n7311 )  ;
assign n8824 =  ( n106 ) & ( n7313 )  ;
assign n8825 =  ( n106 ) & ( n7315 )  ;
assign n8826 =  ( n106 ) & ( n7317 )  ;
assign n8827 =  ( n106 ) & ( n7319 )  ;
assign n8828 =  ( n106 ) & ( n7321 )  ;
assign n8829 =  ( n106 ) & ( n7323 )  ;
assign n8830 =  ( n106 ) & ( n7325 )  ;
assign n8831 =  ( n106 ) & ( n7327 )  ;
assign n8832 =  ( n106 ) & ( n7329 )  ;
assign n8833 =  ( n106 ) & ( n7331 )  ;
assign n8834 =  ( n106 ) & ( n7333 )  ;
assign n8835 =  ( n106 ) & ( n7335 )  ;
assign n8836 =  ( n106 ) & ( n7337 )  ;
assign n8837 =  ( n107 ) & ( n7307 )  ;
assign n8838 =  ( n107 ) & ( n7309 )  ;
assign n8839 =  ( n107 ) & ( n7311 )  ;
assign n8840 =  ( n107 ) & ( n7313 )  ;
assign n8841 =  ( n107 ) & ( n7315 )  ;
assign n8842 =  ( n107 ) & ( n7317 )  ;
assign n8843 =  ( n107 ) & ( n7319 )  ;
assign n8844 =  ( n107 ) & ( n7321 )  ;
assign n8845 =  ( n107 ) & ( n7323 )  ;
assign n8846 =  ( n107 ) & ( n7325 )  ;
assign n8847 =  ( n107 ) & ( n7327 )  ;
assign n8848 =  ( n107 ) & ( n7329 )  ;
assign n8849 =  ( n107 ) & ( n7331 )  ;
assign n8850 =  ( n107 ) & ( n7333 )  ;
assign n8851 =  ( n107 ) & ( n7335 )  ;
assign n8852 =  ( n107 ) & ( n7337 )  ;
assign n8853 =  ( n108 ) & ( n7307 )  ;
assign n8854 =  ( n108 ) & ( n7309 )  ;
assign n8855 =  ( n108 ) & ( n7311 )  ;
assign n8856 =  ( n108 ) & ( n7313 )  ;
assign n8857 =  ( n108 ) & ( n7315 )  ;
assign n8858 =  ( n108 ) & ( n7317 )  ;
assign n8859 =  ( n108 ) & ( n7319 )  ;
assign n8860 =  ( n108 ) & ( n7321 )  ;
assign n8861 =  ( n108 ) & ( n7323 )  ;
assign n8862 =  ( n108 ) & ( n7325 )  ;
assign n8863 =  ( n108 ) & ( n7327 )  ;
assign n8864 =  ( n108 ) & ( n7329 )  ;
assign n8865 =  ( n108 ) & ( n7331 )  ;
assign n8866 =  ( n108 ) & ( n7333 )  ;
assign n8867 =  ( n108 ) & ( n7335 )  ;
assign n8868 =  ( n108 ) & ( n7337 )  ;
assign n8869 =  ( n8868 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n8870 =  ( n8867 ) ? ( VREG_0_1 ) : ( n8869 ) ;
assign n8871 =  ( n8866 ) ? ( VREG_0_2 ) : ( n8870 ) ;
assign n8872 =  ( n8865 ) ? ( VREG_0_3 ) : ( n8871 ) ;
assign n8873 =  ( n8864 ) ? ( VREG_0_4 ) : ( n8872 ) ;
assign n8874 =  ( n8863 ) ? ( VREG_0_5 ) : ( n8873 ) ;
assign n8875 =  ( n8862 ) ? ( VREG_0_6 ) : ( n8874 ) ;
assign n8876 =  ( n8861 ) ? ( VREG_0_7 ) : ( n8875 ) ;
assign n8877 =  ( n8860 ) ? ( VREG_0_8 ) : ( n8876 ) ;
assign n8878 =  ( n8859 ) ? ( VREG_0_9 ) : ( n8877 ) ;
assign n8879 =  ( n8858 ) ? ( VREG_0_10 ) : ( n8878 ) ;
assign n8880 =  ( n8857 ) ? ( VREG_0_11 ) : ( n8879 ) ;
assign n8881 =  ( n8856 ) ? ( VREG_0_12 ) : ( n8880 ) ;
assign n8882 =  ( n8855 ) ? ( VREG_0_13 ) : ( n8881 ) ;
assign n8883 =  ( n8854 ) ? ( VREG_0_14 ) : ( n8882 ) ;
assign n8884 =  ( n8853 ) ? ( VREG_0_15 ) : ( n8883 ) ;
assign n8885 =  ( n8852 ) ? ( VREG_1_0 ) : ( n8884 ) ;
assign n8886 =  ( n8851 ) ? ( VREG_1_1 ) : ( n8885 ) ;
assign n8887 =  ( n8850 ) ? ( VREG_1_2 ) : ( n8886 ) ;
assign n8888 =  ( n8849 ) ? ( VREG_1_3 ) : ( n8887 ) ;
assign n8889 =  ( n8848 ) ? ( VREG_1_4 ) : ( n8888 ) ;
assign n8890 =  ( n8847 ) ? ( VREG_1_5 ) : ( n8889 ) ;
assign n8891 =  ( n8846 ) ? ( VREG_1_6 ) : ( n8890 ) ;
assign n8892 =  ( n8845 ) ? ( VREG_1_7 ) : ( n8891 ) ;
assign n8893 =  ( n8844 ) ? ( VREG_1_8 ) : ( n8892 ) ;
assign n8894 =  ( n8843 ) ? ( VREG_1_9 ) : ( n8893 ) ;
assign n8895 =  ( n8842 ) ? ( VREG_1_10 ) : ( n8894 ) ;
assign n8896 =  ( n8841 ) ? ( VREG_1_11 ) : ( n8895 ) ;
assign n8897 =  ( n8840 ) ? ( VREG_1_12 ) : ( n8896 ) ;
assign n8898 =  ( n8839 ) ? ( VREG_1_13 ) : ( n8897 ) ;
assign n8899 =  ( n8838 ) ? ( VREG_1_14 ) : ( n8898 ) ;
assign n8900 =  ( n8837 ) ? ( VREG_1_15 ) : ( n8899 ) ;
assign n8901 =  ( n8836 ) ? ( VREG_2_0 ) : ( n8900 ) ;
assign n8902 =  ( n8835 ) ? ( VREG_2_1 ) : ( n8901 ) ;
assign n8903 =  ( n8834 ) ? ( VREG_2_2 ) : ( n8902 ) ;
assign n8904 =  ( n8833 ) ? ( VREG_2_3 ) : ( n8903 ) ;
assign n8905 =  ( n8832 ) ? ( VREG_2_4 ) : ( n8904 ) ;
assign n8906 =  ( n8831 ) ? ( VREG_2_5 ) : ( n8905 ) ;
assign n8907 =  ( n8830 ) ? ( VREG_2_6 ) : ( n8906 ) ;
assign n8908 =  ( n8829 ) ? ( VREG_2_7 ) : ( n8907 ) ;
assign n8909 =  ( n8828 ) ? ( VREG_2_8 ) : ( n8908 ) ;
assign n8910 =  ( n8827 ) ? ( VREG_2_9 ) : ( n8909 ) ;
assign n8911 =  ( n8826 ) ? ( VREG_2_10 ) : ( n8910 ) ;
assign n8912 =  ( n8825 ) ? ( VREG_2_11 ) : ( n8911 ) ;
assign n8913 =  ( n8824 ) ? ( VREG_2_12 ) : ( n8912 ) ;
assign n8914 =  ( n8823 ) ? ( VREG_2_13 ) : ( n8913 ) ;
assign n8915 =  ( n8822 ) ? ( VREG_2_14 ) : ( n8914 ) ;
assign n8916 =  ( n8821 ) ? ( VREG_2_15 ) : ( n8915 ) ;
assign n8917 =  ( n8820 ) ? ( VREG_3_0 ) : ( n8916 ) ;
assign n8918 =  ( n8819 ) ? ( VREG_3_1 ) : ( n8917 ) ;
assign n8919 =  ( n8818 ) ? ( VREG_3_2 ) : ( n8918 ) ;
assign n8920 =  ( n8817 ) ? ( VREG_3_3 ) : ( n8919 ) ;
assign n8921 =  ( n8816 ) ? ( VREG_3_4 ) : ( n8920 ) ;
assign n8922 =  ( n8815 ) ? ( VREG_3_5 ) : ( n8921 ) ;
assign n8923 =  ( n8814 ) ? ( VREG_3_6 ) : ( n8922 ) ;
assign n8924 =  ( n8813 ) ? ( VREG_3_7 ) : ( n8923 ) ;
assign n8925 =  ( n8812 ) ? ( VREG_3_8 ) : ( n8924 ) ;
assign n8926 =  ( n8811 ) ? ( VREG_3_9 ) : ( n8925 ) ;
assign n8927 =  ( n8810 ) ? ( VREG_3_10 ) : ( n8926 ) ;
assign n8928 =  ( n8809 ) ? ( VREG_3_11 ) : ( n8927 ) ;
assign n8929 =  ( n8808 ) ? ( VREG_3_12 ) : ( n8928 ) ;
assign n8930 =  ( n8807 ) ? ( VREG_3_13 ) : ( n8929 ) ;
assign n8931 =  ( n8806 ) ? ( VREG_3_14 ) : ( n8930 ) ;
assign n8932 =  ( n8805 ) ? ( VREG_3_15 ) : ( n8931 ) ;
assign n8933 =  ( n8804 ) ? ( VREG_4_0 ) : ( n8932 ) ;
assign n8934 =  ( n8803 ) ? ( VREG_4_1 ) : ( n8933 ) ;
assign n8935 =  ( n8802 ) ? ( VREG_4_2 ) : ( n8934 ) ;
assign n8936 =  ( n8801 ) ? ( VREG_4_3 ) : ( n8935 ) ;
assign n8937 =  ( n8800 ) ? ( VREG_4_4 ) : ( n8936 ) ;
assign n8938 =  ( n8799 ) ? ( VREG_4_5 ) : ( n8937 ) ;
assign n8939 =  ( n8798 ) ? ( VREG_4_6 ) : ( n8938 ) ;
assign n8940 =  ( n8797 ) ? ( VREG_4_7 ) : ( n8939 ) ;
assign n8941 =  ( n8796 ) ? ( VREG_4_8 ) : ( n8940 ) ;
assign n8942 =  ( n8795 ) ? ( VREG_4_9 ) : ( n8941 ) ;
assign n8943 =  ( n8794 ) ? ( VREG_4_10 ) : ( n8942 ) ;
assign n8944 =  ( n8793 ) ? ( VREG_4_11 ) : ( n8943 ) ;
assign n8945 =  ( n8792 ) ? ( VREG_4_12 ) : ( n8944 ) ;
assign n8946 =  ( n8791 ) ? ( VREG_4_13 ) : ( n8945 ) ;
assign n8947 =  ( n8790 ) ? ( VREG_4_14 ) : ( n8946 ) ;
assign n8948 =  ( n8789 ) ? ( VREG_4_15 ) : ( n8947 ) ;
assign n8949 =  ( n8788 ) ? ( VREG_5_0 ) : ( n8948 ) ;
assign n8950 =  ( n8787 ) ? ( VREG_5_1 ) : ( n8949 ) ;
assign n8951 =  ( n8786 ) ? ( VREG_5_2 ) : ( n8950 ) ;
assign n8952 =  ( n8785 ) ? ( VREG_5_3 ) : ( n8951 ) ;
assign n8953 =  ( n8784 ) ? ( VREG_5_4 ) : ( n8952 ) ;
assign n8954 =  ( n8783 ) ? ( VREG_5_5 ) : ( n8953 ) ;
assign n8955 =  ( n8782 ) ? ( VREG_5_6 ) : ( n8954 ) ;
assign n8956 =  ( n8781 ) ? ( VREG_5_7 ) : ( n8955 ) ;
assign n8957 =  ( n8780 ) ? ( VREG_5_8 ) : ( n8956 ) ;
assign n8958 =  ( n8779 ) ? ( VREG_5_9 ) : ( n8957 ) ;
assign n8959 =  ( n8778 ) ? ( VREG_5_10 ) : ( n8958 ) ;
assign n8960 =  ( n8777 ) ? ( VREG_5_11 ) : ( n8959 ) ;
assign n8961 =  ( n8776 ) ? ( VREG_5_12 ) : ( n8960 ) ;
assign n8962 =  ( n8775 ) ? ( VREG_5_13 ) : ( n8961 ) ;
assign n8963 =  ( n8774 ) ? ( VREG_5_14 ) : ( n8962 ) ;
assign n8964 =  ( n8773 ) ? ( VREG_5_15 ) : ( n8963 ) ;
assign n8965 =  ( n8772 ) ? ( VREG_6_0 ) : ( n8964 ) ;
assign n8966 =  ( n8771 ) ? ( VREG_6_1 ) : ( n8965 ) ;
assign n8967 =  ( n8770 ) ? ( VREG_6_2 ) : ( n8966 ) ;
assign n8968 =  ( n8769 ) ? ( VREG_6_3 ) : ( n8967 ) ;
assign n8969 =  ( n8768 ) ? ( VREG_6_4 ) : ( n8968 ) ;
assign n8970 =  ( n8767 ) ? ( VREG_6_5 ) : ( n8969 ) ;
assign n8971 =  ( n8766 ) ? ( VREG_6_6 ) : ( n8970 ) ;
assign n8972 =  ( n8765 ) ? ( VREG_6_7 ) : ( n8971 ) ;
assign n8973 =  ( n8764 ) ? ( VREG_6_8 ) : ( n8972 ) ;
assign n8974 =  ( n8763 ) ? ( VREG_6_9 ) : ( n8973 ) ;
assign n8975 =  ( n8762 ) ? ( VREG_6_10 ) : ( n8974 ) ;
assign n8976 =  ( n8761 ) ? ( VREG_6_11 ) : ( n8975 ) ;
assign n8977 =  ( n8760 ) ? ( VREG_6_12 ) : ( n8976 ) ;
assign n8978 =  ( n8759 ) ? ( VREG_6_13 ) : ( n8977 ) ;
assign n8979 =  ( n8758 ) ? ( VREG_6_14 ) : ( n8978 ) ;
assign n8980 =  ( n8757 ) ? ( VREG_6_15 ) : ( n8979 ) ;
assign n8981 =  ( n8756 ) ? ( VREG_7_0 ) : ( n8980 ) ;
assign n8982 =  ( n8755 ) ? ( VREG_7_1 ) : ( n8981 ) ;
assign n8983 =  ( n8754 ) ? ( VREG_7_2 ) : ( n8982 ) ;
assign n8984 =  ( n8753 ) ? ( VREG_7_3 ) : ( n8983 ) ;
assign n8985 =  ( n8752 ) ? ( VREG_7_4 ) : ( n8984 ) ;
assign n8986 =  ( n8751 ) ? ( VREG_7_5 ) : ( n8985 ) ;
assign n8987 =  ( n8750 ) ? ( VREG_7_6 ) : ( n8986 ) ;
assign n8988 =  ( n8749 ) ? ( VREG_7_7 ) : ( n8987 ) ;
assign n8989 =  ( n8748 ) ? ( VREG_7_8 ) : ( n8988 ) ;
assign n8990 =  ( n8747 ) ? ( VREG_7_9 ) : ( n8989 ) ;
assign n8991 =  ( n8746 ) ? ( VREG_7_10 ) : ( n8990 ) ;
assign n8992 =  ( n8745 ) ? ( VREG_7_11 ) : ( n8991 ) ;
assign n8993 =  ( n8744 ) ? ( VREG_7_12 ) : ( n8992 ) ;
assign n8994 =  ( n8743 ) ? ( VREG_7_13 ) : ( n8993 ) ;
assign n8995 =  ( n8742 ) ? ( VREG_7_14 ) : ( n8994 ) ;
assign n8996 =  ( n8741 ) ? ( VREG_7_15 ) : ( n8995 ) ;
assign n8997 =  ( n8740 ) ? ( VREG_8_0 ) : ( n8996 ) ;
assign n8998 =  ( n8739 ) ? ( VREG_8_1 ) : ( n8997 ) ;
assign n8999 =  ( n8738 ) ? ( VREG_8_2 ) : ( n8998 ) ;
assign n9000 =  ( n8737 ) ? ( VREG_8_3 ) : ( n8999 ) ;
assign n9001 =  ( n8736 ) ? ( VREG_8_4 ) : ( n9000 ) ;
assign n9002 =  ( n8735 ) ? ( VREG_8_5 ) : ( n9001 ) ;
assign n9003 =  ( n8734 ) ? ( VREG_8_6 ) : ( n9002 ) ;
assign n9004 =  ( n8733 ) ? ( VREG_8_7 ) : ( n9003 ) ;
assign n9005 =  ( n8732 ) ? ( VREG_8_8 ) : ( n9004 ) ;
assign n9006 =  ( n8731 ) ? ( VREG_8_9 ) : ( n9005 ) ;
assign n9007 =  ( n8730 ) ? ( VREG_8_10 ) : ( n9006 ) ;
assign n9008 =  ( n8729 ) ? ( VREG_8_11 ) : ( n9007 ) ;
assign n9009 =  ( n8728 ) ? ( VREG_8_12 ) : ( n9008 ) ;
assign n9010 =  ( n8727 ) ? ( VREG_8_13 ) : ( n9009 ) ;
assign n9011 =  ( n8726 ) ? ( VREG_8_14 ) : ( n9010 ) ;
assign n9012 =  ( n8725 ) ? ( VREG_8_15 ) : ( n9011 ) ;
assign n9013 =  ( n8724 ) ? ( VREG_9_0 ) : ( n9012 ) ;
assign n9014 =  ( n8723 ) ? ( VREG_9_1 ) : ( n9013 ) ;
assign n9015 =  ( n8722 ) ? ( VREG_9_2 ) : ( n9014 ) ;
assign n9016 =  ( n8721 ) ? ( VREG_9_3 ) : ( n9015 ) ;
assign n9017 =  ( n8720 ) ? ( VREG_9_4 ) : ( n9016 ) ;
assign n9018 =  ( n8719 ) ? ( VREG_9_5 ) : ( n9017 ) ;
assign n9019 =  ( n8718 ) ? ( VREG_9_6 ) : ( n9018 ) ;
assign n9020 =  ( n8717 ) ? ( VREG_9_7 ) : ( n9019 ) ;
assign n9021 =  ( n8716 ) ? ( VREG_9_8 ) : ( n9020 ) ;
assign n9022 =  ( n8715 ) ? ( VREG_9_9 ) : ( n9021 ) ;
assign n9023 =  ( n8714 ) ? ( VREG_9_10 ) : ( n9022 ) ;
assign n9024 =  ( n8713 ) ? ( VREG_9_11 ) : ( n9023 ) ;
assign n9025 =  ( n8712 ) ? ( VREG_9_12 ) : ( n9024 ) ;
assign n9026 =  ( n8711 ) ? ( VREG_9_13 ) : ( n9025 ) ;
assign n9027 =  ( n8710 ) ? ( VREG_9_14 ) : ( n9026 ) ;
assign n9028 =  ( n8709 ) ? ( VREG_9_15 ) : ( n9027 ) ;
assign n9029 =  ( n8708 ) ? ( VREG_10_0 ) : ( n9028 ) ;
assign n9030 =  ( n8707 ) ? ( VREG_10_1 ) : ( n9029 ) ;
assign n9031 =  ( n8706 ) ? ( VREG_10_2 ) : ( n9030 ) ;
assign n9032 =  ( n8705 ) ? ( VREG_10_3 ) : ( n9031 ) ;
assign n9033 =  ( n8704 ) ? ( VREG_10_4 ) : ( n9032 ) ;
assign n9034 =  ( n8703 ) ? ( VREG_10_5 ) : ( n9033 ) ;
assign n9035 =  ( n8702 ) ? ( VREG_10_6 ) : ( n9034 ) ;
assign n9036 =  ( n8701 ) ? ( VREG_10_7 ) : ( n9035 ) ;
assign n9037 =  ( n8700 ) ? ( VREG_10_8 ) : ( n9036 ) ;
assign n9038 =  ( n8699 ) ? ( VREG_10_9 ) : ( n9037 ) ;
assign n9039 =  ( n8698 ) ? ( VREG_10_10 ) : ( n9038 ) ;
assign n9040 =  ( n8697 ) ? ( VREG_10_11 ) : ( n9039 ) ;
assign n9041 =  ( n8696 ) ? ( VREG_10_12 ) : ( n9040 ) ;
assign n9042 =  ( n8695 ) ? ( VREG_10_13 ) : ( n9041 ) ;
assign n9043 =  ( n8694 ) ? ( VREG_10_14 ) : ( n9042 ) ;
assign n9044 =  ( n8693 ) ? ( VREG_10_15 ) : ( n9043 ) ;
assign n9045 =  ( n8692 ) ? ( VREG_11_0 ) : ( n9044 ) ;
assign n9046 =  ( n8691 ) ? ( VREG_11_1 ) : ( n9045 ) ;
assign n9047 =  ( n8690 ) ? ( VREG_11_2 ) : ( n9046 ) ;
assign n9048 =  ( n8689 ) ? ( VREG_11_3 ) : ( n9047 ) ;
assign n9049 =  ( n8688 ) ? ( VREG_11_4 ) : ( n9048 ) ;
assign n9050 =  ( n8687 ) ? ( VREG_11_5 ) : ( n9049 ) ;
assign n9051 =  ( n8686 ) ? ( VREG_11_6 ) : ( n9050 ) ;
assign n9052 =  ( n8685 ) ? ( VREG_11_7 ) : ( n9051 ) ;
assign n9053 =  ( n8684 ) ? ( VREG_11_8 ) : ( n9052 ) ;
assign n9054 =  ( n8683 ) ? ( VREG_11_9 ) : ( n9053 ) ;
assign n9055 =  ( n8682 ) ? ( VREG_11_10 ) : ( n9054 ) ;
assign n9056 =  ( n8681 ) ? ( VREG_11_11 ) : ( n9055 ) ;
assign n9057 =  ( n8680 ) ? ( VREG_11_12 ) : ( n9056 ) ;
assign n9058 =  ( n8679 ) ? ( VREG_11_13 ) : ( n9057 ) ;
assign n9059 =  ( n8678 ) ? ( VREG_11_14 ) : ( n9058 ) ;
assign n9060 =  ( n8677 ) ? ( VREG_11_15 ) : ( n9059 ) ;
assign n9061 =  ( n8676 ) ? ( VREG_12_0 ) : ( n9060 ) ;
assign n9062 =  ( n8675 ) ? ( VREG_12_1 ) : ( n9061 ) ;
assign n9063 =  ( n8674 ) ? ( VREG_12_2 ) : ( n9062 ) ;
assign n9064 =  ( n8673 ) ? ( VREG_12_3 ) : ( n9063 ) ;
assign n9065 =  ( n8672 ) ? ( VREG_12_4 ) : ( n9064 ) ;
assign n9066 =  ( n8671 ) ? ( VREG_12_5 ) : ( n9065 ) ;
assign n9067 =  ( n8670 ) ? ( VREG_12_6 ) : ( n9066 ) ;
assign n9068 =  ( n8669 ) ? ( VREG_12_7 ) : ( n9067 ) ;
assign n9069 =  ( n8668 ) ? ( VREG_12_8 ) : ( n9068 ) ;
assign n9070 =  ( n8667 ) ? ( VREG_12_9 ) : ( n9069 ) ;
assign n9071 =  ( n8666 ) ? ( VREG_12_10 ) : ( n9070 ) ;
assign n9072 =  ( n8665 ) ? ( VREG_12_11 ) : ( n9071 ) ;
assign n9073 =  ( n8664 ) ? ( VREG_12_12 ) : ( n9072 ) ;
assign n9074 =  ( n8663 ) ? ( VREG_12_13 ) : ( n9073 ) ;
assign n9075 =  ( n8662 ) ? ( VREG_12_14 ) : ( n9074 ) ;
assign n9076 =  ( n8661 ) ? ( VREG_12_15 ) : ( n9075 ) ;
assign n9077 =  ( n8660 ) ? ( VREG_13_0 ) : ( n9076 ) ;
assign n9078 =  ( n8659 ) ? ( VREG_13_1 ) : ( n9077 ) ;
assign n9079 =  ( n8658 ) ? ( VREG_13_2 ) : ( n9078 ) ;
assign n9080 =  ( n8657 ) ? ( VREG_13_3 ) : ( n9079 ) ;
assign n9081 =  ( n8656 ) ? ( VREG_13_4 ) : ( n9080 ) ;
assign n9082 =  ( n8655 ) ? ( VREG_13_5 ) : ( n9081 ) ;
assign n9083 =  ( n8654 ) ? ( VREG_13_6 ) : ( n9082 ) ;
assign n9084 =  ( n8653 ) ? ( VREG_13_7 ) : ( n9083 ) ;
assign n9085 =  ( n8652 ) ? ( VREG_13_8 ) : ( n9084 ) ;
assign n9086 =  ( n8651 ) ? ( VREG_13_9 ) : ( n9085 ) ;
assign n9087 =  ( n8650 ) ? ( VREG_13_10 ) : ( n9086 ) ;
assign n9088 =  ( n8649 ) ? ( VREG_13_11 ) : ( n9087 ) ;
assign n9089 =  ( n8648 ) ? ( VREG_13_12 ) : ( n9088 ) ;
assign n9090 =  ( n8647 ) ? ( VREG_13_13 ) : ( n9089 ) ;
assign n9091 =  ( n8646 ) ? ( VREG_13_14 ) : ( n9090 ) ;
assign n9092 =  ( n8645 ) ? ( VREG_13_15 ) : ( n9091 ) ;
assign n9093 =  ( n8644 ) ? ( VREG_14_0 ) : ( n9092 ) ;
assign n9094 =  ( n8643 ) ? ( VREG_14_1 ) : ( n9093 ) ;
assign n9095 =  ( n8642 ) ? ( VREG_14_2 ) : ( n9094 ) ;
assign n9096 =  ( n8641 ) ? ( VREG_14_3 ) : ( n9095 ) ;
assign n9097 =  ( n8640 ) ? ( VREG_14_4 ) : ( n9096 ) ;
assign n9098 =  ( n8639 ) ? ( VREG_14_5 ) : ( n9097 ) ;
assign n9099 =  ( n8638 ) ? ( VREG_14_6 ) : ( n9098 ) ;
assign n9100 =  ( n8637 ) ? ( VREG_14_7 ) : ( n9099 ) ;
assign n9101 =  ( n8636 ) ? ( VREG_14_8 ) : ( n9100 ) ;
assign n9102 =  ( n8635 ) ? ( VREG_14_9 ) : ( n9101 ) ;
assign n9103 =  ( n8634 ) ? ( VREG_14_10 ) : ( n9102 ) ;
assign n9104 =  ( n8633 ) ? ( VREG_14_11 ) : ( n9103 ) ;
assign n9105 =  ( n8632 ) ? ( VREG_14_12 ) : ( n9104 ) ;
assign n9106 =  ( n8631 ) ? ( VREG_14_13 ) : ( n9105 ) ;
assign n9107 =  ( n8630 ) ? ( VREG_14_14 ) : ( n9106 ) ;
assign n9108 =  ( n8629 ) ? ( VREG_14_15 ) : ( n9107 ) ;
assign n9109 =  ( n8628 ) ? ( VREG_15_0 ) : ( n9108 ) ;
assign n9110 =  ( n8627 ) ? ( VREG_15_1 ) : ( n9109 ) ;
assign n9111 =  ( n8626 ) ? ( VREG_15_2 ) : ( n9110 ) ;
assign n9112 =  ( n8625 ) ? ( VREG_15_3 ) : ( n9111 ) ;
assign n9113 =  ( n8624 ) ? ( VREG_15_4 ) : ( n9112 ) ;
assign n9114 =  ( n8623 ) ? ( VREG_15_5 ) : ( n9113 ) ;
assign n9115 =  ( n8622 ) ? ( VREG_15_6 ) : ( n9114 ) ;
assign n9116 =  ( n8621 ) ? ( VREG_15_7 ) : ( n9115 ) ;
assign n9117 =  ( n8620 ) ? ( VREG_15_8 ) : ( n9116 ) ;
assign n9118 =  ( n8619 ) ? ( VREG_15_9 ) : ( n9117 ) ;
assign n9119 =  ( n8618 ) ? ( VREG_15_10 ) : ( n9118 ) ;
assign n9120 =  ( n8617 ) ? ( VREG_15_11 ) : ( n9119 ) ;
assign n9121 =  ( n8616 ) ? ( VREG_15_12 ) : ( n9120 ) ;
assign n9122 =  ( n8615 ) ? ( VREG_15_13 ) : ( n9121 ) ;
assign n9123 =  ( n8614 ) ? ( VREG_15_14 ) : ( n9122 ) ;
assign n9124 =  ( n8613 ) ? ( VREG_15_15 ) : ( n9123 ) ;
assign n9125 =  ( n8612 ) ? ( VREG_16_0 ) : ( n9124 ) ;
assign n9126 =  ( n8611 ) ? ( VREG_16_1 ) : ( n9125 ) ;
assign n9127 =  ( n8610 ) ? ( VREG_16_2 ) : ( n9126 ) ;
assign n9128 =  ( n8609 ) ? ( VREG_16_3 ) : ( n9127 ) ;
assign n9129 =  ( n8608 ) ? ( VREG_16_4 ) : ( n9128 ) ;
assign n9130 =  ( n8607 ) ? ( VREG_16_5 ) : ( n9129 ) ;
assign n9131 =  ( n8606 ) ? ( VREG_16_6 ) : ( n9130 ) ;
assign n9132 =  ( n8605 ) ? ( VREG_16_7 ) : ( n9131 ) ;
assign n9133 =  ( n8604 ) ? ( VREG_16_8 ) : ( n9132 ) ;
assign n9134 =  ( n8603 ) ? ( VREG_16_9 ) : ( n9133 ) ;
assign n9135 =  ( n8602 ) ? ( VREG_16_10 ) : ( n9134 ) ;
assign n9136 =  ( n8601 ) ? ( VREG_16_11 ) : ( n9135 ) ;
assign n9137 =  ( n8600 ) ? ( VREG_16_12 ) : ( n9136 ) ;
assign n9138 =  ( n8599 ) ? ( VREG_16_13 ) : ( n9137 ) ;
assign n9139 =  ( n8598 ) ? ( VREG_16_14 ) : ( n9138 ) ;
assign n9140 =  ( n8597 ) ? ( VREG_16_15 ) : ( n9139 ) ;
assign n9141 =  ( n8596 ) ? ( VREG_17_0 ) : ( n9140 ) ;
assign n9142 =  ( n8595 ) ? ( VREG_17_1 ) : ( n9141 ) ;
assign n9143 =  ( n8594 ) ? ( VREG_17_2 ) : ( n9142 ) ;
assign n9144 =  ( n8593 ) ? ( VREG_17_3 ) : ( n9143 ) ;
assign n9145 =  ( n8592 ) ? ( VREG_17_4 ) : ( n9144 ) ;
assign n9146 =  ( n8591 ) ? ( VREG_17_5 ) : ( n9145 ) ;
assign n9147 =  ( n8590 ) ? ( VREG_17_6 ) : ( n9146 ) ;
assign n9148 =  ( n8589 ) ? ( VREG_17_7 ) : ( n9147 ) ;
assign n9149 =  ( n8588 ) ? ( VREG_17_8 ) : ( n9148 ) ;
assign n9150 =  ( n8587 ) ? ( VREG_17_9 ) : ( n9149 ) ;
assign n9151 =  ( n8586 ) ? ( VREG_17_10 ) : ( n9150 ) ;
assign n9152 =  ( n8585 ) ? ( VREG_17_11 ) : ( n9151 ) ;
assign n9153 =  ( n8584 ) ? ( VREG_17_12 ) : ( n9152 ) ;
assign n9154 =  ( n8583 ) ? ( VREG_17_13 ) : ( n9153 ) ;
assign n9155 =  ( n8582 ) ? ( VREG_17_14 ) : ( n9154 ) ;
assign n9156 =  ( n8581 ) ? ( VREG_17_15 ) : ( n9155 ) ;
assign n9157 =  ( n8580 ) ? ( VREG_18_0 ) : ( n9156 ) ;
assign n9158 =  ( n8579 ) ? ( VREG_18_1 ) : ( n9157 ) ;
assign n9159 =  ( n8578 ) ? ( VREG_18_2 ) : ( n9158 ) ;
assign n9160 =  ( n8577 ) ? ( VREG_18_3 ) : ( n9159 ) ;
assign n9161 =  ( n8576 ) ? ( VREG_18_4 ) : ( n9160 ) ;
assign n9162 =  ( n8575 ) ? ( VREG_18_5 ) : ( n9161 ) ;
assign n9163 =  ( n8574 ) ? ( VREG_18_6 ) : ( n9162 ) ;
assign n9164 =  ( n8573 ) ? ( VREG_18_7 ) : ( n9163 ) ;
assign n9165 =  ( n8572 ) ? ( VREG_18_8 ) : ( n9164 ) ;
assign n9166 =  ( n8571 ) ? ( VREG_18_9 ) : ( n9165 ) ;
assign n9167 =  ( n8570 ) ? ( VREG_18_10 ) : ( n9166 ) ;
assign n9168 =  ( n8569 ) ? ( VREG_18_11 ) : ( n9167 ) ;
assign n9169 =  ( n8568 ) ? ( VREG_18_12 ) : ( n9168 ) ;
assign n9170 =  ( n8567 ) ? ( VREG_18_13 ) : ( n9169 ) ;
assign n9171 =  ( n8566 ) ? ( VREG_18_14 ) : ( n9170 ) ;
assign n9172 =  ( n8565 ) ? ( VREG_18_15 ) : ( n9171 ) ;
assign n9173 =  ( n8564 ) ? ( VREG_19_0 ) : ( n9172 ) ;
assign n9174 =  ( n8563 ) ? ( VREG_19_1 ) : ( n9173 ) ;
assign n9175 =  ( n8562 ) ? ( VREG_19_2 ) : ( n9174 ) ;
assign n9176 =  ( n8561 ) ? ( VREG_19_3 ) : ( n9175 ) ;
assign n9177 =  ( n8560 ) ? ( VREG_19_4 ) : ( n9176 ) ;
assign n9178 =  ( n8559 ) ? ( VREG_19_5 ) : ( n9177 ) ;
assign n9179 =  ( n8558 ) ? ( VREG_19_6 ) : ( n9178 ) ;
assign n9180 =  ( n8557 ) ? ( VREG_19_7 ) : ( n9179 ) ;
assign n9181 =  ( n8556 ) ? ( VREG_19_8 ) : ( n9180 ) ;
assign n9182 =  ( n8555 ) ? ( VREG_19_9 ) : ( n9181 ) ;
assign n9183 =  ( n8554 ) ? ( VREG_19_10 ) : ( n9182 ) ;
assign n9184 =  ( n8553 ) ? ( VREG_19_11 ) : ( n9183 ) ;
assign n9185 =  ( n8552 ) ? ( VREG_19_12 ) : ( n9184 ) ;
assign n9186 =  ( n8551 ) ? ( VREG_19_13 ) : ( n9185 ) ;
assign n9187 =  ( n8550 ) ? ( VREG_19_14 ) : ( n9186 ) ;
assign n9188 =  ( n8549 ) ? ( VREG_19_15 ) : ( n9187 ) ;
assign n9189 =  ( n8548 ) ? ( VREG_20_0 ) : ( n9188 ) ;
assign n9190 =  ( n8547 ) ? ( VREG_20_1 ) : ( n9189 ) ;
assign n9191 =  ( n8546 ) ? ( VREG_20_2 ) : ( n9190 ) ;
assign n9192 =  ( n8545 ) ? ( VREG_20_3 ) : ( n9191 ) ;
assign n9193 =  ( n8544 ) ? ( VREG_20_4 ) : ( n9192 ) ;
assign n9194 =  ( n8543 ) ? ( VREG_20_5 ) : ( n9193 ) ;
assign n9195 =  ( n8542 ) ? ( VREG_20_6 ) : ( n9194 ) ;
assign n9196 =  ( n8541 ) ? ( VREG_20_7 ) : ( n9195 ) ;
assign n9197 =  ( n8540 ) ? ( VREG_20_8 ) : ( n9196 ) ;
assign n9198 =  ( n8539 ) ? ( VREG_20_9 ) : ( n9197 ) ;
assign n9199 =  ( n8538 ) ? ( VREG_20_10 ) : ( n9198 ) ;
assign n9200 =  ( n8537 ) ? ( VREG_20_11 ) : ( n9199 ) ;
assign n9201 =  ( n8536 ) ? ( VREG_20_12 ) : ( n9200 ) ;
assign n9202 =  ( n8535 ) ? ( VREG_20_13 ) : ( n9201 ) ;
assign n9203 =  ( n8534 ) ? ( VREG_20_14 ) : ( n9202 ) ;
assign n9204 =  ( n8533 ) ? ( VREG_20_15 ) : ( n9203 ) ;
assign n9205 =  ( n8532 ) ? ( VREG_21_0 ) : ( n9204 ) ;
assign n9206 =  ( n8531 ) ? ( VREG_21_1 ) : ( n9205 ) ;
assign n9207 =  ( n8530 ) ? ( VREG_21_2 ) : ( n9206 ) ;
assign n9208 =  ( n8529 ) ? ( VREG_21_3 ) : ( n9207 ) ;
assign n9209 =  ( n8528 ) ? ( VREG_21_4 ) : ( n9208 ) ;
assign n9210 =  ( n8527 ) ? ( VREG_21_5 ) : ( n9209 ) ;
assign n9211 =  ( n8526 ) ? ( VREG_21_6 ) : ( n9210 ) ;
assign n9212 =  ( n8525 ) ? ( VREG_21_7 ) : ( n9211 ) ;
assign n9213 =  ( n8524 ) ? ( VREG_21_8 ) : ( n9212 ) ;
assign n9214 =  ( n8523 ) ? ( VREG_21_9 ) : ( n9213 ) ;
assign n9215 =  ( n8522 ) ? ( VREG_21_10 ) : ( n9214 ) ;
assign n9216 =  ( n8521 ) ? ( VREG_21_11 ) : ( n9215 ) ;
assign n9217 =  ( n8520 ) ? ( VREG_21_12 ) : ( n9216 ) ;
assign n9218 =  ( n8519 ) ? ( VREG_21_13 ) : ( n9217 ) ;
assign n9219 =  ( n8518 ) ? ( VREG_21_14 ) : ( n9218 ) ;
assign n9220 =  ( n8517 ) ? ( VREG_21_15 ) : ( n9219 ) ;
assign n9221 =  ( n8516 ) ? ( VREG_22_0 ) : ( n9220 ) ;
assign n9222 =  ( n8515 ) ? ( VREG_22_1 ) : ( n9221 ) ;
assign n9223 =  ( n8514 ) ? ( VREG_22_2 ) : ( n9222 ) ;
assign n9224 =  ( n8513 ) ? ( VREG_22_3 ) : ( n9223 ) ;
assign n9225 =  ( n8512 ) ? ( VREG_22_4 ) : ( n9224 ) ;
assign n9226 =  ( n8511 ) ? ( VREG_22_5 ) : ( n9225 ) ;
assign n9227 =  ( n8510 ) ? ( VREG_22_6 ) : ( n9226 ) ;
assign n9228 =  ( n8509 ) ? ( VREG_22_7 ) : ( n9227 ) ;
assign n9229 =  ( n8508 ) ? ( VREG_22_8 ) : ( n9228 ) ;
assign n9230 =  ( n8507 ) ? ( VREG_22_9 ) : ( n9229 ) ;
assign n9231 =  ( n8506 ) ? ( VREG_22_10 ) : ( n9230 ) ;
assign n9232 =  ( n8505 ) ? ( VREG_22_11 ) : ( n9231 ) ;
assign n9233 =  ( n8504 ) ? ( VREG_22_12 ) : ( n9232 ) ;
assign n9234 =  ( n8503 ) ? ( VREG_22_13 ) : ( n9233 ) ;
assign n9235 =  ( n8502 ) ? ( VREG_22_14 ) : ( n9234 ) ;
assign n9236 =  ( n8501 ) ? ( VREG_22_15 ) : ( n9235 ) ;
assign n9237 =  ( n8500 ) ? ( VREG_23_0 ) : ( n9236 ) ;
assign n9238 =  ( n8499 ) ? ( VREG_23_1 ) : ( n9237 ) ;
assign n9239 =  ( n8498 ) ? ( VREG_23_2 ) : ( n9238 ) ;
assign n9240 =  ( n8497 ) ? ( VREG_23_3 ) : ( n9239 ) ;
assign n9241 =  ( n8496 ) ? ( VREG_23_4 ) : ( n9240 ) ;
assign n9242 =  ( n8495 ) ? ( VREG_23_5 ) : ( n9241 ) ;
assign n9243 =  ( n8494 ) ? ( VREG_23_6 ) : ( n9242 ) ;
assign n9244 =  ( n8493 ) ? ( VREG_23_7 ) : ( n9243 ) ;
assign n9245 =  ( n8492 ) ? ( VREG_23_8 ) : ( n9244 ) ;
assign n9246 =  ( n8491 ) ? ( VREG_23_9 ) : ( n9245 ) ;
assign n9247 =  ( n8490 ) ? ( VREG_23_10 ) : ( n9246 ) ;
assign n9248 =  ( n8489 ) ? ( VREG_23_11 ) : ( n9247 ) ;
assign n9249 =  ( n8488 ) ? ( VREG_23_12 ) : ( n9248 ) ;
assign n9250 =  ( n8487 ) ? ( VREG_23_13 ) : ( n9249 ) ;
assign n9251 =  ( n8486 ) ? ( VREG_23_14 ) : ( n9250 ) ;
assign n9252 =  ( n8485 ) ? ( VREG_23_15 ) : ( n9251 ) ;
assign n9253 =  ( n8484 ) ? ( VREG_24_0 ) : ( n9252 ) ;
assign n9254 =  ( n8483 ) ? ( VREG_24_1 ) : ( n9253 ) ;
assign n9255 =  ( n8482 ) ? ( VREG_24_2 ) : ( n9254 ) ;
assign n9256 =  ( n8481 ) ? ( VREG_24_3 ) : ( n9255 ) ;
assign n9257 =  ( n8480 ) ? ( VREG_24_4 ) : ( n9256 ) ;
assign n9258 =  ( n8479 ) ? ( VREG_24_5 ) : ( n9257 ) ;
assign n9259 =  ( n8478 ) ? ( VREG_24_6 ) : ( n9258 ) ;
assign n9260 =  ( n8477 ) ? ( VREG_24_7 ) : ( n9259 ) ;
assign n9261 =  ( n8476 ) ? ( VREG_24_8 ) : ( n9260 ) ;
assign n9262 =  ( n8475 ) ? ( VREG_24_9 ) : ( n9261 ) ;
assign n9263 =  ( n8474 ) ? ( VREG_24_10 ) : ( n9262 ) ;
assign n9264 =  ( n8473 ) ? ( VREG_24_11 ) : ( n9263 ) ;
assign n9265 =  ( n8472 ) ? ( VREG_24_12 ) : ( n9264 ) ;
assign n9266 =  ( n8471 ) ? ( VREG_24_13 ) : ( n9265 ) ;
assign n9267 =  ( n8470 ) ? ( VREG_24_14 ) : ( n9266 ) ;
assign n9268 =  ( n8469 ) ? ( VREG_24_15 ) : ( n9267 ) ;
assign n9269 =  ( n8468 ) ? ( VREG_25_0 ) : ( n9268 ) ;
assign n9270 =  ( n8467 ) ? ( VREG_25_1 ) : ( n9269 ) ;
assign n9271 =  ( n8466 ) ? ( VREG_25_2 ) : ( n9270 ) ;
assign n9272 =  ( n8465 ) ? ( VREG_25_3 ) : ( n9271 ) ;
assign n9273 =  ( n8464 ) ? ( VREG_25_4 ) : ( n9272 ) ;
assign n9274 =  ( n8463 ) ? ( VREG_25_5 ) : ( n9273 ) ;
assign n9275 =  ( n8462 ) ? ( VREG_25_6 ) : ( n9274 ) ;
assign n9276 =  ( n8461 ) ? ( VREG_25_7 ) : ( n9275 ) ;
assign n9277 =  ( n8460 ) ? ( VREG_25_8 ) : ( n9276 ) ;
assign n9278 =  ( n8459 ) ? ( VREG_25_9 ) : ( n9277 ) ;
assign n9279 =  ( n8458 ) ? ( VREG_25_10 ) : ( n9278 ) ;
assign n9280 =  ( n8457 ) ? ( VREG_25_11 ) : ( n9279 ) ;
assign n9281 =  ( n8456 ) ? ( VREG_25_12 ) : ( n9280 ) ;
assign n9282 =  ( n8455 ) ? ( VREG_25_13 ) : ( n9281 ) ;
assign n9283 =  ( n8454 ) ? ( VREG_25_14 ) : ( n9282 ) ;
assign n9284 =  ( n8453 ) ? ( VREG_25_15 ) : ( n9283 ) ;
assign n9285 =  ( n8452 ) ? ( VREG_26_0 ) : ( n9284 ) ;
assign n9286 =  ( n8451 ) ? ( VREG_26_1 ) : ( n9285 ) ;
assign n9287 =  ( n8450 ) ? ( VREG_26_2 ) : ( n9286 ) ;
assign n9288 =  ( n8449 ) ? ( VREG_26_3 ) : ( n9287 ) ;
assign n9289 =  ( n8448 ) ? ( VREG_26_4 ) : ( n9288 ) ;
assign n9290 =  ( n8447 ) ? ( VREG_26_5 ) : ( n9289 ) ;
assign n9291 =  ( n8446 ) ? ( VREG_26_6 ) : ( n9290 ) ;
assign n9292 =  ( n8445 ) ? ( VREG_26_7 ) : ( n9291 ) ;
assign n9293 =  ( n8444 ) ? ( VREG_26_8 ) : ( n9292 ) ;
assign n9294 =  ( n8443 ) ? ( VREG_26_9 ) : ( n9293 ) ;
assign n9295 =  ( n8442 ) ? ( VREG_26_10 ) : ( n9294 ) ;
assign n9296 =  ( n8441 ) ? ( VREG_26_11 ) : ( n9295 ) ;
assign n9297 =  ( n8440 ) ? ( VREG_26_12 ) : ( n9296 ) ;
assign n9298 =  ( n8439 ) ? ( VREG_26_13 ) : ( n9297 ) ;
assign n9299 =  ( n8438 ) ? ( VREG_26_14 ) : ( n9298 ) ;
assign n9300 =  ( n8437 ) ? ( VREG_26_15 ) : ( n9299 ) ;
assign n9301 =  ( n8436 ) ? ( VREG_27_0 ) : ( n9300 ) ;
assign n9302 =  ( n8435 ) ? ( VREG_27_1 ) : ( n9301 ) ;
assign n9303 =  ( n8434 ) ? ( VREG_27_2 ) : ( n9302 ) ;
assign n9304 =  ( n8433 ) ? ( VREG_27_3 ) : ( n9303 ) ;
assign n9305 =  ( n8432 ) ? ( VREG_27_4 ) : ( n9304 ) ;
assign n9306 =  ( n8431 ) ? ( VREG_27_5 ) : ( n9305 ) ;
assign n9307 =  ( n8430 ) ? ( VREG_27_6 ) : ( n9306 ) ;
assign n9308 =  ( n8429 ) ? ( VREG_27_7 ) : ( n9307 ) ;
assign n9309 =  ( n8428 ) ? ( VREG_27_8 ) : ( n9308 ) ;
assign n9310 =  ( n8427 ) ? ( VREG_27_9 ) : ( n9309 ) ;
assign n9311 =  ( n8426 ) ? ( VREG_27_10 ) : ( n9310 ) ;
assign n9312 =  ( n8425 ) ? ( VREG_27_11 ) : ( n9311 ) ;
assign n9313 =  ( n8424 ) ? ( VREG_27_12 ) : ( n9312 ) ;
assign n9314 =  ( n8423 ) ? ( VREG_27_13 ) : ( n9313 ) ;
assign n9315 =  ( n8422 ) ? ( VREG_27_14 ) : ( n9314 ) ;
assign n9316 =  ( n8421 ) ? ( VREG_27_15 ) : ( n9315 ) ;
assign n9317 =  ( n8420 ) ? ( VREG_28_0 ) : ( n9316 ) ;
assign n9318 =  ( n8419 ) ? ( VREG_28_1 ) : ( n9317 ) ;
assign n9319 =  ( n8418 ) ? ( VREG_28_2 ) : ( n9318 ) ;
assign n9320 =  ( n8417 ) ? ( VREG_28_3 ) : ( n9319 ) ;
assign n9321 =  ( n8416 ) ? ( VREG_28_4 ) : ( n9320 ) ;
assign n9322 =  ( n8415 ) ? ( VREG_28_5 ) : ( n9321 ) ;
assign n9323 =  ( n8414 ) ? ( VREG_28_6 ) : ( n9322 ) ;
assign n9324 =  ( n8413 ) ? ( VREG_28_7 ) : ( n9323 ) ;
assign n9325 =  ( n8412 ) ? ( VREG_28_8 ) : ( n9324 ) ;
assign n9326 =  ( n8411 ) ? ( VREG_28_9 ) : ( n9325 ) ;
assign n9327 =  ( n8410 ) ? ( VREG_28_10 ) : ( n9326 ) ;
assign n9328 =  ( n8409 ) ? ( VREG_28_11 ) : ( n9327 ) ;
assign n9329 =  ( n8408 ) ? ( VREG_28_12 ) : ( n9328 ) ;
assign n9330 =  ( n8407 ) ? ( VREG_28_13 ) : ( n9329 ) ;
assign n9331 =  ( n8406 ) ? ( VREG_28_14 ) : ( n9330 ) ;
assign n9332 =  ( n8405 ) ? ( VREG_28_15 ) : ( n9331 ) ;
assign n9333 =  ( n8404 ) ? ( VREG_29_0 ) : ( n9332 ) ;
assign n9334 =  ( n8403 ) ? ( VREG_29_1 ) : ( n9333 ) ;
assign n9335 =  ( n8402 ) ? ( VREG_29_2 ) : ( n9334 ) ;
assign n9336 =  ( n8401 ) ? ( VREG_29_3 ) : ( n9335 ) ;
assign n9337 =  ( n8400 ) ? ( VREG_29_4 ) : ( n9336 ) ;
assign n9338 =  ( n8399 ) ? ( VREG_29_5 ) : ( n9337 ) ;
assign n9339 =  ( n8398 ) ? ( VREG_29_6 ) : ( n9338 ) ;
assign n9340 =  ( n8397 ) ? ( VREG_29_7 ) : ( n9339 ) ;
assign n9341 =  ( n8396 ) ? ( VREG_29_8 ) : ( n9340 ) ;
assign n9342 =  ( n8395 ) ? ( VREG_29_9 ) : ( n9341 ) ;
assign n9343 =  ( n8394 ) ? ( VREG_29_10 ) : ( n9342 ) ;
assign n9344 =  ( n8393 ) ? ( VREG_29_11 ) : ( n9343 ) ;
assign n9345 =  ( n8392 ) ? ( VREG_29_12 ) : ( n9344 ) ;
assign n9346 =  ( n8391 ) ? ( VREG_29_13 ) : ( n9345 ) ;
assign n9347 =  ( n8390 ) ? ( VREG_29_14 ) : ( n9346 ) ;
assign n9348 =  ( n8389 ) ? ( VREG_29_15 ) : ( n9347 ) ;
assign n9349 =  ( n8388 ) ? ( VREG_30_0 ) : ( n9348 ) ;
assign n9350 =  ( n8387 ) ? ( VREG_30_1 ) : ( n9349 ) ;
assign n9351 =  ( n8386 ) ? ( VREG_30_2 ) : ( n9350 ) ;
assign n9352 =  ( n8385 ) ? ( VREG_30_3 ) : ( n9351 ) ;
assign n9353 =  ( n8384 ) ? ( VREG_30_4 ) : ( n9352 ) ;
assign n9354 =  ( n8383 ) ? ( VREG_30_5 ) : ( n9353 ) ;
assign n9355 =  ( n8382 ) ? ( VREG_30_6 ) : ( n9354 ) ;
assign n9356 =  ( n8381 ) ? ( VREG_30_7 ) : ( n9355 ) ;
assign n9357 =  ( n8380 ) ? ( VREG_30_8 ) : ( n9356 ) ;
assign n9358 =  ( n8379 ) ? ( VREG_30_9 ) : ( n9357 ) ;
assign n9359 =  ( n8378 ) ? ( VREG_30_10 ) : ( n9358 ) ;
assign n9360 =  ( n8377 ) ? ( VREG_30_11 ) : ( n9359 ) ;
assign n9361 =  ( n8376 ) ? ( VREG_30_12 ) : ( n9360 ) ;
assign n9362 =  ( n8375 ) ? ( VREG_30_13 ) : ( n9361 ) ;
assign n9363 =  ( n8374 ) ? ( VREG_30_14 ) : ( n9362 ) ;
assign n9364 =  ( n8373 ) ? ( VREG_30_15 ) : ( n9363 ) ;
assign n9365 =  ( n8372 ) ? ( VREG_31_0 ) : ( n9364 ) ;
assign n9366 =  ( n8371 ) ? ( VREG_31_1 ) : ( n9365 ) ;
assign n9367 =  ( n8370 ) ? ( VREG_31_2 ) : ( n9366 ) ;
assign n9368 =  ( n8369 ) ? ( VREG_31_3 ) : ( n9367 ) ;
assign n9369 =  ( n8368 ) ? ( VREG_31_4 ) : ( n9368 ) ;
assign n9370 =  ( n8367 ) ? ( VREG_31_5 ) : ( n9369 ) ;
assign n9371 =  ( n8366 ) ? ( VREG_31_6 ) : ( n9370 ) ;
assign n9372 =  ( n8365 ) ? ( VREG_31_7 ) : ( n9371 ) ;
assign n9373 =  ( n8364 ) ? ( VREG_31_8 ) : ( n9372 ) ;
assign n9374 =  ( n8363 ) ? ( VREG_31_9 ) : ( n9373 ) ;
assign n9375 =  ( n8362 ) ? ( VREG_31_10 ) : ( n9374 ) ;
assign n9376 =  ( n8361 ) ? ( VREG_31_11 ) : ( n9375 ) ;
assign n9377 =  ( n8360 ) ? ( VREG_31_12 ) : ( n9376 ) ;
assign n9378 =  ( n8359 ) ? ( VREG_31_13 ) : ( n9377 ) ;
assign n9379 =  ( n8358 ) ? ( VREG_31_14 ) : ( n9378 ) ;
assign n9380 =  ( n8357 ) ? ( VREG_31_15 ) : ( n9379 ) ;
assign n9381 =  ( n8346 ) + ( n9380 )  ;
assign n9382 =  ( n8346 ) - ( n9380 )  ;
assign n9383 =  ( n8346 ) & ( n9380 )  ;
assign n9384 =  ( n8346 ) | ( n9380 )  ;
assign n9385 =  ( ( n8346 ) * ( n9380 ))  ;
assign n9386 =  ( n148 ) ? ( n9385 ) : ( VREG_0_11 ) ;
assign n9387 =  ( n146 ) ? ( n9384 ) : ( n9386 ) ;
assign n9388 =  ( n144 ) ? ( n9383 ) : ( n9387 ) ;
assign n9389 =  ( n142 ) ? ( n9382 ) : ( n9388 ) ;
assign n9390 =  ( n10 ) ? ( n9381 ) : ( n9389 ) ;
assign n9391 = n3030[11:11] ;
assign n9392 =  ( n9391 ) == ( 1'd0 )  ;
assign n9393 =  ( n9392 ) ? ( VREG_0_11 ) : ( n8356 ) ;
assign n9394 =  ( n9392 ) ? ( VREG_0_11 ) : ( n9390 ) ;
assign n9395 =  ( n3034 ) ? ( n9394 ) : ( VREG_0_11 ) ;
assign n9396 =  ( n2965 ) ? ( n9393 ) : ( n9395 ) ;
assign n9397 =  ( n1930 ) ? ( n9390 ) : ( n9396 ) ;
assign n9398 =  ( n879 ) ? ( n8356 ) : ( n9397 ) ;
assign n9399 =  ( n8346 ) + ( n164 )  ;
assign n9400 =  ( n8346 ) - ( n164 )  ;
assign n9401 =  ( n8346 ) & ( n164 )  ;
assign n9402 =  ( n8346 ) | ( n164 )  ;
assign n9403 =  ( ( n8346 ) * ( n164 ))  ;
assign n9404 =  ( n172 ) ? ( n9403 ) : ( VREG_0_11 ) ;
assign n9405 =  ( n170 ) ? ( n9402 ) : ( n9404 ) ;
assign n9406 =  ( n168 ) ? ( n9401 ) : ( n9405 ) ;
assign n9407 =  ( n166 ) ? ( n9400 ) : ( n9406 ) ;
assign n9408 =  ( n162 ) ? ( n9399 ) : ( n9407 ) ;
assign n9409 =  ( n8346 ) + ( n180 )  ;
assign n9410 =  ( n8346 ) - ( n180 )  ;
assign n9411 =  ( n8346 ) & ( n180 )  ;
assign n9412 =  ( n8346 ) | ( n180 )  ;
assign n9413 =  ( ( n8346 ) * ( n180 ))  ;
assign n9414 =  ( n172 ) ? ( n9413 ) : ( VREG_0_11 ) ;
assign n9415 =  ( n170 ) ? ( n9412 ) : ( n9414 ) ;
assign n9416 =  ( n168 ) ? ( n9411 ) : ( n9415 ) ;
assign n9417 =  ( n166 ) ? ( n9410 ) : ( n9416 ) ;
assign n9418 =  ( n162 ) ? ( n9409 ) : ( n9417 ) ;
assign n9419 =  ( n9392 ) ? ( VREG_0_11 ) : ( n9418 ) ;
assign n9420 =  ( n3051 ) ? ( n9419 ) : ( VREG_0_11 ) ;
assign n9421 =  ( n3040 ) ? ( n9408 ) : ( n9420 ) ;
assign n9422 =  ( n192 ) ? ( VREG_0_11 ) : ( VREG_0_11 ) ;
assign n9423 =  ( n157 ) ? ( n9421 ) : ( n9422 ) ;
assign n9424 =  ( n6 ) ? ( n9398 ) : ( n9423 ) ;
assign n9425 =  ( n4 ) ? ( n9424 ) : ( VREG_0_11 ) ;
assign n9426 =  ( 32'd12 ) == ( 32'd15 )  ;
assign n9427 =  ( n12 ) & ( n9426 )  ;
assign n9428 =  ( 32'd12 ) == ( 32'd14 )  ;
assign n9429 =  ( n12 ) & ( n9428 )  ;
assign n9430 =  ( 32'd12 ) == ( 32'd13 )  ;
assign n9431 =  ( n12 ) & ( n9430 )  ;
assign n9432 =  ( 32'd12 ) == ( 32'd12 )  ;
assign n9433 =  ( n12 ) & ( n9432 )  ;
assign n9434 =  ( 32'd12 ) == ( 32'd11 )  ;
assign n9435 =  ( n12 ) & ( n9434 )  ;
assign n9436 =  ( 32'd12 ) == ( 32'd10 )  ;
assign n9437 =  ( n12 ) & ( n9436 )  ;
assign n9438 =  ( 32'd12 ) == ( 32'd9 )  ;
assign n9439 =  ( n12 ) & ( n9438 )  ;
assign n9440 =  ( 32'd12 ) == ( 32'd8 )  ;
assign n9441 =  ( n12 ) & ( n9440 )  ;
assign n9442 =  ( 32'd12 ) == ( 32'd7 )  ;
assign n9443 =  ( n12 ) & ( n9442 )  ;
assign n9444 =  ( 32'd12 ) == ( 32'd6 )  ;
assign n9445 =  ( n12 ) & ( n9444 )  ;
assign n9446 =  ( 32'd12 ) == ( 32'd5 )  ;
assign n9447 =  ( n12 ) & ( n9446 )  ;
assign n9448 =  ( 32'd12 ) == ( 32'd4 )  ;
assign n9449 =  ( n12 ) & ( n9448 )  ;
assign n9450 =  ( 32'd12 ) == ( 32'd3 )  ;
assign n9451 =  ( n12 ) & ( n9450 )  ;
assign n9452 =  ( 32'd12 ) == ( 32'd2 )  ;
assign n9453 =  ( n12 ) & ( n9452 )  ;
assign n9454 =  ( 32'd12 ) == ( 32'd1 )  ;
assign n9455 =  ( n12 ) & ( n9454 )  ;
assign n9456 =  ( 32'd12 ) == ( 32'd0 )  ;
assign n9457 =  ( n12 ) & ( n9456 )  ;
assign n9458 =  ( n13 ) & ( n9426 )  ;
assign n9459 =  ( n13 ) & ( n9428 )  ;
assign n9460 =  ( n13 ) & ( n9430 )  ;
assign n9461 =  ( n13 ) & ( n9432 )  ;
assign n9462 =  ( n13 ) & ( n9434 )  ;
assign n9463 =  ( n13 ) & ( n9436 )  ;
assign n9464 =  ( n13 ) & ( n9438 )  ;
assign n9465 =  ( n13 ) & ( n9440 )  ;
assign n9466 =  ( n13 ) & ( n9442 )  ;
assign n9467 =  ( n13 ) & ( n9444 )  ;
assign n9468 =  ( n13 ) & ( n9446 )  ;
assign n9469 =  ( n13 ) & ( n9448 )  ;
assign n9470 =  ( n13 ) & ( n9450 )  ;
assign n9471 =  ( n13 ) & ( n9452 )  ;
assign n9472 =  ( n13 ) & ( n9454 )  ;
assign n9473 =  ( n13 ) & ( n9456 )  ;
assign n9474 =  ( n14 ) & ( n9426 )  ;
assign n9475 =  ( n14 ) & ( n9428 )  ;
assign n9476 =  ( n14 ) & ( n9430 )  ;
assign n9477 =  ( n14 ) & ( n9432 )  ;
assign n9478 =  ( n14 ) & ( n9434 )  ;
assign n9479 =  ( n14 ) & ( n9436 )  ;
assign n9480 =  ( n14 ) & ( n9438 )  ;
assign n9481 =  ( n14 ) & ( n9440 )  ;
assign n9482 =  ( n14 ) & ( n9442 )  ;
assign n9483 =  ( n14 ) & ( n9444 )  ;
assign n9484 =  ( n14 ) & ( n9446 )  ;
assign n9485 =  ( n14 ) & ( n9448 )  ;
assign n9486 =  ( n14 ) & ( n9450 )  ;
assign n9487 =  ( n14 ) & ( n9452 )  ;
assign n9488 =  ( n14 ) & ( n9454 )  ;
assign n9489 =  ( n14 ) & ( n9456 )  ;
assign n9490 =  ( n15 ) & ( n9426 )  ;
assign n9491 =  ( n15 ) & ( n9428 )  ;
assign n9492 =  ( n15 ) & ( n9430 )  ;
assign n9493 =  ( n15 ) & ( n9432 )  ;
assign n9494 =  ( n15 ) & ( n9434 )  ;
assign n9495 =  ( n15 ) & ( n9436 )  ;
assign n9496 =  ( n15 ) & ( n9438 )  ;
assign n9497 =  ( n15 ) & ( n9440 )  ;
assign n9498 =  ( n15 ) & ( n9442 )  ;
assign n9499 =  ( n15 ) & ( n9444 )  ;
assign n9500 =  ( n15 ) & ( n9446 )  ;
assign n9501 =  ( n15 ) & ( n9448 )  ;
assign n9502 =  ( n15 ) & ( n9450 )  ;
assign n9503 =  ( n15 ) & ( n9452 )  ;
assign n9504 =  ( n15 ) & ( n9454 )  ;
assign n9505 =  ( n15 ) & ( n9456 )  ;
assign n9506 =  ( n16 ) & ( n9426 )  ;
assign n9507 =  ( n16 ) & ( n9428 )  ;
assign n9508 =  ( n16 ) & ( n9430 )  ;
assign n9509 =  ( n16 ) & ( n9432 )  ;
assign n9510 =  ( n16 ) & ( n9434 )  ;
assign n9511 =  ( n16 ) & ( n9436 )  ;
assign n9512 =  ( n16 ) & ( n9438 )  ;
assign n9513 =  ( n16 ) & ( n9440 )  ;
assign n9514 =  ( n16 ) & ( n9442 )  ;
assign n9515 =  ( n16 ) & ( n9444 )  ;
assign n9516 =  ( n16 ) & ( n9446 )  ;
assign n9517 =  ( n16 ) & ( n9448 )  ;
assign n9518 =  ( n16 ) & ( n9450 )  ;
assign n9519 =  ( n16 ) & ( n9452 )  ;
assign n9520 =  ( n16 ) & ( n9454 )  ;
assign n9521 =  ( n16 ) & ( n9456 )  ;
assign n9522 =  ( n17 ) & ( n9426 )  ;
assign n9523 =  ( n17 ) & ( n9428 )  ;
assign n9524 =  ( n17 ) & ( n9430 )  ;
assign n9525 =  ( n17 ) & ( n9432 )  ;
assign n9526 =  ( n17 ) & ( n9434 )  ;
assign n9527 =  ( n17 ) & ( n9436 )  ;
assign n9528 =  ( n17 ) & ( n9438 )  ;
assign n9529 =  ( n17 ) & ( n9440 )  ;
assign n9530 =  ( n17 ) & ( n9442 )  ;
assign n9531 =  ( n17 ) & ( n9444 )  ;
assign n9532 =  ( n17 ) & ( n9446 )  ;
assign n9533 =  ( n17 ) & ( n9448 )  ;
assign n9534 =  ( n17 ) & ( n9450 )  ;
assign n9535 =  ( n17 ) & ( n9452 )  ;
assign n9536 =  ( n17 ) & ( n9454 )  ;
assign n9537 =  ( n17 ) & ( n9456 )  ;
assign n9538 =  ( n18 ) & ( n9426 )  ;
assign n9539 =  ( n18 ) & ( n9428 )  ;
assign n9540 =  ( n18 ) & ( n9430 )  ;
assign n9541 =  ( n18 ) & ( n9432 )  ;
assign n9542 =  ( n18 ) & ( n9434 )  ;
assign n9543 =  ( n18 ) & ( n9436 )  ;
assign n9544 =  ( n18 ) & ( n9438 )  ;
assign n9545 =  ( n18 ) & ( n9440 )  ;
assign n9546 =  ( n18 ) & ( n9442 )  ;
assign n9547 =  ( n18 ) & ( n9444 )  ;
assign n9548 =  ( n18 ) & ( n9446 )  ;
assign n9549 =  ( n18 ) & ( n9448 )  ;
assign n9550 =  ( n18 ) & ( n9450 )  ;
assign n9551 =  ( n18 ) & ( n9452 )  ;
assign n9552 =  ( n18 ) & ( n9454 )  ;
assign n9553 =  ( n18 ) & ( n9456 )  ;
assign n9554 =  ( n19 ) & ( n9426 )  ;
assign n9555 =  ( n19 ) & ( n9428 )  ;
assign n9556 =  ( n19 ) & ( n9430 )  ;
assign n9557 =  ( n19 ) & ( n9432 )  ;
assign n9558 =  ( n19 ) & ( n9434 )  ;
assign n9559 =  ( n19 ) & ( n9436 )  ;
assign n9560 =  ( n19 ) & ( n9438 )  ;
assign n9561 =  ( n19 ) & ( n9440 )  ;
assign n9562 =  ( n19 ) & ( n9442 )  ;
assign n9563 =  ( n19 ) & ( n9444 )  ;
assign n9564 =  ( n19 ) & ( n9446 )  ;
assign n9565 =  ( n19 ) & ( n9448 )  ;
assign n9566 =  ( n19 ) & ( n9450 )  ;
assign n9567 =  ( n19 ) & ( n9452 )  ;
assign n9568 =  ( n19 ) & ( n9454 )  ;
assign n9569 =  ( n19 ) & ( n9456 )  ;
assign n9570 =  ( n20 ) & ( n9426 )  ;
assign n9571 =  ( n20 ) & ( n9428 )  ;
assign n9572 =  ( n20 ) & ( n9430 )  ;
assign n9573 =  ( n20 ) & ( n9432 )  ;
assign n9574 =  ( n20 ) & ( n9434 )  ;
assign n9575 =  ( n20 ) & ( n9436 )  ;
assign n9576 =  ( n20 ) & ( n9438 )  ;
assign n9577 =  ( n20 ) & ( n9440 )  ;
assign n9578 =  ( n20 ) & ( n9442 )  ;
assign n9579 =  ( n20 ) & ( n9444 )  ;
assign n9580 =  ( n20 ) & ( n9446 )  ;
assign n9581 =  ( n20 ) & ( n9448 )  ;
assign n9582 =  ( n20 ) & ( n9450 )  ;
assign n9583 =  ( n20 ) & ( n9452 )  ;
assign n9584 =  ( n20 ) & ( n9454 )  ;
assign n9585 =  ( n20 ) & ( n9456 )  ;
assign n9586 =  ( n21 ) & ( n9426 )  ;
assign n9587 =  ( n21 ) & ( n9428 )  ;
assign n9588 =  ( n21 ) & ( n9430 )  ;
assign n9589 =  ( n21 ) & ( n9432 )  ;
assign n9590 =  ( n21 ) & ( n9434 )  ;
assign n9591 =  ( n21 ) & ( n9436 )  ;
assign n9592 =  ( n21 ) & ( n9438 )  ;
assign n9593 =  ( n21 ) & ( n9440 )  ;
assign n9594 =  ( n21 ) & ( n9442 )  ;
assign n9595 =  ( n21 ) & ( n9444 )  ;
assign n9596 =  ( n21 ) & ( n9446 )  ;
assign n9597 =  ( n21 ) & ( n9448 )  ;
assign n9598 =  ( n21 ) & ( n9450 )  ;
assign n9599 =  ( n21 ) & ( n9452 )  ;
assign n9600 =  ( n21 ) & ( n9454 )  ;
assign n9601 =  ( n21 ) & ( n9456 )  ;
assign n9602 =  ( n22 ) & ( n9426 )  ;
assign n9603 =  ( n22 ) & ( n9428 )  ;
assign n9604 =  ( n22 ) & ( n9430 )  ;
assign n9605 =  ( n22 ) & ( n9432 )  ;
assign n9606 =  ( n22 ) & ( n9434 )  ;
assign n9607 =  ( n22 ) & ( n9436 )  ;
assign n9608 =  ( n22 ) & ( n9438 )  ;
assign n9609 =  ( n22 ) & ( n9440 )  ;
assign n9610 =  ( n22 ) & ( n9442 )  ;
assign n9611 =  ( n22 ) & ( n9444 )  ;
assign n9612 =  ( n22 ) & ( n9446 )  ;
assign n9613 =  ( n22 ) & ( n9448 )  ;
assign n9614 =  ( n22 ) & ( n9450 )  ;
assign n9615 =  ( n22 ) & ( n9452 )  ;
assign n9616 =  ( n22 ) & ( n9454 )  ;
assign n9617 =  ( n22 ) & ( n9456 )  ;
assign n9618 =  ( n23 ) & ( n9426 )  ;
assign n9619 =  ( n23 ) & ( n9428 )  ;
assign n9620 =  ( n23 ) & ( n9430 )  ;
assign n9621 =  ( n23 ) & ( n9432 )  ;
assign n9622 =  ( n23 ) & ( n9434 )  ;
assign n9623 =  ( n23 ) & ( n9436 )  ;
assign n9624 =  ( n23 ) & ( n9438 )  ;
assign n9625 =  ( n23 ) & ( n9440 )  ;
assign n9626 =  ( n23 ) & ( n9442 )  ;
assign n9627 =  ( n23 ) & ( n9444 )  ;
assign n9628 =  ( n23 ) & ( n9446 )  ;
assign n9629 =  ( n23 ) & ( n9448 )  ;
assign n9630 =  ( n23 ) & ( n9450 )  ;
assign n9631 =  ( n23 ) & ( n9452 )  ;
assign n9632 =  ( n23 ) & ( n9454 )  ;
assign n9633 =  ( n23 ) & ( n9456 )  ;
assign n9634 =  ( n24 ) & ( n9426 )  ;
assign n9635 =  ( n24 ) & ( n9428 )  ;
assign n9636 =  ( n24 ) & ( n9430 )  ;
assign n9637 =  ( n24 ) & ( n9432 )  ;
assign n9638 =  ( n24 ) & ( n9434 )  ;
assign n9639 =  ( n24 ) & ( n9436 )  ;
assign n9640 =  ( n24 ) & ( n9438 )  ;
assign n9641 =  ( n24 ) & ( n9440 )  ;
assign n9642 =  ( n24 ) & ( n9442 )  ;
assign n9643 =  ( n24 ) & ( n9444 )  ;
assign n9644 =  ( n24 ) & ( n9446 )  ;
assign n9645 =  ( n24 ) & ( n9448 )  ;
assign n9646 =  ( n24 ) & ( n9450 )  ;
assign n9647 =  ( n24 ) & ( n9452 )  ;
assign n9648 =  ( n24 ) & ( n9454 )  ;
assign n9649 =  ( n24 ) & ( n9456 )  ;
assign n9650 =  ( n25 ) & ( n9426 )  ;
assign n9651 =  ( n25 ) & ( n9428 )  ;
assign n9652 =  ( n25 ) & ( n9430 )  ;
assign n9653 =  ( n25 ) & ( n9432 )  ;
assign n9654 =  ( n25 ) & ( n9434 )  ;
assign n9655 =  ( n25 ) & ( n9436 )  ;
assign n9656 =  ( n25 ) & ( n9438 )  ;
assign n9657 =  ( n25 ) & ( n9440 )  ;
assign n9658 =  ( n25 ) & ( n9442 )  ;
assign n9659 =  ( n25 ) & ( n9444 )  ;
assign n9660 =  ( n25 ) & ( n9446 )  ;
assign n9661 =  ( n25 ) & ( n9448 )  ;
assign n9662 =  ( n25 ) & ( n9450 )  ;
assign n9663 =  ( n25 ) & ( n9452 )  ;
assign n9664 =  ( n25 ) & ( n9454 )  ;
assign n9665 =  ( n25 ) & ( n9456 )  ;
assign n9666 =  ( n26 ) & ( n9426 )  ;
assign n9667 =  ( n26 ) & ( n9428 )  ;
assign n9668 =  ( n26 ) & ( n9430 )  ;
assign n9669 =  ( n26 ) & ( n9432 )  ;
assign n9670 =  ( n26 ) & ( n9434 )  ;
assign n9671 =  ( n26 ) & ( n9436 )  ;
assign n9672 =  ( n26 ) & ( n9438 )  ;
assign n9673 =  ( n26 ) & ( n9440 )  ;
assign n9674 =  ( n26 ) & ( n9442 )  ;
assign n9675 =  ( n26 ) & ( n9444 )  ;
assign n9676 =  ( n26 ) & ( n9446 )  ;
assign n9677 =  ( n26 ) & ( n9448 )  ;
assign n9678 =  ( n26 ) & ( n9450 )  ;
assign n9679 =  ( n26 ) & ( n9452 )  ;
assign n9680 =  ( n26 ) & ( n9454 )  ;
assign n9681 =  ( n26 ) & ( n9456 )  ;
assign n9682 =  ( n27 ) & ( n9426 )  ;
assign n9683 =  ( n27 ) & ( n9428 )  ;
assign n9684 =  ( n27 ) & ( n9430 )  ;
assign n9685 =  ( n27 ) & ( n9432 )  ;
assign n9686 =  ( n27 ) & ( n9434 )  ;
assign n9687 =  ( n27 ) & ( n9436 )  ;
assign n9688 =  ( n27 ) & ( n9438 )  ;
assign n9689 =  ( n27 ) & ( n9440 )  ;
assign n9690 =  ( n27 ) & ( n9442 )  ;
assign n9691 =  ( n27 ) & ( n9444 )  ;
assign n9692 =  ( n27 ) & ( n9446 )  ;
assign n9693 =  ( n27 ) & ( n9448 )  ;
assign n9694 =  ( n27 ) & ( n9450 )  ;
assign n9695 =  ( n27 ) & ( n9452 )  ;
assign n9696 =  ( n27 ) & ( n9454 )  ;
assign n9697 =  ( n27 ) & ( n9456 )  ;
assign n9698 =  ( n28 ) & ( n9426 )  ;
assign n9699 =  ( n28 ) & ( n9428 )  ;
assign n9700 =  ( n28 ) & ( n9430 )  ;
assign n9701 =  ( n28 ) & ( n9432 )  ;
assign n9702 =  ( n28 ) & ( n9434 )  ;
assign n9703 =  ( n28 ) & ( n9436 )  ;
assign n9704 =  ( n28 ) & ( n9438 )  ;
assign n9705 =  ( n28 ) & ( n9440 )  ;
assign n9706 =  ( n28 ) & ( n9442 )  ;
assign n9707 =  ( n28 ) & ( n9444 )  ;
assign n9708 =  ( n28 ) & ( n9446 )  ;
assign n9709 =  ( n28 ) & ( n9448 )  ;
assign n9710 =  ( n28 ) & ( n9450 )  ;
assign n9711 =  ( n28 ) & ( n9452 )  ;
assign n9712 =  ( n28 ) & ( n9454 )  ;
assign n9713 =  ( n28 ) & ( n9456 )  ;
assign n9714 =  ( n29 ) & ( n9426 )  ;
assign n9715 =  ( n29 ) & ( n9428 )  ;
assign n9716 =  ( n29 ) & ( n9430 )  ;
assign n9717 =  ( n29 ) & ( n9432 )  ;
assign n9718 =  ( n29 ) & ( n9434 )  ;
assign n9719 =  ( n29 ) & ( n9436 )  ;
assign n9720 =  ( n29 ) & ( n9438 )  ;
assign n9721 =  ( n29 ) & ( n9440 )  ;
assign n9722 =  ( n29 ) & ( n9442 )  ;
assign n9723 =  ( n29 ) & ( n9444 )  ;
assign n9724 =  ( n29 ) & ( n9446 )  ;
assign n9725 =  ( n29 ) & ( n9448 )  ;
assign n9726 =  ( n29 ) & ( n9450 )  ;
assign n9727 =  ( n29 ) & ( n9452 )  ;
assign n9728 =  ( n29 ) & ( n9454 )  ;
assign n9729 =  ( n29 ) & ( n9456 )  ;
assign n9730 =  ( n30 ) & ( n9426 )  ;
assign n9731 =  ( n30 ) & ( n9428 )  ;
assign n9732 =  ( n30 ) & ( n9430 )  ;
assign n9733 =  ( n30 ) & ( n9432 )  ;
assign n9734 =  ( n30 ) & ( n9434 )  ;
assign n9735 =  ( n30 ) & ( n9436 )  ;
assign n9736 =  ( n30 ) & ( n9438 )  ;
assign n9737 =  ( n30 ) & ( n9440 )  ;
assign n9738 =  ( n30 ) & ( n9442 )  ;
assign n9739 =  ( n30 ) & ( n9444 )  ;
assign n9740 =  ( n30 ) & ( n9446 )  ;
assign n9741 =  ( n30 ) & ( n9448 )  ;
assign n9742 =  ( n30 ) & ( n9450 )  ;
assign n9743 =  ( n30 ) & ( n9452 )  ;
assign n9744 =  ( n30 ) & ( n9454 )  ;
assign n9745 =  ( n30 ) & ( n9456 )  ;
assign n9746 =  ( n31 ) & ( n9426 )  ;
assign n9747 =  ( n31 ) & ( n9428 )  ;
assign n9748 =  ( n31 ) & ( n9430 )  ;
assign n9749 =  ( n31 ) & ( n9432 )  ;
assign n9750 =  ( n31 ) & ( n9434 )  ;
assign n9751 =  ( n31 ) & ( n9436 )  ;
assign n9752 =  ( n31 ) & ( n9438 )  ;
assign n9753 =  ( n31 ) & ( n9440 )  ;
assign n9754 =  ( n31 ) & ( n9442 )  ;
assign n9755 =  ( n31 ) & ( n9444 )  ;
assign n9756 =  ( n31 ) & ( n9446 )  ;
assign n9757 =  ( n31 ) & ( n9448 )  ;
assign n9758 =  ( n31 ) & ( n9450 )  ;
assign n9759 =  ( n31 ) & ( n9452 )  ;
assign n9760 =  ( n31 ) & ( n9454 )  ;
assign n9761 =  ( n31 ) & ( n9456 )  ;
assign n9762 =  ( n32 ) & ( n9426 )  ;
assign n9763 =  ( n32 ) & ( n9428 )  ;
assign n9764 =  ( n32 ) & ( n9430 )  ;
assign n9765 =  ( n32 ) & ( n9432 )  ;
assign n9766 =  ( n32 ) & ( n9434 )  ;
assign n9767 =  ( n32 ) & ( n9436 )  ;
assign n9768 =  ( n32 ) & ( n9438 )  ;
assign n9769 =  ( n32 ) & ( n9440 )  ;
assign n9770 =  ( n32 ) & ( n9442 )  ;
assign n9771 =  ( n32 ) & ( n9444 )  ;
assign n9772 =  ( n32 ) & ( n9446 )  ;
assign n9773 =  ( n32 ) & ( n9448 )  ;
assign n9774 =  ( n32 ) & ( n9450 )  ;
assign n9775 =  ( n32 ) & ( n9452 )  ;
assign n9776 =  ( n32 ) & ( n9454 )  ;
assign n9777 =  ( n32 ) & ( n9456 )  ;
assign n9778 =  ( n33 ) & ( n9426 )  ;
assign n9779 =  ( n33 ) & ( n9428 )  ;
assign n9780 =  ( n33 ) & ( n9430 )  ;
assign n9781 =  ( n33 ) & ( n9432 )  ;
assign n9782 =  ( n33 ) & ( n9434 )  ;
assign n9783 =  ( n33 ) & ( n9436 )  ;
assign n9784 =  ( n33 ) & ( n9438 )  ;
assign n9785 =  ( n33 ) & ( n9440 )  ;
assign n9786 =  ( n33 ) & ( n9442 )  ;
assign n9787 =  ( n33 ) & ( n9444 )  ;
assign n9788 =  ( n33 ) & ( n9446 )  ;
assign n9789 =  ( n33 ) & ( n9448 )  ;
assign n9790 =  ( n33 ) & ( n9450 )  ;
assign n9791 =  ( n33 ) & ( n9452 )  ;
assign n9792 =  ( n33 ) & ( n9454 )  ;
assign n9793 =  ( n33 ) & ( n9456 )  ;
assign n9794 =  ( n34 ) & ( n9426 )  ;
assign n9795 =  ( n34 ) & ( n9428 )  ;
assign n9796 =  ( n34 ) & ( n9430 )  ;
assign n9797 =  ( n34 ) & ( n9432 )  ;
assign n9798 =  ( n34 ) & ( n9434 )  ;
assign n9799 =  ( n34 ) & ( n9436 )  ;
assign n9800 =  ( n34 ) & ( n9438 )  ;
assign n9801 =  ( n34 ) & ( n9440 )  ;
assign n9802 =  ( n34 ) & ( n9442 )  ;
assign n9803 =  ( n34 ) & ( n9444 )  ;
assign n9804 =  ( n34 ) & ( n9446 )  ;
assign n9805 =  ( n34 ) & ( n9448 )  ;
assign n9806 =  ( n34 ) & ( n9450 )  ;
assign n9807 =  ( n34 ) & ( n9452 )  ;
assign n9808 =  ( n34 ) & ( n9454 )  ;
assign n9809 =  ( n34 ) & ( n9456 )  ;
assign n9810 =  ( n35 ) & ( n9426 )  ;
assign n9811 =  ( n35 ) & ( n9428 )  ;
assign n9812 =  ( n35 ) & ( n9430 )  ;
assign n9813 =  ( n35 ) & ( n9432 )  ;
assign n9814 =  ( n35 ) & ( n9434 )  ;
assign n9815 =  ( n35 ) & ( n9436 )  ;
assign n9816 =  ( n35 ) & ( n9438 )  ;
assign n9817 =  ( n35 ) & ( n9440 )  ;
assign n9818 =  ( n35 ) & ( n9442 )  ;
assign n9819 =  ( n35 ) & ( n9444 )  ;
assign n9820 =  ( n35 ) & ( n9446 )  ;
assign n9821 =  ( n35 ) & ( n9448 )  ;
assign n9822 =  ( n35 ) & ( n9450 )  ;
assign n9823 =  ( n35 ) & ( n9452 )  ;
assign n9824 =  ( n35 ) & ( n9454 )  ;
assign n9825 =  ( n35 ) & ( n9456 )  ;
assign n9826 =  ( n36 ) & ( n9426 )  ;
assign n9827 =  ( n36 ) & ( n9428 )  ;
assign n9828 =  ( n36 ) & ( n9430 )  ;
assign n9829 =  ( n36 ) & ( n9432 )  ;
assign n9830 =  ( n36 ) & ( n9434 )  ;
assign n9831 =  ( n36 ) & ( n9436 )  ;
assign n9832 =  ( n36 ) & ( n9438 )  ;
assign n9833 =  ( n36 ) & ( n9440 )  ;
assign n9834 =  ( n36 ) & ( n9442 )  ;
assign n9835 =  ( n36 ) & ( n9444 )  ;
assign n9836 =  ( n36 ) & ( n9446 )  ;
assign n9837 =  ( n36 ) & ( n9448 )  ;
assign n9838 =  ( n36 ) & ( n9450 )  ;
assign n9839 =  ( n36 ) & ( n9452 )  ;
assign n9840 =  ( n36 ) & ( n9454 )  ;
assign n9841 =  ( n36 ) & ( n9456 )  ;
assign n9842 =  ( n37 ) & ( n9426 )  ;
assign n9843 =  ( n37 ) & ( n9428 )  ;
assign n9844 =  ( n37 ) & ( n9430 )  ;
assign n9845 =  ( n37 ) & ( n9432 )  ;
assign n9846 =  ( n37 ) & ( n9434 )  ;
assign n9847 =  ( n37 ) & ( n9436 )  ;
assign n9848 =  ( n37 ) & ( n9438 )  ;
assign n9849 =  ( n37 ) & ( n9440 )  ;
assign n9850 =  ( n37 ) & ( n9442 )  ;
assign n9851 =  ( n37 ) & ( n9444 )  ;
assign n9852 =  ( n37 ) & ( n9446 )  ;
assign n9853 =  ( n37 ) & ( n9448 )  ;
assign n9854 =  ( n37 ) & ( n9450 )  ;
assign n9855 =  ( n37 ) & ( n9452 )  ;
assign n9856 =  ( n37 ) & ( n9454 )  ;
assign n9857 =  ( n37 ) & ( n9456 )  ;
assign n9858 =  ( n38 ) & ( n9426 )  ;
assign n9859 =  ( n38 ) & ( n9428 )  ;
assign n9860 =  ( n38 ) & ( n9430 )  ;
assign n9861 =  ( n38 ) & ( n9432 )  ;
assign n9862 =  ( n38 ) & ( n9434 )  ;
assign n9863 =  ( n38 ) & ( n9436 )  ;
assign n9864 =  ( n38 ) & ( n9438 )  ;
assign n9865 =  ( n38 ) & ( n9440 )  ;
assign n9866 =  ( n38 ) & ( n9442 )  ;
assign n9867 =  ( n38 ) & ( n9444 )  ;
assign n9868 =  ( n38 ) & ( n9446 )  ;
assign n9869 =  ( n38 ) & ( n9448 )  ;
assign n9870 =  ( n38 ) & ( n9450 )  ;
assign n9871 =  ( n38 ) & ( n9452 )  ;
assign n9872 =  ( n38 ) & ( n9454 )  ;
assign n9873 =  ( n38 ) & ( n9456 )  ;
assign n9874 =  ( n39 ) & ( n9426 )  ;
assign n9875 =  ( n39 ) & ( n9428 )  ;
assign n9876 =  ( n39 ) & ( n9430 )  ;
assign n9877 =  ( n39 ) & ( n9432 )  ;
assign n9878 =  ( n39 ) & ( n9434 )  ;
assign n9879 =  ( n39 ) & ( n9436 )  ;
assign n9880 =  ( n39 ) & ( n9438 )  ;
assign n9881 =  ( n39 ) & ( n9440 )  ;
assign n9882 =  ( n39 ) & ( n9442 )  ;
assign n9883 =  ( n39 ) & ( n9444 )  ;
assign n9884 =  ( n39 ) & ( n9446 )  ;
assign n9885 =  ( n39 ) & ( n9448 )  ;
assign n9886 =  ( n39 ) & ( n9450 )  ;
assign n9887 =  ( n39 ) & ( n9452 )  ;
assign n9888 =  ( n39 ) & ( n9454 )  ;
assign n9889 =  ( n39 ) & ( n9456 )  ;
assign n9890 =  ( n40 ) & ( n9426 )  ;
assign n9891 =  ( n40 ) & ( n9428 )  ;
assign n9892 =  ( n40 ) & ( n9430 )  ;
assign n9893 =  ( n40 ) & ( n9432 )  ;
assign n9894 =  ( n40 ) & ( n9434 )  ;
assign n9895 =  ( n40 ) & ( n9436 )  ;
assign n9896 =  ( n40 ) & ( n9438 )  ;
assign n9897 =  ( n40 ) & ( n9440 )  ;
assign n9898 =  ( n40 ) & ( n9442 )  ;
assign n9899 =  ( n40 ) & ( n9444 )  ;
assign n9900 =  ( n40 ) & ( n9446 )  ;
assign n9901 =  ( n40 ) & ( n9448 )  ;
assign n9902 =  ( n40 ) & ( n9450 )  ;
assign n9903 =  ( n40 ) & ( n9452 )  ;
assign n9904 =  ( n40 ) & ( n9454 )  ;
assign n9905 =  ( n40 ) & ( n9456 )  ;
assign n9906 =  ( n41 ) & ( n9426 )  ;
assign n9907 =  ( n41 ) & ( n9428 )  ;
assign n9908 =  ( n41 ) & ( n9430 )  ;
assign n9909 =  ( n41 ) & ( n9432 )  ;
assign n9910 =  ( n41 ) & ( n9434 )  ;
assign n9911 =  ( n41 ) & ( n9436 )  ;
assign n9912 =  ( n41 ) & ( n9438 )  ;
assign n9913 =  ( n41 ) & ( n9440 )  ;
assign n9914 =  ( n41 ) & ( n9442 )  ;
assign n9915 =  ( n41 ) & ( n9444 )  ;
assign n9916 =  ( n41 ) & ( n9446 )  ;
assign n9917 =  ( n41 ) & ( n9448 )  ;
assign n9918 =  ( n41 ) & ( n9450 )  ;
assign n9919 =  ( n41 ) & ( n9452 )  ;
assign n9920 =  ( n41 ) & ( n9454 )  ;
assign n9921 =  ( n41 ) & ( n9456 )  ;
assign n9922 =  ( n42 ) & ( n9426 )  ;
assign n9923 =  ( n42 ) & ( n9428 )  ;
assign n9924 =  ( n42 ) & ( n9430 )  ;
assign n9925 =  ( n42 ) & ( n9432 )  ;
assign n9926 =  ( n42 ) & ( n9434 )  ;
assign n9927 =  ( n42 ) & ( n9436 )  ;
assign n9928 =  ( n42 ) & ( n9438 )  ;
assign n9929 =  ( n42 ) & ( n9440 )  ;
assign n9930 =  ( n42 ) & ( n9442 )  ;
assign n9931 =  ( n42 ) & ( n9444 )  ;
assign n9932 =  ( n42 ) & ( n9446 )  ;
assign n9933 =  ( n42 ) & ( n9448 )  ;
assign n9934 =  ( n42 ) & ( n9450 )  ;
assign n9935 =  ( n42 ) & ( n9452 )  ;
assign n9936 =  ( n42 ) & ( n9454 )  ;
assign n9937 =  ( n42 ) & ( n9456 )  ;
assign n9938 =  ( n43 ) & ( n9426 )  ;
assign n9939 =  ( n43 ) & ( n9428 )  ;
assign n9940 =  ( n43 ) & ( n9430 )  ;
assign n9941 =  ( n43 ) & ( n9432 )  ;
assign n9942 =  ( n43 ) & ( n9434 )  ;
assign n9943 =  ( n43 ) & ( n9436 )  ;
assign n9944 =  ( n43 ) & ( n9438 )  ;
assign n9945 =  ( n43 ) & ( n9440 )  ;
assign n9946 =  ( n43 ) & ( n9442 )  ;
assign n9947 =  ( n43 ) & ( n9444 )  ;
assign n9948 =  ( n43 ) & ( n9446 )  ;
assign n9949 =  ( n43 ) & ( n9448 )  ;
assign n9950 =  ( n43 ) & ( n9450 )  ;
assign n9951 =  ( n43 ) & ( n9452 )  ;
assign n9952 =  ( n43 ) & ( n9454 )  ;
assign n9953 =  ( n43 ) & ( n9456 )  ;
assign n9954 =  ( n9953 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n9955 =  ( n9952 ) ? ( VREG_0_1 ) : ( n9954 ) ;
assign n9956 =  ( n9951 ) ? ( VREG_0_2 ) : ( n9955 ) ;
assign n9957 =  ( n9950 ) ? ( VREG_0_3 ) : ( n9956 ) ;
assign n9958 =  ( n9949 ) ? ( VREG_0_4 ) : ( n9957 ) ;
assign n9959 =  ( n9948 ) ? ( VREG_0_5 ) : ( n9958 ) ;
assign n9960 =  ( n9947 ) ? ( VREG_0_6 ) : ( n9959 ) ;
assign n9961 =  ( n9946 ) ? ( VREG_0_7 ) : ( n9960 ) ;
assign n9962 =  ( n9945 ) ? ( VREG_0_8 ) : ( n9961 ) ;
assign n9963 =  ( n9944 ) ? ( VREG_0_9 ) : ( n9962 ) ;
assign n9964 =  ( n9943 ) ? ( VREG_0_10 ) : ( n9963 ) ;
assign n9965 =  ( n9942 ) ? ( VREG_0_11 ) : ( n9964 ) ;
assign n9966 =  ( n9941 ) ? ( VREG_0_12 ) : ( n9965 ) ;
assign n9967 =  ( n9940 ) ? ( VREG_0_13 ) : ( n9966 ) ;
assign n9968 =  ( n9939 ) ? ( VREG_0_14 ) : ( n9967 ) ;
assign n9969 =  ( n9938 ) ? ( VREG_0_15 ) : ( n9968 ) ;
assign n9970 =  ( n9937 ) ? ( VREG_1_0 ) : ( n9969 ) ;
assign n9971 =  ( n9936 ) ? ( VREG_1_1 ) : ( n9970 ) ;
assign n9972 =  ( n9935 ) ? ( VREG_1_2 ) : ( n9971 ) ;
assign n9973 =  ( n9934 ) ? ( VREG_1_3 ) : ( n9972 ) ;
assign n9974 =  ( n9933 ) ? ( VREG_1_4 ) : ( n9973 ) ;
assign n9975 =  ( n9932 ) ? ( VREG_1_5 ) : ( n9974 ) ;
assign n9976 =  ( n9931 ) ? ( VREG_1_6 ) : ( n9975 ) ;
assign n9977 =  ( n9930 ) ? ( VREG_1_7 ) : ( n9976 ) ;
assign n9978 =  ( n9929 ) ? ( VREG_1_8 ) : ( n9977 ) ;
assign n9979 =  ( n9928 ) ? ( VREG_1_9 ) : ( n9978 ) ;
assign n9980 =  ( n9927 ) ? ( VREG_1_10 ) : ( n9979 ) ;
assign n9981 =  ( n9926 ) ? ( VREG_1_11 ) : ( n9980 ) ;
assign n9982 =  ( n9925 ) ? ( VREG_1_12 ) : ( n9981 ) ;
assign n9983 =  ( n9924 ) ? ( VREG_1_13 ) : ( n9982 ) ;
assign n9984 =  ( n9923 ) ? ( VREG_1_14 ) : ( n9983 ) ;
assign n9985 =  ( n9922 ) ? ( VREG_1_15 ) : ( n9984 ) ;
assign n9986 =  ( n9921 ) ? ( VREG_2_0 ) : ( n9985 ) ;
assign n9987 =  ( n9920 ) ? ( VREG_2_1 ) : ( n9986 ) ;
assign n9988 =  ( n9919 ) ? ( VREG_2_2 ) : ( n9987 ) ;
assign n9989 =  ( n9918 ) ? ( VREG_2_3 ) : ( n9988 ) ;
assign n9990 =  ( n9917 ) ? ( VREG_2_4 ) : ( n9989 ) ;
assign n9991 =  ( n9916 ) ? ( VREG_2_5 ) : ( n9990 ) ;
assign n9992 =  ( n9915 ) ? ( VREG_2_6 ) : ( n9991 ) ;
assign n9993 =  ( n9914 ) ? ( VREG_2_7 ) : ( n9992 ) ;
assign n9994 =  ( n9913 ) ? ( VREG_2_8 ) : ( n9993 ) ;
assign n9995 =  ( n9912 ) ? ( VREG_2_9 ) : ( n9994 ) ;
assign n9996 =  ( n9911 ) ? ( VREG_2_10 ) : ( n9995 ) ;
assign n9997 =  ( n9910 ) ? ( VREG_2_11 ) : ( n9996 ) ;
assign n9998 =  ( n9909 ) ? ( VREG_2_12 ) : ( n9997 ) ;
assign n9999 =  ( n9908 ) ? ( VREG_2_13 ) : ( n9998 ) ;
assign n10000 =  ( n9907 ) ? ( VREG_2_14 ) : ( n9999 ) ;
assign n10001 =  ( n9906 ) ? ( VREG_2_15 ) : ( n10000 ) ;
assign n10002 =  ( n9905 ) ? ( VREG_3_0 ) : ( n10001 ) ;
assign n10003 =  ( n9904 ) ? ( VREG_3_1 ) : ( n10002 ) ;
assign n10004 =  ( n9903 ) ? ( VREG_3_2 ) : ( n10003 ) ;
assign n10005 =  ( n9902 ) ? ( VREG_3_3 ) : ( n10004 ) ;
assign n10006 =  ( n9901 ) ? ( VREG_3_4 ) : ( n10005 ) ;
assign n10007 =  ( n9900 ) ? ( VREG_3_5 ) : ( n10006 ) ;
assign n10008 =  ( n9899 ) ? ( VREG_3_6 ) : ( n10007 ) ;
assign n10009 =  ( n9898 ) ? ( VREG_3_7 ) : ( n10008 ) ;
assign n10010 =  ( n9897 ) ? ( VREG_3_8 ) : ( n10009 ) ;
assign n10011 =  ( n9896 ) ? ( VREG_3_9 ) : ( n10010 ) ;
assign n10012 =  ( n9895 ) ? ( VREG_3_10 ) : ( n10011 ) ;
assign n10013 =  ( n9894 ) ? ( VREG_3_11 ) : ( n10012 ) ;
assign n10014 =  ( n9893 ) ? ( VREG_3_12 ) : ( n10013 ) ;
assign n10015 =  ( n9892 ) ? ( VREG_3_13 ) : ( n10014 ) ;
assign n10016 =  ( n9891 ) ? ( VREG_3_14 ) : ( n10015 ) ;
assign n10017 =  ( n9890 ) ? ( VREG_3_15 ) : ( n10016 ) ;
assign n10018 =  ( n9889 ) ? ( VREG_4_0 ) : ( n10017 ) ;
assign n10019 =  ( n9888 ) ? ( VREG_4_1 ) : ( n10018 ) ;
assign n10020 =  ( n9887 ) ? ( VREG_4_2 ) : ( n10019 ) ;
assign n10021 =  ( n9886 ) ? ( VREG_4_3 ) : ( n10020 ) ;
assign n10022 =  ( n9885 ) ? ( VREG_4_4 ) : ( n10021 ) ;
assign n10023 =  ( n9884 ) ? ( VREG_4_5 ) : ( n10022 ) ;
assign n10024 =  ( n9883 ) ? ( VREG_4_6 ) : ( n10023 ) ;
assign n10025 =  ( n9882 ) ? ( VREG_4_7 ) : ( n10024 ) ;
assign n10026 =  ( n9881 ) ? ( VREG_4_8 ) : ( n10025 ) ;
assign n10027 =  ( n9880 ) ? ( VREG_4_9 ) : ( n10026 ) ;
assign n10028 =  ( n9879 ) ? ( VREG_4_10 ) : ( n10027 ) ;
assign n10029 =  ( n9878 ) ? ( VREG_4_11 ) : ( n10028 ) ;
assign n10030 =  ( n9877 ) ? ( VREG_4_12 ) : ( n10029 ) ;
assign n10031 =  ( n9876 ) ? ( VREG_4_13 ) : ( n10030 ) ;
assign n10032 =  ( n9875 ) ? ( VREG_4_14 ) : ( n10031 ) ;
assign n10033 =  ( n9874 ) ? ( VREG_4_15 ) : ( n10032 ) ;
assign n10034 =  ( n9873 ) ? ( VREG_5_0 ) : ( n10033 ) ;
assign n10035 =  ( n9872 ) ? ( VREG_5_1 ) : ( n10034 ) ;
assign n10036 =  ( n9871 ) ? ( VREG_5_2 ) : ( n10035 ) ;
assign n10037 =  ( n9870 ) ? ( VREG_5_3 ) : ( n10036 ) ;
assign n10038 =  ( n9869 ) ? ( VREG_5_4 ) : ( n10037 ) ;
assign n10039 =  ( n9868 ) ? ( VREG_5_5 ) : ( n10038 ) ;
assign n10040 =  ( n9867 ) ? ( VREG_5_6 ) : ( n10039 ) ;
assign n10041 =  ( n9866 ) ? ( VREG_5_7 ) : ( n10040 ) ;
assign n10042 =  ( n9865 ) ? ( VREG_5_8 ) : ( n10041 ) ;
assign n10043 =  ( n9864 ) ? ( VREG_5_9 ) : ( n10042 ) ;
assign n10044 =  ( n9863 ) ? ( VREG_5_10 ) : ( n10043 ) ;
assign n10045 =  ( n9862 ) ? ( VREG_5_11 ) : ( n10044 ) ;
assign n10046 =  ( n9861 ) ? ( VREG_5_12 ) : ( n10045 ) ;
assign n10047 =  ( n9860 ) ? ( VREG_5_13 ) : ( n10046 ) ;
assign n10048 =  ( n9859 ) ? ( VREG_5_14 ) : ( n10047 ) ;
assign n10049 =  ( n9858 ) ? ( VREG_5_15 ) : ( n10048 ) ;
assign n10050 =  ( n9857 ) ? ( VREG_6_0 ) : ( n10049 ) ;
assign n10051 =  ( n9856 ) ? ( VREG_6_1 ) : ( n10050 ) ;
assign n10052 =  ( n9855 ) ? ( VREG_6_2 ) : ( n10051 ) ;
assign n10053 =  ( n9854 ) ? ( VREG_6_3 ) : ( n10052 ) ;
assign n10054 =  ( n9853 ) ? ( VREG_6_4 ) : ( n10053 ) ;
assign n10055 =  ( n9852 ) ? ( VREG_6_5 ) : ( n10054 ) ;
assign n10056 =  ( n9851 ) ? ( VREG_6_6 ) : ( n10055 ) ;
assign n10057 =  ( n9850 ) ? ( VREG_6_7 ) : ( n10056 ) ;
assign n10058 =  ( n9849 ) ? ( VREG_6_8 ) : ( n10057 ) ;
assign n10059 =  ( n9848 ) ? ( VREG_6_9 ) : ( n10058 ) ;
assign n10060 =  ( n9847 ) ? ( VREG_6_10 ) : ( n10059 ) ;
assign n10061 =  ( n9846 ) ? ( VREG_6_11 ) : ( n10060 ) ;
assign n10062 =  ( n9845 ) ? ( VREG_6_12 ) : ( n10061 ) ;
assign n10063 =  ( n9844 ) ? ( VREG_6_13 ) : ( n10062 ) ;
assign n10064 =  ( n9843 ) ? ( VREG_6_14 ) : ( n10063 ) ;
assign n10065 =  ( n9842 ) ? ( VREG_6_15 ) : ( n10064 ) ;
assign n10066 =  ( n9841 ) ? ( VREG_7_0 ) : ( n10065 ) ;
assign n10067 =  ( n9840 ) ? ( VREG_7_1 ) : ( n10066 ) ;
assign n10068 =  ( n9839 ) ? ( VREG_7_2 ) : ( n10067 ) ;
assign n10069 =  ( n9838 ) ? ( VREG_7_3 ) : ( n10068 ) ;
assign n10070 =  ( n9837 ) ? ( VREG_7_4 ) : ( n10069 ) ;
assign n10071 =  ( n9836 ) ? ( VREG_7_5 ) : ( n10070 ) ;
assign n10072 =  ( n9835 ) ? ( VREG_7_6 ) : ( n10071 ) ;
assign n10073 =  ( n9834 ) ? ( VREG_7_7 ) : ( n10072 ) ;
assign n10074 =  ( n9833 ) ? ( VREG_7_8 ) : ( n10073 ) ;
assign n10075 =  ( n9832 ) ? ( VREG_7_9 ) : ( n10074 ) ;
assign n10076 =  ( n9831 ) ? ( VREG_7_10 ) : ( n10075 ) ;
assign n10077 =  ( n9830 ) ? ( VREG_7_11 ) : ( n10076 ) ;
assign n10078 =  ( n9829 ) ? ( VREG_7_12 ) : ( n10077 ) ;
assign n10079 =  ( n9828 ) ? ( VREG_7_13 ) : ( n10078 ) ;
assign n10080 =  ( n9827 ) ? ( VREG_7_14 ) : ( n10079 ) ;
assign n10081 =  ( n9826 ) ? ( VREG_7_15 ) : ( n10080 ) ;
assign n10082 =  ( n9825 ) ? ( VREG_8_0 ) : ( n10081 ) ;
assign n10083 =  ( n9824 ) ? ( VREG_8_1 ) : ( n10082 ) ;
assign n10084 =  ( n9823 ) ? ( VREG_8_2 ) : ( n10083 ) ;
assign n10085 =  ( n9822 ) ? ( VREG_8_3 ) : ( n10084 ) ;
assign n10086 =  ( n9821 ) ? ( VREG_8_4 ) : ( n10085 ) ;
assign n10087 =  ( n9820 ) ? ( VREG_8_5 ) : ( n10086 ) ;
assign n10088 =  ( n9819 ) ? ( VREG_8_6 ) : ( n10087 ) ;
assign n10089 =  ( n9818 ) ? ( VREG_8_7 ) : ( n10088 ) ;
assign n10090 =  ( n9817 ) ? ( VREG_8_8 ) : ( n10089 ) ;
assign n10091 =  ( n9816 ) ? ( VREG_8_9 ) : ( n10090 ) ;
assign n10092 =  ( n9815 ) ? ( VREG_8_10 ) : ( n10091 ) ;
assign n10093 =  ( n9814 ) ? ( VREG_8_11 ) : ( n10092 ) ;
assign n10094 =  ( n9813 ) ? ( VREG_8_12 ) : ( n10093 ) ;
assign n10095 =  ( n9812 ) ? ( VREG_8_13 ) : ( n10094 ) ;
assign n10096 =  ( n9811 ) ? ( VREG_8_14 ) : ( n10095 ) ;
assign n10097 =  ( n9810 ) ? ( VREG_8_15 ) : ( n10096 ) ;
assign n10098 =  ( n9809 ) ? ( VREG_9_0 ) : ( n10097 ) ;
assign n10099 =  ( n9808 ) ? ( VREG_9_1 ) : ( n10098 ) ;
assign n10100 =  ( n9807 ) ? ( VREG_9_2 ) : ( n10099 ) ;
assign n10101 =  ( n9806 ) ? ( VREG_9_3 ) : ( n10100 ) ;
assign n10102 =  ( n9805 ) ? ( VREG_9_4 ) : ( n10101 ) ;
assign n10103 =  ( n9804 ) ? ( VREG_9_5 ) : ( n10102 ) ;
assign n10104 =  ( n9803 ) ? ( VREG_9_6 ) : ( n10103 ) ;
assign n10105 =  ( n9802 ) ? ( VREG_9_7 ) : ( n10104 ) ;
assign n10106 =  ( n9801 ) ? ( VREG_9_8 ) : ( n10105 ) ;
assign n10107 =  ( n9800 ) ? ( VREG_9_9 ) : ( n10106 ) ;
assign n10108 =  ( n9799 ) ? ( VREG_9_10 ) : ( n10107 ) ;
assign n10109 =  ( n9798 ) ? ( VREG_9_11 ) : ( n10108 ) ;
assign n10110 =  ( n9797 ) ? ( VREG_9_12 ) : ( n10109 ) ;
assign n10111 =  ( n9796 ) ? ( VREG_9_13 ) : ( n10110 ) ;
assign n10112 =  ( n9795 ) ? ( VREG_9_14 ) : ( n10111 ) ;
assign n10113 =  ( n9794 ) ? ( VREG_9_15 ) : ( n10112 ) ;
assign n10114 =  ( n9793 ) ? ( VREG_10_0 ) : ( n10113 ) ;
assign n10115 =  ( n9792 ) ? ( VREG_10_1 ) : ( n10114 ) ;
assign n10116 =  ( n9791 ) ? ( VREG_10_2 ) : ( n10115 ) ;
assign n10117 =  ( n9790 ) ? ( VREG_10_3 ) : ( n10116 ) ;
assign n10118 =  ( n9789 ) ? ( VREG_10_4 ) : ( n10117 ) ;
assign n10119 =  ( n9788 ) ? ( VREG_10_5 ) : ( n10118 ) ;
assign n10120 =  ( n9787 ) ? ( VREG_10_6 ) : ( n10119 ) ;
assign n10121 =  ( n9786 ) ? ( VREG_10_7 ) : ( n10120 ) ;
assign n10122 =  ( n9785 ) ? ( VREG_10_8 ) : ( n10121 ) ;
assign n10123 =  ( n9784 ) ? ( VREG_10_9 ) : ( n10122 ) ;
assign n10124 =  ( n9783 ) ? ( VREG_10_10 ) : ( n10123 ) ;
assign n10125 =  ( n9782 ) ? ( VREG_10_11 ) : ( n10124 ) ;
assign n10126 =  ( n9781 ) ? ( VREG_10_12 ) : ( n10125 ) ;
assign n10127 =  ( n9780 ) ? ( VREG_10_13 ) : ( n10126 ) ;
assign n10128 =  ( n9779 ) ? ( VREG_10_14 ) : ( n10127 ) ;
assign n10129 =  ( n9778 ) ? ( VREG_10_15 ) : ( n10128 ) ;
assign n10130 =  ( n9777 ) ? ( VREG_11_0 ) : ( n10129 ) ;
assign n10131 =  ( n9776 ) ? ( VREG_11_1 ) : ( n10130 ) ;
assign n10132 =  ( n9775 ) ? ( VREG_11_2 ) : ( n10131 ) ;
assign n10133 =  ( n9774 ) ? ( VREG_11_3 ) : ( n10132 ) ;
assign n10134 =  ( n9773 ) ? ( VREG_11_4 ) : ( n10133 ) ;
assign n10135 =  ( n9772 ) ? ( VREG_11_5 ) : ( n10134 ) ;
assign n10136 =  ( n9771 ) ? ( VREG_11_6 ) : ( n10135 ) ;
assign n10137 =  ( n9770 ) ? ( VREG_11_7 ) : ( n10136 ) ;
assign n10138 =  ( n9769 ) ? ( VREG_11_8 ) : ( n10137 ) ;
assign n10139 =  ( n9768 ) ? ( VREG_11_9 ) : ( n10138 ) ;
assign n10140 =  ( n9767 ) ? ( VREG_11_10 ) : ( n10139 ) ;
assign n10141 =  ( n9766 ) ? ( VREG_11_11 ) : ( n10140 ) ;
assign n10142 =  ( n9765 ) ? ( VREG_11_12 ) : ( n10141 ) ;
assign n10143 =  ( n9764 ) ? ( VREG_11_13 ) : ( n10142 ) ;
assign n10144 =  ( n9763 ) ? ( VREG_11_14 ) : ( n10143 ) ;
assign n10145 =  ( n9762 ) ? ( VREG_11_15 ) : ( n10144 ) ;
assign n10146 =  ( n9761 ) ? ( VREG_12_0 ) : ( n10145 ) ;
assign n10147 =  ( n9760 ) ? ( VREG_12_1 ) : ( n10146 ) ;
assign n10148 =  ( n9759 ) ? ( VREG_12_2 ) : ( n10147 ) ;
assign n10149 =  ( n9758 ) ? ( VREG_12_3 ) : ( n10148 ) ;
assign n10150 =  ( n9757 ) ? ( VREG_12_4 ) : ( n10149 ) ;
assign n10151 =  ( n9756 ) ? ( VREG_12_5 ) : ( n10150 ) ;
assign n10152 =  ( n9755 ) ? ( VREG_12_6 ) : ( n10151 ) ;
assign n10153 =  ( n9754 ) ? ( VREG_12_7 ) : ( n10152 ) ;
assign n10154 =  ( n9753 ) ? ( VREG_12_8 ) : ( n10153 ) ;
assign n10155 =  ( n9752 ) ? ( VREG_12_9 ) : ( n10154 ) ;
assign n10156 =  ( n9751 ) ? ( VREG_12_10 ) : ( n10155 ) ;
assign n10157 =  ( n9750 ) ? ( VREG_12_11 ) : ( n10156 ) ;
assign n10158 =  ( n9749 ) ? ( VREG_12_12 ) : ( n10157 ) ;
assign n10159 =  ( n9748 ) ? ( VREG_12_13 ) : ( n10158 ) ;
assign n10160 =  ( n9747 ) ? ( VREG_12_14 ) : ( n10159 ) ;
assign n10161 =  ( n9746 ) ? ( VREG_12_15 ) : ( n10160 ) ;
assign n10162 =  ( n9745 ) ? ( VREG_13_0 ) : ( n10161 ) ;
assign n10163 =  ( n9744 ) ? ( VREG_13_1 ) : ( n10162 ) ;
assign n10164 =  ( n9743 ) ? ( VREG_13_2 ) : ( n10163 ) ;
assign n10165 =  ( n9742 ) ? ( VREG_13_3 ) : ( n10164 ) ;
assign n10166 =  ( n9741 ) ? ( VREG_13_4 ) : ( n10165 ) ;
assign n10167 =  ( n9740 ) ? ( VREG_13_5 ) : ( n10166 ) ;
assign n10168 =  ( n9739 ) ? ( VREG_13_6 ) : ( n10167 ) ;
assign n10169 =  ( n9738 ) ? ( VREG_13_7 ) : ( n10168 ) ;
assign n10170 =  ( n9737 ) ? ( VREG_13_8 ) : ( n10169 ) ;
assign n10171 =  ( n9736 ) ? ( VREG_13_9 ) : ( n10170 ) ;
assign n10172 =  ( n9735 ) ? ( VREG_13_10 ) : ( n10171 ) ;
assign n10173 =  ( n9734 ) ? ( VREG_13_11 ) : ( n10172 ) ;
assign n10174 =  ( n9733 ) ? ( VREG_13_12 ) : ( n10173 ) ;
assign n10175 =  ( n9732 ) ? ( VREG_13_13 ) : ( n10174 ) ;
assign n10176 =  ( n9731 ) ? ( VREG_13_14 ) : ( n10175 ) ;
assign n10177 =  ( n9730 ) ? ( VREG_13_15 ) : ( n10176 ) ;
assign n10178 =  ( n9729 ) ? ( VREG_14_0 ) : ( n10177 ) ;
assign n10179 =  ( n9728 ) ? ( VREG_14_1 ) : ( n10178 ) ;
assign n10180 =  ( n9727 ) ? ( VREG_14_2 ) : ( n10179 ) ;
assign n10181 =  ( n9726 ) ? ( VREG_14_3 ) : ( n10180 ) ;
assign n10182 =  ( n9725 ) ? ( VREG_14_4 ) : ( n10181 ) ;
assign n10183 =  ( n9724 ) ? ( VREG_14_5 ) : ( n10182 ) ;
assign n10184 =  ( n9723 ) ? ( VREG_14_6 ) : ( n10183 ) ;
assign n10185 =  ( n9722 ) ? ( VREG_14_7 ) : ( n10184 ) ;
assign n10186 =  ( n9721 ) ? ( VREG_14_8 ) : ( n10185 ) ;
assign n10187 =  ( n9720 ) ? ( VREG_14_9 ) : ( n10186 ) ;
assign n10188 =  ( n9719 ) ? ( VREG_14_10 ) : ( n10187 ) ;
assign n10189 =  ( n9718 ) ? ( VREG_14_11 ) : ( n10188 ) ;
assign n10190 =  ( n9717 ) ? ( VREG_14_12 ) : ( n10189 ) ;
assign n10191 =  ( n9716 ) ? ( VREG_14_13 ) : ( n10190 ) ;
assign n10192 =  ( n9715 ) ? ( VREG_14_14 ) : ( n10191 ) ;
assign n10193 =  ( n9714 ) ? ( VREG_14_15 ) : ( n10192 ) ;
assign n10194 =  ( n9713 ) ? ( VREG_15_0 ) : ( n10193 ) ;
assign n10195 =  ( n9712 ) ? ( VREG_15_1 ) : ( n10194 ) ;
assign n10196 =  ( n9711 ) ? ( VREG_15_2 ) : ( n10195 ) ;
assign n10197 =  ( n9710 ) ? ( VREG_15_3 ) : ( n10196 ) ;
assign n10198 =  ( n9709 ) ? ( VREG_15_4 ) : ( n10197 ) ;
assign n10199 =  ( n9708 ) ? ( VREG_15_5 ) : ( n10198 ) ;
assign n10200 =  ( n9707 ) ? ( VREG_15_6 ) : ( n10199 ) ;
assign n10201 =  ( n9706 ) ? ( VREG_15_7 ) : ( n10200 ) ;
assign n10202 =  ( n9705 ) ? ( VREG_15_8 ) : ( n10201 ) ;
assign n10203 =  ( n9704 ) ? ( VREG_15_9 ) : ( n10202 ) ;
assign n10204 =  ( n9703 ) ? ( VREG_15_10 ) : ( n10203 ) ;
assign n10205 =  ( n9702 ) ? ( VREG_15_11 ) : ( n10204 ) ;
assign n10206 =  ( n9701 ) ? ( VREG_15_12 ) : ( n10205 ) ;
assign n10207 =  ( n9700 ) ? ( VREG_15_13 ) : ( n10206 ) ;
assign n10208 =  ( n9699 ) ? ( VREG_15_14 ) : ( n10207 ) ;
assign n10209 =  ( n9698 ) ? ( VREG_15_15 ) : ( n10208 ) ;
assign n10210 =  ( n9697 ) ? ( VREG_16_0 ) : ( n10209 ) ;
assign n10211 =  ( n9696 ) ? ( VREG_16_1 ) : ( n10210 ) ;
assign n10212 =  ( n9695 ) ? ( VREG_16_2 ) : ( n10211 ) ;
assign n10213 =  ( n9694 ) ? ( VREG_16_3 ) : ( n10212 ) ;
assign n10214 =  ( n9693 ) ? ( VREG_16_4 ) : ( n10213 ) ;
assign n10215 =  ( n9692 ) ? ( VREG_16_5 ) : ( n10214 ) ;
assign n10216 =  ( n9691 ) ? ( VREG_16_6 ) : ( n10215 ) ;
assign n10217 =  ( n9690 ) ? ( VREG_16_7 ) : ( n10216 ) ;
assign n10218 =  ( n9689 ) ? ( VREG_16_8 ) : ( n10217 ) ;
assign n10219 =  ( n9688 ) ? ( VREG_16_9 ) : ( n10218 ) ;
assign n10220 =  ( n9687 ) ? ( VREG_16_10 ) : ( n10219 ) ;
assign n10221 =  ( n9686 ) ? ( VREG_16_11 ) : ( n10220 ) ;
assign n10222 =  ( n9685 ) ? ( VREG_16_12 ) : ( n10221 ) ;
assign n10223 =  ( n9684 ) ? ( VREG_16_13 ) : ( n10222 ) ;
assign n10224 =  ( n9683 ) ? ( VREG_16_14 ) : ( n10223 ) ;
assign n10225 =  ( n9682 ) ? ( VREG_16_15 ) : ( n10224 ) ;
assign n10226 =  ( n9681 ) ? ( VREG_17_0 ) : ( n10225 ) ;
assign n10227 =  ( n9680 ) ? ( VREG_17_1 ) : ( n10226 ) ;
assign n10228 =  ( n9679 ) ? ( VREG_17_2 ) : ( n10227 ) ;
assign n10229 =  ( n9678 ) ? ( VREG_17_3 ) : ( n10228 ) ;
assign n10230 =  ( n9677 ) ? ( VREG_17_4 ) : ( n10229 ) ;
assign n10231 =  ( n9676 ) ? ( VREG_17_5 ) : ( n10230 ) ;
assign n10232 =  ( n9675 ) ? ( VREG_17_6 ) : ( n10231 ) ;
assign n10233 =  ( n9674 ) ? ( VREG_17_7 ) : ( n10232 ) ;
assign n10234 =  ( n9673 ) ? ( VREG_17_8 ) : ( n10233 ) ;
assign n10235 =  ( n9672 ) ? ( VREG_17_9 ) : ( n10234 ) ;
assign n10236 =  ( n9671 ) ? ( VREG_17_10 ) : ( n10235 ) ;
assign n10237 =  ( n9670 ) ? ( VREG_17_11 ) : ( n10236 ) ;
assign n10238 =  ( n9669 ) ? ( VREG_17_12 ) : ( n10237 ) ;
assign n10239 =  ( n9668 ) ? ( VREG_17_13 ) : ( n10238 ) ;
assign n10240 =  ( n9667 ) ? ( VREG_17_14 ) : ( n10239 ) ;
assign n10241 =  ( n9666 ) ? ( VREG_17_15 ) : ( n10240 ) ;
assign n10242 =  ( n9665 ) ? ( VREG_18_0 ) : ( n10241 ) ;
assign n10243 =  ( n9664 ) ? ( VREG_18_1 ) : ( n10242 ) ;
assign n10244 =  ( n9663 ) ? ( VREG_18_2 ) : ( n10243 ) ;
assign n10245 =  ( n9662 ) ? ( VREG_18_3 ) : ( n10244 ) ;
assign n10246 =  ( n9661 ) ? ( VREG_18_4 ) : ( n10245 ) ;
assign n10247 =  ( n9660 ) ? ( VREG_18_5 ) : ( n10246 ) ;
assign n10248 =  ( n9659 ) ? ( VREG_18_6 ) : ( n10247 ) ;
assign n10249 =  ( n9658 ) ? ( VREG_18_7 ) : ( n10248 ) ;
assign n10250 =  ( n9657 ) ? ( VREG_18_8 ) : ( n10249 ) ;
assign n10251 =  ( n9656 ) ? ( VREG_18_9 ) : ( n10250 ) ;
assign n10252 =  ( n9655 ) ? ( VREG_18_10 ) : ( n10251 ) ;
assign n10253 =  ( n9654 ) ? ( VREG_18_11 ) : ( n10252 ) ;
assign n10254 =  ( n9653 ) ? ( VREG_18_12 ) : ( n10253 ) ;
assign n10255 =  ( n9652 ) ? ( VREG_18_13 ) : ( n10254 ) ;
assign n10256 =  ( n9651 ) ? ( VREG_18_14 ) : ( n10255 ) ;
assign n10257 =  ( n9650 ) ? ( VREG_18_15 ) : ( n10256 ) ;
assign n10258 =  ( n9649 ) ? ( VREG_19_0 ) : ( n10257 ) ;
assign n10259 =  ( n9648 ) ? ( VREG_19_1 ) : ( n10258 ) ;
assign n10260 =  ( n9647 ) ? ( VREG_19_2 ) : ( n10259 ) ;
assign n10261 =  ( n9646 ) ? ( VREG_19_3 ) : ( n10260 ) ;
assign n10262 =  ( n9645 ) ? ( VREG_19_4 ) : ( n10261 ) ;
assign n10263 =  ( n9644 ) ? ( VREG_19_5 ) : ( n10262 ) ;
assign n10264 =  ( n9643 ) ? ( VREG_19_6 ) : ( n10263 ) ;
assign n10265 =  ( n9642 ) ? ( VREG_19_7 ) : ( n10264 ) ;
assign n10266 =  ( n9641 ) ? ( VREG_19_8 ) : ( n10265 ) ;
assign n10267 =  ( n9640 ) ? ( VREG_19_9 ) : ( n10266 ) ;
assign n10268 =  ( n9639 ) ? ( VREG_19_10 ) : ( n10267 ) ;
assign n10269 =  ( n9638 ) ? ( VREG_19_11 ) : ( n10268 ) ;
assign n10270 =  ( n9637 ) ? ( VREG_19_12 ) : ( n10269 ) ;
assign n10271 =  ( n9636 ) ? ( VREG_19_13 ) : ( n10270 ) ;
assign n10272 =  ( n9635 ) ? ( VREG_19_14 ) : ( n10271 ) ;
assign n10273 =  ( n9634 ) ? ( VREG_19_15 ) : ( n10272 ) ;
assign n10274 =  ( n9633 ) ? ( VREG_20_0 ) : ( n10273 ) ;
assign n10275 =  ( n9632 ) ? ( VREG_20_1 ) : ( n10274 ) ;
assign n10276 =  ( n9631 ) ? ( VREG_20_2 ) : ( n10275 ) ;
assign n10277 =  ( n9630 ) ? ( VREG_20_3 ) : ( n10276 ) ;
assign n10278 =  ( n9629 ) ? ( VREG_20_4 ) : ( n10277 ) ;
assign n10279 =  ( n9628 ) ? ( VREG_20_5 ) : ( n10278 ) ;
assign n10280 =  ( n9627 ) ? ( VREG_20_6 ) : ( n10279 ) ;
assign n10281 =  ( n9626 ) ? ( VREG_20_7 ) : ( n10280 ) ;
assign n10282 =  ( n9625 ) ? ( VREG_20_8 ) : ( n10281 ) ;
assign n10283 =  ( n9624 ) ? ( VREG_20_9 ) : ( n10282 ) ;
assign n10284 =  ( n9623 ) ? ( VREG_20_10 ) : ( n10283 ) ;
assign n10285 =  ( n9622 ) ? ( VREG_20_11 ) : ( n10284 ) ;
assign n10286 =  ( n9621 ) ? ( VREG_20_12 ) : ( n10285 ) ;
assign n10287 =  ( n9620 ) ? ( VREG_20_13 ) : ( n10286 ) ;
assign n10288 =  ( n9619 ) ? ( VREG_20_14 ) : ( n10287 ) ;
assign n10289 =  ( n9618 ) ? ( VREG_20_15 ) : ( n10288 ) ;
assign n10290 =  ( n9617 ) ? ( VREG_21_0 ) : ( n10289 ) ;
assign n10291 =  ( n9616 ) ? ( VREG_21_1 ) : ( n10290 ) ;
assign n10292 =  ( n9615 ) ? ( VREG_21_2 ) : ( n10291 ) ;
assign n10293 =  ( n9614 ) ? ( VREG_21_3 ) : ( n10292 ) ;
assign n10294 =  ( n9613 ) ? ( VREG_21_4 ) : ( n10293 ) ;
assign n10295 =  ( n9612 ) ? ( VREG_21_5 ) : ( n10294 ) ;
assign n10296 =  ( n9611 ) ? ( VREG_21_6 ) : ( n10295 ) ;
assign n10297 =  ( n9610 ) ? ( VREG_21_7 ) : ( n10296 ) ;
assign n10298 =  ( n9609 ) ? ( VREG_21_8 ) : ( n10297 ) ;
assign n10299 =  ( n9608 ) ? ( VREG_21_9 ) : ( n10298 ) ;
assign n10300 =  ( n9607 ) ? ( VREG_21_10 ) : ( n10299 ) ;
assign n10301 =  ( n9606 ) ? ( VREG_21_11 ) : ( n10300 ) ;
assign n10302 =  ( n9605 ) ? ( VREG_21_12 ) : ( n10301 ) ;
assign n10303 =  ( n9604 ) ? ( VREG_21_13 ) : ( n10302 ) ;
assign n10304 =  ( n9603 ) ? ( VREG_21_14 ) : ( n10303 ) ;
assign n10305 =  ( n9602 ) ? ( VREG_21_15 ) : ( n10304 ) ;
assign n10306 =  ( n9601 ) ? ( VREG_22_0 ) : ( n10305 ) ;
assign n10307 =  ( n9600 ) ? ( VREG_22_1 ) : ( n10306 ) ;
assign n10308 =  ( n9599 ) ? ( VREG_22_2 ) : ( n10307 ) ;
assign n10309 =  ( n9598 ) ? ( VREG_22_3 ) : ( n10308 ) ;
assign n10310 =  ( n9597 ) ? ( VREG_22_4 ) : ( n10309 ) ;
assign n10311 =  ( n9596 ) ? ( VREG_22_5 ) : ( n10310 ) ;
assign n10312 =  ( n9595 ) ? ( VREG_22_6 ) : ( n10311 ) ;
assign n10313 =  ( n9594 ) ? ( VREG_22_7 ) : ( n10312 ) ;
assign n10314 =  ( n9593 ) ? ( VREG_22_8 ) : ( n10313 ) ;
assign n10315 =  ( n9592 ) ? ( VREG_22_9 ) : ( n10314 ) ;
assign n10316 =  ( n9591 ) ? ( VREG_22_10 ) : ( n10315 ) ;
assign n10317 =  ( n9590 ) ? ( VREG_22_11 ) : ( n10316 ) ;
assign n10318 =  ( n9589 ) ? ( VREG_22_12 ) : ( n10317 ) ;
assign n10319 =  ( n9588 ) ? ( VREG_22_13 ) : ( n10318 ) ;
assign n10320 =  ( n9587 ) ? ( VREG_22_14 ) : ( n10319 ) ;
assign n10321 =  ( n9586 ) ? ( VREG_22_15 ) : ( n10320 ) ;
assign n10322 =  ( n9585 ) ? ( VREG_23_0 ) : ( n10321 ) ;
assign n10323 =  ( n9584 ) ? ( VREG_23_1 ) : ( n10322 ) ;
assign n10324 =  ( n9583 ) ? ( VREG_23_2 ) : ( n10323 ) ;
assign n10325 =  ( n9582 ) ? ( VREG_23_3 ) : ( n10324 ) ;
assign n10326 =  ( n9581 ) ? ( VREG_23_4 ) : ( n10325 ) ;
assign n10327 =  ( n9580 ) ? ( VREG_23_5 ) : ( n10326 ) ;
assign n10328 =  ( n9579 ) ? ( VREG_23_6 ) : ( n10327 ) ;
assign n10329 =  ( n9578 ) ? ( VREG_23_7 ) : ( n10328 ) ;
assign n10330 =  ( n9577 ) ? ( VREG_23_8 ) : ( n10329 ) ;
assign n10331 =  ( n9576 ) ? ( VREG_23_9 ) : ( n10330 ) ;
assign n10332 =  ( n9575 ) ? ( VREG_23_10 ) : ( n10331 ) ;
assign n10333 =  ( n9574 ) ? ( VREG_23_11 ) : ( n10332 ) ;
assign n10334 =  ( n9573 ) ? ( VREG_23_12 ) : ( n10333 ) ;
assign n10335 =  ( n9572 ) ? ( VREG_23_13 ) : ( n10334 ) ;
assign n10336 =  ( n9571 ) ? ( VREG_23_14 ) : ( n10335 ) ;
assign n10337 =  ( n9570 ) ? ( VREG_23_15 ) : ( n10336 ) ;
assign n10338 =  ( n9569 ) ? ( VREG_24_0 ) : ( n10337 ) ;
assign n10339 =  ( n9568 ) ? ( VREG_24_1 ) : ( n10338 ) ;
assign n10340 =  ( n9567 ) ? ( VREG_24_2 ) : ( n10339 ) ;
assign n10341 =  ( n9566 ) ? ( VREG_24_3 ) : ( n10340 ) ;
assign n10342 =  ( n9565 ) ? ( VREG_24_4 ) : ( n10341 ) ;
assign n10343 =  ( n9564 ) ? ( VREG_24_5 ) : ( n10342 ) ;
assign n10344 =  ( n9563 ) ? ( VREG_24_6 ) : ( n10343 ) ;
assign n10345 =  ( n9562 ) ? ( VREG_24_7 ) : ( n10344 ) ;
assign n10346 =  ( n9561 ) ? ( VREG_24_8 ) : ( n10345 ) ;
assign n10347 =  ( n9560 ) ? ( VREG_24_9 ) : ( n10346 ) ;
assign n10348 =  ( n9559 ) ? ( VREG_24_10 ) : ( n10347 ) ;
assign n10349 =  ( n9558 ) ? ( VREG_24_11 ) : ( n10348 ) ;
assign n10350 =  ( n9557 ) ? ( VREG_24_12 ) : ( n10349 ) ;
assign n10351 =  ( n9556 ) ? ( VREG_24_13 ) : ( n10350 ) ;
assign n10352 =  ( n9555 ) ? ( VREG_24_14 ) : ( n10351 ) ;
assign n10353 =  ( n9554 ) ? ( VREG_24_15 ) : ( n10352 ) ;
assign n10354 =  ( n9553 ) ? ( VREG_25_0 ) : ( n10353 ) ;
assign n10355 =  ( n9552 ) ? ( VREG_25_1 ) : ( n10354 ) ;
assign n10356 =  ( n9551 ) ? ( VREG_25_2 ) : ( n10355 ) ;
assign n10357 =  ( n9550 ) ? ( VREG_25_3 ) : ( n10356 ) ;
assign n10358 =  ( n9549 ) ? ( VREG_25_4 ) : ( n10357 ) ;
assign n10359 =  ( n9548 ) ? ( VREG_25_5 ) : ( n10358 ) ;
assign n10360 =  ( n9547 ) ? ( VREG_25_6 ) : ( n10359 ) ;
assign n10361 =  ( n9546 ) ? ( VREG_25_7 ) : ( n10360 ) ;
assign n10362 =  ( n9545 ) ? ( VREG_25_8 ) : ( n10361 ) ;
assign n10363 =  ( n9544 ) ? ( VREG_25_9 ) : ( n10362 ) ;
assign n10364 =  ( n9543 ) ? ( VREG_25_10 ) : ( n10363 ) ;
assign n10365 =  ( n9542 ) ? ( VREG_25_11 ) : ( n10364 ) ;
assign n10366 =  ( n9541 ) ? ( VREG_25_12 ) : ( n10365 ) ;
assign n10367 =  ( n9540 ) ? ( VREG_25_13 ) : ( n10366 ) ;
assign n10368 =  ( n9539 ) ? ( VREG_25_14 ) : ( n10367 ) ;
assign n10369 =  ( n9538 ) ? ( VREG_25_15 ) : ( n10368 ) ;
assign n10370 =  ( n9537 ) ? ( VREG_26_0 ) : ( n10369 ) ;
assign n10371 =  ( n9536 ) ? ( VREG_26_1 ) : ( n10370 ) ;
assign n10372 =  ( n9535 ) ? ( VREG_26_2 ) : ( n10371 ) ;
assign n10373 =  ( n9534 ) ? ( VREG_26_3 ) : ( n10372 ) ;
assign n10374 =  ( n9533 ) ? ( VREG_26_4 ) : ( n10373 ) ;
assign n10375 =  ( n9532 ) ? ( VREG_26_5 ) : ( n10374 ) ;
assign n10376 =  ( n9531 ) ? ( VREG_26_6 ) : ( n10375 ) ;
assign n10377 =  ( n9530 ) ? ( VREG_26_7 ) : ( n10376 ) ;
assign n10378 =  ( n9529 ) ? ( VREG_26_8 ) : ( n10377 ) ;
assign n10379 =  ( n9528 ) ? ( VREG_26_9 ) : ( n10378 ) ;
assign n10380 =  ( n9527 ) ? ( VREG_26_10 ) : ( n10379 ) ;
assign n10381 =  ( n9526 ) ? ( VREG_26_11 ) : ( n10380 ) ;
assign n10382 =  ( n9525 ) ? ( VREG_26_12 ) : ( n10381 ) ;
assign n10383 =  ( n9524 ) ? ( VREG_26_13 ) : ( n10382 ) ;
assign n10384 =  ( n9523 ) ? ( VREG_26_14 ) : ( n10383 ) ;
assign n10385 =  ( n9522 ) ? ( VREG_26_15 ) : ( n10384 ) ;
assign n10386 =  ( n9521 ) ? ( VREG_27_0 ) : ( n10385 ) ;
assign n10387 =  ( n9520 ) ? ( VREG_27_1 ) : ( n10386 ) ;
assign n10388 =  ( n9519 ) ? ( VREG_27_2 ) : ( n10387 ) ;
assign n10389 =  ( n9518 ) ? ( VREG_27_3 ) : ( n10388 ) ;
assign n10390 =  ( n9517 ) ? ( VREG_27_4 ) : ( n10389 ) ;
assign n10391 =  ( n9516 ) ? ( VREG_27_5 ) : ( n10390 ) ;
assign n10392 =  ( n9515 ) ? ( VREG_27_6 ) : ( n10391 ) ;
assign n10393 =  ( n9514 ) ? ( VREG_27_7 ) : ( n10392 ) ;
assign n10394 =  ( n9513 ) ? ( VREG_27_8 ) : ( n10393 ) ;
assign n10395 =  ( n9512 ) ? ( VREG_27_9 ) : ( n10394 ) ;
assign n10396 =  ( n9511 ) ? ( VREG_27_10 ) : ( n10395 ) ;
assign n10397 =  ( n9510 ) ? ( VREG_27_11 ) : ( n10396 ) ;
assign n10398 =  ( n9509 ) ? ( VREG_27_12 ) : ( n10397 ) ;
assign n10399 =  ( n9508 ) ? ( VREG_27_13 ) : ( n10398 ) ;
assign n10400 =  ( n9507 ) ? ( VREG_27_14 ) : ( n10399 ) ;
assign n10401 =  ( n9506 ) ? ( VREG_27_15 ) : ( n10400 ) ;
assign n10402 =  ( n9505 ) ? ( VREG_28_0 ) : ( n10401 ) ;
assign n10403 =  ( n9504 ) ? ( VREG_28_1 ) : ( n10402 ) ;
assign n10404 =  ( n9503 ) ? ( VREG_28_2 ) : ( n10403 ) ;
assign n10405 =  ( n9502 ) ? ( VREG_28_3 ) : ( n10404 ) ;
assign n10406 =  ( n9501 ) ? ( VREG_28_4 ) : ( n10405 ) ;
assign n10407 =  ( n9500 ) ? ( VREG_28_5 ) : ( n10406 ) ;
assign n10408 =  ( n9499 ) ? ( VREG_28_6 ) : ( n10407 ) ;
assign n10409 =  ( n9498 ) ? ( VREG_28_7 ) : ( n10408 ) ;
assign n10410 =  ( n9497 ) ? ( VREG_28_8 ) : ( n10409 ) ;
assign n10411 =  ( n9496 ) ? ( VREG_28_9 ) : ( n10410 ) ;
assign n10412 =  ( n9495 ) ? ( VREG_28_10 ) : ( n10411 ) ;
assign n10413 =  ( n9494 ) ? ( VREG_28_11 ) : ( n10412 ) ;
assign n10414 =  ( n9493 ) ? ( VREG_28_12 ) : ( n10413 ) ;
assign n10415 =  ( n9492 ) ? ( VREG_28_13 ) : ( n10414 ) ;
assign n10416 =  ( n9491 ) ? ( VREG_28_14 ) : ( n10415 ) ;
assign n10417 =  ( n9490 ) ? ( VREG_28_15 ) : ( n10416 ) ;
assign n10418 =  ( n9489 ) ? ( VREG_29_0 ) : ( n10417 ) ;
assign n10419 =  ( n9488 ) ? ( VREG_29_1 ) : ( n10418 ) ;
assign n10420 =  ( n9487 ) ? ( VREG_29_2 ) : ( n10419 ) ;
assign n10421 =  ( n9486 ) ? ( VREG_29_3 ) : ( n10420 ) ;
assign n10422 =  ( n9485 ) ? ( VREG_29_4 ) : ( n10421 ) ;
assign n10423 =  ( n9484 ) ? ( VREG_29_5 ) : ( n10422 ) ;
assign n10424 =  ( n9483 ) ? ( VREG_29_6 ) : ( n10423 ) ;
assign n10425 =  ( n9482 ) ? ( VREG_29_7 ) : ( n10424 ) ;
assign n10426 =  ( n9481 ) ? ( VREG_29_8 ) : ( n10425 ) ;
assign n10427 =  ( n9480 ) ? ( VREG_29_9 ) : ( n10426 ) ;
assign n10428 =  ( n9479 ) ? ( VREG_29_10 ) : ( n10427 ) ;
assign n10429 =  ( n9478 ) ? ( VREG_29_11 ) : ( n10428 ) ;
assign n10430 =  ( n9477 ) ? ( VREG_29_12 ) : ( n10429 ) ;
assign n10431 =  ( n9476 ) ? ( VREG_29_13 ) : ( n10430 ) ;
assign n10432 =  ( n9475 ) ? ( VREG_29_14 ) : ( n10431 ) ;
assign n10433 =  ( n9474 ) ? ( VREG_29_15 ) : ( n10432 ) ;
assign n10434 =  ( n9473 ) ? ( VREG_30_0 ) : ( n10433 ) ;
assign n10435 =  ( n9472 ) ? ( VREG_30_1 ) : ( n10434 ) ;
assign n10436 =  ( n9471 ) ? ( VREG_30_2 ) : ( n10435 ) ;
assign n10437 =  ( n9470 ) ? ( VREG_30_3 ) : ( n10436 ) ;
assign n10438 =  ( n9469 ) ? ( VREG_30_4 ) : ( n10437 ) ;
assign n10439 =  ( n9468 ) ? ( VREG_30_5 ) : ( n10438 ) ;
assign n10440 =  ( n9467 ) ? ( VREG_30_6 ) : ( n10439 ) ;
assign n10441 =  ( n9466 ) ? ( VREG_30_7 ) : ( n10440 ) ;
assign n10442 =  ( n9465 ) ? ( VREG_30_8 ) : ( n10441 ) ;
assign n10443 =  ( n9464 ) ? ( VREG_30_9 ) : ( n10442 ) ;
assign n10444 =  ( n9463 ) ? ( VREG_30_10 ) : ( n10443 ) ;
assign n10445 =  ( n9462 ) ? ( VREG_30_11 ) : ( n10444 ) ;
assign n10446 =  ( n9461 ) ? ( VREG_30_12 ) : ( n10445 ) ;
assign n10447 =  ( n9460 ) ? ( VREG_30_13 ) : ( n10446 ) ;
assign n10448 =  ( n9459 ) ? ( VREG_30_14 ) : ( n10447 ) ;
assign n10449 =  ( n9458 ) ? ( VREG_30_15 ) : ( n10448 ) ;
assign n10450 =  ( n9457 ) ? ( VREG_31_0 ) : ( n10449 ) ;
assign n10451 =  ( n9455 ) ? ( VREG_31_1 ) : ( n10450 ) ;
assign n10452 =  ( n9453 ) ? ( VREG_31_2 ) : ( n10451 ) ;
assign n10453 =  ( n9451 ) ? ( VREG_31_3 ) : ( n10452 ) ;
assign n10454 =  ( n9449 ) ? ( VREG_31_4 ) : ( n10453 ) ;
assign n10455 =  ( n9447 ) ? ( VREG_31_5 ) : ( n10454 ) ;
assign n10456 =  ( n9445 ) ? ( VREG_31_6 ) : ( n10455 ) ;
assign n10457 =  ( n9443 ) ? ( VREG_31_7 ) : ( n10456 ) ;
assign n10458 =  ( n9441 ) ? ( VREG_31_8 ) : ( n10457 ) ;
assign n10459 =  ( n9439 ) ? ( VREG_31_9 ) : ( n10458 ) ;
assign n10460 =  ( n9437 ) ? ( VREG_31_10 ) : ( n10459 ) ;
assign n10461 =  ( n9435 ) ? ( VREG_31_11 ) : ( n10460 ) ;
assign n10462 =  ( n9433 ) ? ( VREG_31_12 ) : ( n10461 ) ;
assign n10463 =  ( n9431 ) ? ( VREG_31_13 ) : ( n10462 ) ;
assign n10464 =  ( n9429 ) ? ( VREG_31_14 ) : ( n10463 ) ;
assign n10465 =  ( n9427 ) ? ( VREG_31_15 ) : ( n10464 ) ;
assign n10466 =  ( n10465 ) + ( n140 )  ;
assign n10467 =  ( n10465 ) - ( n140 )  ;
assign n10468 =  ( n10465 ) & ( n140 )  ;
assign n10469 =  ( n10465 ) | ( n140 )  ;
assign n10470 =  ( ( n10465 ) * ( n140 ))  ;
assign n10471 =  ( n148 ) ? ( n10470 ) : ( VREG_0_12 ) ;
assign n10472 =  ( n146 ) ? ( n10469 ) : ( n10471 ) ;
assign n10473 =  ( n144 ) ? ( n10468 ) : ( n10472 ) ;
assign n10474 =  ( n142 ) ? ( n10467 ) : ( n10473 ) ;
assign n10475 =  ( n10 ) ? ( n10466 ) : ( n10474 ) ;
assign n10476 =  ( n77 ) & ( n9426 )  ;
assign n10477 =  ( n77 ) & ( n9428 )  ;
assign n10478 =  ( n77 ) & ( n9430 )  ;
assign n10479 =  ( n77 ) & ( n9432 )  ;
assign n10480 =  ( n77 ) & ( n9434 )  ;
assign n10481 =  ( n77 ) & ( n9436 )  ;
assign n10482 =  ( n77 ) & ( n9438 )  ;
assign n10483 =  ( n77 ) & ( n9440 )  ;
assign n10484 =  ( n77 ) & ( n9442 )  ;
assign n10485 =  ( n77 ) & ( n9444 )  ;
assign n10486 =  ( n77 ) & ( n9446 )  ;
assign n10487 =  ( n77 ) & ( n9448 )  ;
assign n10488 =  ( n77 ) & ( n9450 )  ;
assign n10489 =  ( n77 ) & ( n9452 )  ;
assign n10490 =  ( n77 ) & ( n9454 )  ;
assign n10491 =  ( n77 ) & ( n9456 )  ;
assign n10492 =  ( n78 ) & ( n9426 )  ;
assign n10493 =  ( n78 ) & ( n9428 )  ;
assign n10494 =  ( n78 ) & ( n9430 )  ;
assign n10495 =  ( n78 ) & ( n9432 )  ;
assign n10496 =  ( n78 ) & ( n9434 )  ;
assign n10497 =  ( n78 ) & ( n9436 )  ;
assign n10498 =  ( n78 ) & ( n9438 )  ;
assign n10499 =  ( n78 ) & ( n9440 )  ;
assign n10500 =  ( n78 ) & ( n9442 )  ;
assign n10501 =  ( n78 ) & ( n9444 )  ;
assign n10502 =  ( n78 ) & ( n9446 )  ;
assign n10503 =  ( n78 ) & ( n9448 )  ;
assign n10504 =  ( n78 ) & ( n9450 )  ;
assign n10505 =  ( n78 ) & ( n9452 )  ;
assign n10506 =  ( n78 ) & ( n9454 )  ;
assign n10507 =  ( n78 ) & ( n9456 )  ;
assign n10508 =  ( n79 ) & ( n9426 )  ;
assign n10509 =  ( n79 ) & ( n9428 )  ;
assign n10510 =  ( n79 ) & ( n9430 )  ;
assign n10511 =  ( n79 ) & ( n9432 )  ;
assign n10512 =  ( n79 ) & ( n9434 )  ;
assign n10513 =  ( n79 ) & ( n9436 )  ;
assign n10514 =  ( n79 ) & ( n9438 )  ;
assign n10515 =  ( n79 ) & ( n9440 )  ;
assign n10516 =  ( n79 ) & ( n9442 )  ;
assign n10517 =  ( n79 ) & ( n9444 )  ;
assign n10518 =  ( n79 ) & ( n9446 )  ;
assign n10519 =  ( n79 ) & ( n9448 )  ;
assign n10520 =  ( n79 ) & ( n9450 )  ;
assign n10521 =  ( n79 ) & ( n9452 )  ;
assign n10522 =  ( n79 ) & ( n9454 )  ;
assign n10523 =  ( n79 ) & ( n9456 )  ;
assign n10524 =  ( n80 ) & ( n9426 )  ;
assign n10525 =  ( n80 ) & ( n9428 )  ;
assign n10526 =  ( n80 ) & ( n9430 )  ;
assign n10527 =  ( n80 ) & ( n9432 )  ;
assign n10528 =  ( n80 ) & ( n9434 )  ;
assign n10529 =  ( n80 ) & ( n9436 )  ;
assign n10530 =  ( n80 ) & ( n9438 )  ;
assign n10531 =  ( n80 ) & ( n9440 )  ;
assign n10532 =  ( n80 ) & ( n9442 )  ;
assign n10533 =  ( n80 ) & ( n9444 )  ;
assign n10534 =  ( n80 ) & ( n9446 )  ;
assign n10535 =  ( n80 ) & ( n9448 )  ;
assign n10536 =  ( n80 ) & ( n9450 )  ;
assign n10537 =  ( n80 ) & ( n9452 )  ;
assign n10538 =  ( n80 ) & ( n9454 )  ;
assign n10539 =  ( n80 ) & ( n9456 )  ;
assign n10540 =  ( n81 ) & ( n9426 )  ;
assign n10541 =  ( n81 ) & ( n9428 )  ;
assign n10542 =  ( n81 ) & ( n9430 )  ;
assign n10543 =  ( n81 ) & ( n9432 )  ;
assign n10544 =  ( n81 ) & ( n9434 )  ;
assign n10545 =  ( n81 ) & ( n9436 )  ;
assign n10546 =  ( n81 ) & ( n9438 )  ;
assign n10547 =  ( n81 ) & ( n9440 )  ;
assign n10548 =  ( n81 ) & ( n9442 )  ;
assign n10549 =  ( n81 ) & ( n9444 )  ;
assign n10550 =  ( n81 ) & ( n9446 )  ;
assign n10551 =  ( n81 ) & ( n9448 )  ;
assign n10552 =  ( n81 ) & ( n9450 )  ;
assign n10553 =  ( n81 ) & ( n9452 )  ;
assign n10554 =  ( n81 ) & ( n9454 )  ;
assign n10555 =  ( n81 ) & ( n9456 )  ;
assign n10556 =  ( n82 ) & ( n9426 )  ;
assign n10557 =  ( n82 ) & ( n9428 )  ;
assign n10558 =  ( n82 ) & ( n9430 )  ;
assign n10559 =  ( n82 ) & ( n9432 )  ;
assign n10560 =  ( n82 ) & ( n9434 )  ;
assign n10561 =  ( n82 ) & ( n9436 )  ;
assign n10562 =  ( n82 ) & ( n9438 )  ;
assign n10563 =  ( n82 ) & ( n9440 )  ;
assign n10564 =  ( n82 ) & ( n9442 )  ;
assign n10565 =  ( n82 ) & ( n9444 )  ;
assign n10566 =  ( n82 ) & ( n9446 )  ;
assign n10567 =  ( n82 ) & ( n9448 )  ;
assign n10568 =  ( n82 ) & ( n9450 )  ;
assign n10569 =  ( n82 ) & ( n9452 )  ;
assign n10570 =  ( n82 ) & ( n9454 )  ;
assign n10571 =  ( n82 ) & ( n9456 )  ;
assign n10572 =  ( n83 ) & ( n9426 )  ;
assign n10573 =  ( n83 ) & ( n9428 )  ;
assign n10574 =  ( n83 ) & ( n9430 )  ;
assign n10575 =  ( n83 ) & ( n9432 )  ;
assign n10576 =  ( n83 ) & ( n9434 )  ;
assign n10577 =  ( n83 ) & ( n9436 )  ;
assign n10578 =  ( n83 ) & ( n9438 )  ;
assign n10579 =  ( n83 ) & ( n9440 )  ;
assign n10580 =  ( n83 ) & ( n9442 )  ;
assign n10581 =  ( n83 ) & ( n9444 )  ;
assign n10582 =  ( n83 ) & ( n9446 )  ;
assign n10583 =  ( n83 ) & ( n9448 )  ;
assign n10584 =  ( n83 ) & ( n9450 )  ;
assign n10585 =  ( n83 ) & ( n9452 )  ;
assign n10586 =  ( n83 ) & ( n9454 )  ;
assign n10587 =  ( n83 ) & ( n9456 )  ;
assign n10588 =  ( n84 ) & ( n9426 )  ;
assign n10589 =  ( n84 ) & ( n9428 )  ;
assign n10590 =  ( n84 ) & ( n9430 )  ;
assign n10591 =  ( n84 ) & ( n9432 )  ;
assign n10592 =  ( n84 ) & ( n9434 )  ;
assign n10593 =  ( n84 ) & ( n9436 )  ;
assign n10594 =  ( n84 ) & ( n9438 )  ;
assign n10595 =  ( n84 ) & ( n9440 )  ;
assign n10596 =  ( n84 ) & ( n9442 )  ;
assign n10597 =  ( n84 ) & ( n9444 )  ;
assign n10598 =  ( n84 ) & ( n9446 )  ;
assign n10599 =  ( n84 ) & ( n9448 )  ;
assign n10600 =  ( n84 ) & ( n9450 )  ;
assign n10601 =  ( n84 ) & ( n9452 )  ;
assign n10602 =  ( n84 ) & ( n9454 )  ;
assign n10603 =  ( n84 ) & ( n9456 )  ;
assign n10604 =  ( n85 ) & ( n9426 )  ;
assign n10605 =  ( n85 ) & ( n9428 )  ;
assign n10606 =  ( n85 ) & ( n9430 )  ;
assign n10607 =  ( n85 ) & ( n9432 )  ;
assign n10608 =  ( n85 ) & ( n9434 )  ;
assign n10609 =  ( n85 ) & ( n9436 )  ;
assign n10610 =  ( n85 ) & ( n9438 )  ;
assign n10611 =  ( n85 ) & ( n9440 )  ;
assign n10612 =  ( n85 ) & ( n9442 )  ;
assign n10613 =  ( n85 ) & ( n9444 )  ;
assign n10614 =  ( n85 ) & ( n9446 )  ;
assign n10615 =  ( n85 ) & ( n9448 )  ;
assign n10616 =  ( n85 ) & ( n9450 )  ;
assign n10617 =  ( n85 ) & ( n9452 )  ;
assign n10618 =  ( n85 ) & ( n9454 )  ;
assign n10619 =  ( n85 ) & ( n9456 )  ;
assign n10620 =  ( n86 ) & ( n9426 )  ;
assign n10621 =  ( n86 ) & ( n9428 )  ;
assign n10622 =  ( n86 ) & ( n9430 )  ;
assign n10623 =  ( n86 ) & ( n9432 )  ;
assign n10624 =  ( n86 ) & ( n9434 )  ;
assign n10625 =  ( n86 ) & ( n9436 )  ;
assign n10626 =  ( n86 ) & ( n9438 )  ;
assign n10627 =  ( n86 ) & ( n9440 )  ;
assign n10628 =  ( n86 ) & ( n9442 )  ;
assign n10629 =  ( n86 ) & ( n9444 )  ;
assign n10630 =  ( n86 ) & ( n9446 )  ;
assign n10631 =  ( n86 ) & ( n9448 )  ;
assign n10632 =  ( n86 ) & ( n9450 )  ;
assign n10633 =  ( n86 ) & ( n9452 )  ;
assign n10634 =  ( n86 ) & ( n9454 )  ;
assign n10635 =  ( n86 ) & ( n9456 )  ;
assign n10636 =  ( n87 ) & ( n9426 )  ;
assign n10637 =  ( n87 ) & ( n9428 )  ;
assign n10638 =  ( n87 ) & ( n9430 )  ;
assign n10639 =  ( n87 ) & ( n9432 )  ;
assign n10640 =  ( n87 ) & ( n9434 )  ;
assign n10641 =  ( n87 ) & ( n9436 )  ;
assign n10642 =  ( n87 ) & ( n9438 )  ;
assign n10643 =  ( n87 ) & ( n9440 )  ;
assign n10644 =  ( n87 ) & ( n9442 )  ;
assign n10645 =  ( n87 ) & ( n9444 )  ;
assign n10646 =  ( n87 ) & ( n9446 )  ;
assign n10647 =  ( n87 ) & ( n9448 )  ;
assign n10648 =  ( n87 ) & ( n9450 )  ;
assign n10649 =  ( n87 ) & ( n9452 )  ;
assign n10650 =  ( n87 ) & ( n9454 )  ;
assign n10651 =  ( n87 ) & ( n9456 )  ;
assign n10652 =  ( n88 ) & ( n9426 )  ;
assign n10653 =  ( n88 ) & ( n9428 )  ;
assign n10654 =  ( n88 ) & ( n9430 )  ;
assign n10655 =  ( n88 ) & ( n9432 )  ;
assign n10656 =  ( n88 ) & ( n9434 )  ;
assign n10657 =  ( n88 ) & ( n9436 )  ;
assign n10658 =  ( n88 ) & ( n9438 )  ;
assign n10659 =  ( n88 ) & ( n9440 )  ;
assign n10660 =  ( n88 ) & ( n9442 )  ;
assign n10661 =  ( n88 ) & ( n9444 )  ;
assign n10662 =  ( n88 ) & ( n9446 )  ;
assign n10663 =  ( n88 ) & ( n9448 )  ;
assign n10664 =  ( n88 ) & ( n9450 )  ;
assign n10665 =  ( n88 ) & ( n9452 )  ;
assign n10666 =  ( n88 ) & ( n9454 )  ;
assign n10667 =  ( n88 ) & ( n9456 )  ;
assign n10668 =  ( n89 ) & ( n9426 )  ;
assign n10669 =  ( n89 ) & ( n9428 )  ;
assign n10670 =  ( n89 ) & ( n9430 )  ;
assign n10671 =  ( n89 ) & ( n9432 )  ;
assign n10672 =  ( n89 ) & ( n9434 )  ;
assign n10673 =  ( n89 ) & ( n9436 )  ;
assign n10674 =  ( n89 ) & ( n9438 )  ;
assign n10675 =  ( n89 ) & ( n9440 )  ;
assign n10676 =  ( n89 ) & ( n9442 )  ;
assign n10677 =  ( n89 ) & ( n9444 )  ;
assign n10678 =  ( n89 ) & ( n9446 )  ;
assign n10679 =  ( n89 ) & ( n9448 )  ;
assign n10680 =  ( n89 ) & ( n9450 )  ;
assign n10681 =  ( n89 ) & ( n9452 )  ;
assign n10682 =  ( n89 ) & ( n9454 )  ;
assign n10683 =  ( n89 ) & ( n9456 )  ;
assign n10684 =  ( n90 ) & ( n9426 )  ;
assign n10685 =  ( n90 ) & ( n9428 )  ;
assign n10686 =  ( n90 ) & ( n9430 )  ;
assign n10687 =  ( n90 ) & ( n9432 )  ;
assign n10688 =  ( n90 ) & ( n9434 )  ;
assign n10689 =  ( n90 ) & ( n9436 )  ;
assign n10690 =  ( n90 ) & ( n9438 )  ;
assign n10691 =  ( n90 ) & ( n9440 )  ;
assign n10692 =  ( n90 ) & ( n9442 )  ;
assign n10693 =  ( n90 ) & ( n9444 )  ;
assign n10694 =  ( n90 ) & ( n9446 )  ;
assign n10695 =  ( n90 ) & ( n9448 )  ;
assign n10696 =  ( n90 ) & ( n9450 )  ;
assign n10697 =  ( n90 ) & ( n9452 )  ;
assign n10698 =  ( n90 ) & ( n9454 )  ;
assign n10699 =  ( n90 ) & ( n9456 )  ;
assign n10700 =  ( n91 ) & ( n9426 )  ;
assign n10701 =  ( n91 ) & ( n9428 )  ;
assign n10702 =  ( n91 ) & ( n9430 )  ;
assign n10703 =  ( n91 ) & ( n9432 )  ;
assign n10704 =  ( n91 ) & ( n9434 )  ;
assign n10705 =  ( n91 ) & ( n9436 )  ;
assign n10706 =  ( n91 ) & ( n9438 )  ;
assign n10707 =  ( n91 ) & ( n9440 )  ;
assign n10708 =  ( n91 ) & ( n9442 )  ;
assign n10709 =  ( n91 ) & ( n9444 )  ;
assign n10710 =  ( n91 ) & ( n9446 )  ;
assign n10711 =  ( n91 ) & ( n9448 )  ;
assign n10712 =  ( n91 ) & ( n9450 )  ;
assign n10713 =  ( n91 ) & ( n9452 )  ;
assign n10714 =  ( n91 ) & ( n9454 )  ;
assign n10715 =  ( n91 ) & ( n9456 )  ;
assign n10716 =  ( n92 ) & ( n9426 )  ;
assign n10717 =  ( n92 ) & ( n9428 )  ;
assign n10718 =  ( n92 ) & ( n9430 )  ;
assign n10719 =  ( n92 ) & ( n9432 )  ;
assign n10720 =  ( n92 ) & ( n9434 )  ;
assign n10721 =  ( n92 ) & ( n9436 )  ;
assign n10722 =  ( n92 ) & ( n9438 )  ;
assign n10723 =  ( n92 ) & ( n9440 )  ;
assign n10724 =  ( n92 ) & ( n9442 )  ;
assign n10725 =  ( n92 ) & ( n9444 )  ;
assign n10726 =  ( n92 ) & ( n9446 )  ;
assign n10727 =  ( n92 ) & ( n9448 )  ;
assign n10728 =  ( n92 ) & ( n9450 )  ;
assign n10729 =  ( n92 ) & ( n9452 )  ;
assign n10730 =  ( n92 ) & ( n9454 )  ;
assign n10731 =  ( n92 ) & ( n9456 )  ;
assign n10732 =  ( n93 ) & ( n9426 )  ;
assign n10733 =  ( n93 ) & ( n9428 )  ;
assign n10734 =  ( n93 ) & ( n9430 )  ;
assign n10735 =  ( n93 ) & ( n9432 )  ;
assign n10736 =  ( n93 ) & ( n9434 )  ;
assign n10737 =  ( n93 ) & ( n9436 )  ;
assign n10738 =  ( n93 ) & ( n9438 )  ;
assign n10739 =  ( n93 ) & ( n9440 )  ;
assign n10740 =  ( n93 ) & ( n9442 )  ;
assign n10741 =  ( n93 ) & ( n9444 )  ;
assign n10742 =  ( n93 ) & ( n9446 )  ;
assign n10743 =  ( n93 ) & ( n9448 )  ;
assign n10744 =  ( n93 ) & ( n9450 )  ;
assign n10745 =  ( n93 ) & ( n9452 )  ;
assign n10746 =  ( n93 ) & ( n9454 )  ;
assign n10747 =  ( n93 ) & ( n9456 )  ;
assign n10748 =  ( n94 ) & ( n9426 )  ;
assign n10749 =  ( n94 ) & ( n9428 )  ;
assign n10750 =  ( n94 ) & ( n9430 )  ;
assign n10751 =  ( n94 ) & ( n9432 )  ;
assign n10752 =  ( n94 ) & ( n9434 )  ;
assign n10753 =  ( n94 ) & ( n9436 )  ;
assign n10754 =  ( n94 ) & ( n9438 )  ;
assign n10755 =  ( n94 ) & ( n9440 )  ;
assign n10756 =  ( n94 ) & ( n9442 )  ;
assign n10757 =  ( n94 ) & ( n9444 )  ;
assign n10758 =  ( n94 ) & ( n9446 )  ;
assign n10759 =  ( n94 ) & ( n9448 )  ;
assign n10760 =  ( n94 ) & ( n9450 )  ;
assign n10761 =  ( n94 ) & ( n9452 )  ;
assign n10762 =  ( n94 ) & ( n9454 )  ;
assign n10763 =  ( n94 ) & ( n9456 )  ;
assign n10764 =  ( n95 ) & ( n9426 )  ;
assign n10765 =  ( n95 ) & ( n9428 )  ;
assign n10766 =  ( n95 ) & ( n9430 )  ;
assign n10767 =  ( n95 ) & ( n9432 )  ;
assign n10768 =  ( n95 ) & ( n9434 )  ;
assign n10769 =  ( n95 ) & ( n9436 )  ;
assign n10770 =  ( n95 ) & ( n9438 )  ;
assign n10771 =  ( n95 ) & ( n9440 )  ;
assign n10772 =  ( n95 ) & ( n9442 )  ;
assign n10773 =  ( n95 ) & ( n9444 )  ;
assign n10774 =  ( n95 ) & ( n9446 )  ;
assign n10775 =  ( n95 ) & ( n9448 )  ;
assign n10776 =  ( n95 ) & ( n9450 )  ;
assign n10777 =  ( n95 ) & ( n9452 )  ;
assign n10778 =  ( n95 ) & ( n9454 )  ;
assign n10779 =  ( n95 ) & ( n9456 )  ;
assign n10780 =  ( n96 ) & ( n9426 )  ;
assign n10781 =  ( n96 ) & ( n9428 )  ;
assign n10782 =  ( n96 ) & ( n9430 )  ;
assign n10783 =  ( n96 ) & ( n9432 )  ;
assign n10784 =  ( n96 ) & ( n9434 )  ;
assign n10785 =  ( n96 ) & ( n9436 )  ;
assign n10786 =  ( n96 ) & ( n9438 )  ;
assign n10787 =  ( n96 ) & ( n9440 )  ;
assign n10788 =  ( n96 ) & ( n9442 )  ;
assign n10789 =  ( n96 ) & ( n9444 )  ;
assign n10790 =  ( n96 ) & ( n9446 )  ;
assign n10791 =  ( n96 ) & ( n9448 )  ;
assign n10792 =  ( n96 ) & ( n9450 )  ;
assign n10793 =  ( n96 ) & ( n9452 )  ;
assign n10794 =  ( n96 ) & ( n9454 )  ;
assign n10795 =  ( n96 ) & ( n9456 )  ;
assign n10796 =  ( n97 ) & ( n9426 )  ;
assign n10797 =  ( n97 ) & ( n9428 )  ;
assign n10798 =  ( n97 ) & ( n9430 )  ;
assign n10799 =  ( n97 ) & ( n9432 )  ;
assign n10800 =  ( n97 ) & ( n9434 )  ;
assign n10801 =  ( n97 ) & ( n9436 )  ;
assign n10802 =  ( n97 ) & ( n9438 )  ;
assign n10803 =  ( n97 ) & ( n9440 )  ;
assign n10804 =  ( n97 ) & ( n9442 )  ;
assign n10805 =  ( n97 ) & ( n9444 )  ;
assign n10806 =  ( n97 ) & ( n9446 )  ;
assign n10807 =  ( n97 ) & ( n9448 )  ;
assign n10808 =  ( n97 ) & ( n9450 )  ;
assign n10809 =  ( n97 ) & ( n9452 )  ;
assign n10810 =  ( n97 ) & ( n9454 )  ;
assign n10811 =  ( n97 ) & ( n9456 )  ;
assign n10812 =  ( n98 ) & ( n9426 )  ;
assign n10813 =  ( n98 ) & ( n9428 )  ;
assign n10814 =  ( n98 ) & ( n9430 )  ;
assign n10815 =  ( n98 ) & ( n9432 )  ;
assign n10816 =  ( n98 ) & ( n9434 )  ;
assign n10817 =  ( n98 ) & ( n9436 )  ;
assign n10818 =  ( n98 ) & ( n9438 )  ;
assign n10819 =  ( n98 ) & ( n9440 )  ;
assign n10820 =  ( n98 ) & ( n9442 )  ;
assign n10821 =  ( n98 ) & ( n9444 )  ;
assign n10822 =  ( n98 ) & ( n9446 )  ;
assign n10823 =  ( n98 ) & ( n9448 )  ;
assign n10824 =  ( n98 ) & ( n9450 )  ;
assign n10825 =  ( n98 ) & ( n9452 )  ;
assign n10826 =  ( n98 ) & ( n9454 )  ;
assign n10827 =  ( n98 ) & ( n9456 )  ;
assign n10828 =  ( n99 ) & ( n9426 )  ;
assign n10829 =  ( n99 ) & ( n9428 )  ;
assign n10830 =  ( n99 ) & ( n9430 )  ;
assign n10831 =  ( n99 ) & ( n9432 )  ;
assign n10832 =  ( n99 ) & ( n9434 )  ;
assign n10833 =  ( n99 ) & ( n9436 )  ;
assign n10834 =  ( n99 ) & ( n9438 )  ;
assign n10835 =  ( n99 ) & ( n9440 )  ;
assign n10836 =  ( n99 ) & ( n9442 )  ;
assign n10837 =  ( n99 ) & ( n9444 )  ;
assign n10838 =  ( n99 ) & ( n9446 )  ;
assign n10839 =  ( n99 ) & ( n9448 )  ;
assign n10840 =  ( n99 ) & ( n9450 )  ;
assign n10841 =  ( n99 ) & ( n9452 )  ;
assign n10842 =  ( n99 ) & ( n9454 )  ;
assign n10843 =  ( n99 ) & ( n9456 )  ;
assign n10844 =  ( n100 ) & ( n9426 )  ;
assign n10845 =  ( n100 ) & ( n9428 )  ;
assign n10846 =  ( n100 ) & ( n9430 )  ;
assign n10847 =  ( n100 ) & ( n9432 )  ;
assign n10848 =  ( n100 ) & ( n9434 )  ;
assign n10849 =  ( n100 ) & ( n9436 )  ;
assign n10850 =  ( n100 ) & ( n9438 )  ;
assign n10851 =  ( n100 ) & ( n9440 )  ;
assign n10852 =  ( n100 ) & ( n9442 )  ;
assign n10853 =  ( n100 ) & ( n9444 )  ;
assign n10854 =  ( n100 ) & ( n9446 )  ;
assign n10855 =  ( n100 ) & ( n9448 )  ;
assign n10856 =  ( n100 ) & ( n9450 )  ;
assign n10857 =  ( n100 ) & ( n9452 )  ;
assign n10858 =  ( n100 ) & ( n9454 )  ;
assign n10859 =  ( n100 ) & ( n9456 )  ;
assign n10860 =  ( n101 ) & ( n9426 )  ;
assign n10861 =  ( n101 ) & ( n9428 )  ;
assign n10862 =  ( n101 ) & ( n9430 )  ;
assign n10863 =  ( n101 ) & ( n9432 )  ;
assign n10864 =  ( n101 ) & ( n9434 )  ;
assign n10865 =  ( n101 ) & ( n9436 )  ;
assign n10866 =  ( n101 ) & ( n9438 )  ;
assign n10867 =  ( n101 ) & ( n9440 )  ;
assign n10868 =  ( n101 ) & ( n9442 )  ;
assign n10869 =  ( n101 ) & ( n9444 )  ;
assign n10870 =  ( n101 ) & ( n9446 )  ;
assign n10871 =  ( n101 ) & ( n9448 )  ;
assign n10872 =  ( n101 ) & ( n9450 )  ;
assign n10873 =  ( n101 ) & ( n9452 )  ;
assign n10874 =  ( n101 ) & ( n9454 )  ;
assign n10875 =  ( n101 ) & ( n9456 )  ;
assign n10876 =  ( n102 ) & ( n9426 )  ;
assign n10877 =  ( n102 ) & ( n9428 )  ;
assign n10878 =  ( n102 ) & ( n9430 )  ;
assign n10879 =  ( n102 ) & ( n9432 )  ;
assign n10880 =  ( n102 ) & ( n9434 )  ;
assign n10881 =  ( n102 ) & ( n9436 )  ;
assign n10882 =  ( n102 ) & ( n9438 )  ;
assign n10883 =  ( n102 ) & ( n9440 )  ;
assign n10884 =  ( n102 ) & ( n9442 )  ;
assign n10885 =  ( n102 ) & ( n9444 )  ;
assign n10886 =  ( n102 ) & ( n9446 )  ;
assign n10887 =  ( n102 ) & ( n9448 )  ;
assign n10888 =  ( n102 ) & ( n9450 )  ;
assign n10889 =  ( n102 ) & ( n9452 )  ;
assign n10890 =  ( n102 ) & ( n9454 )  ;
assign n10891 =  ( n102 ) & ( n9456 )  ;
assign n10892 =  ( n103 ) & ( n9426 )  ;
assign n10893 =  ( n103 ) & ( n9428 )  ;
assign n10894 =  ( n103 ) & ( n9430 )  ;
assign n10895 =  ( n103 ) & ( n9432 )  ;
assign n10896 =  ( n103 ) & ( n9434 )  ;
assign n10897 =  ( n103 ) & ( n9436 )  ;
assign n10898 =  ( n103 ) & ( n9438 )  ;
assign n10899 =  ( n103 ) & ( n9440 )  ;
assign n10900 =  ( n103 ) & ( n9442 )  ;
assign n10901 =  ( n103 ) & ( n9444 )  ;
assign n10902 =  ( n103 ) & ( n9446 )  ;
assign n10903 =  ( n103 ) & ( n9448 )  ;
assign n10904 =  ( n103 ) & ( n9450 )  ;
assign n10905 =  ( n103 ) & ( n9452 )  ;
assign n10906 =  ( n103 ) & ( n9454 )  ;
assign n10907 =  ( n103 ) & ( n9456 )  ;
assign n10908 =  ( n104 ) & ( n9426 )  ;
assign n10909 =  ( n104 ) & ( n9428 )  ;
assign n10910 =  ( n104 ) & ( n9430 )  ;
assign n10911 =  ( n104 ) & ( n9432 )  ;
assign n10912 =  ( n104 ) & ( n9434 )  ;
assign n10913 =  ( n104 ) & ( n9436 )  ;
assign n10914 =  ( n104 ) & ( n9438 )  ;
assign n10915 =  ( n104 ) & ( n9440 )  ;
assign n10916 =  ( n104 ) & ( n9442 )  ;
assign n10917 =  ( n104 ) & ( n9444 )  ;
assign n10918 =  ( n104 ) & ( n9446 )  ;
assign n10919 =  ( n104 ) & ( n9448 )  ;
assign n10920 =  ( n104 ) & ( n9450 )  ;
assign n10921 =  ( n104 ) & ( n9452 )  ;
assign n10922 =  ( n104 ) & ( n9454 )  ;
assign n10923 =  ( n104 ) & ( n9456 )  ;
assign n10924 =  ( n105 ) & ( n9426 )  ;
assign n10925 =  ( n105 ) & ( n9428 )  ;
assign n10926 =  ( n105 ) & ( n9430 )  ;
assign n10927 =  ( n105 ) & ( n9432 )  ;
assign n10928 =  ( n105 ) & ( n9434 )  ;
assign n10929 =  ( n105 ) & ( n9436 )  ;
assign n10930 =  ( n105 ) & ( n9438 )  ;
assign n10931 =  ( n105 ) & ( n9440 )  ;
assign n10932 =  ( n105 ) & ( n9442 )  ;
assign n10933 =  ( n105 ) & ( n9444 )  ;
assign n10934 =  ( n105 ) & ( n9446 )  ;
assign n10935 =  ( n105 ) & ( n9448 )  ;
assign n10936 =  ( n105 ) & ( n9450 )  ;
assign n10937 =  ( n105 ) & ( n9452 )  ;
assign n10938 =  ( n105 ) & ( n9454 )  ;
assign n10939 =  ( n105 ) & ( n9456 )  ;
assign n10940 =  ( n106 ) & ( n9426 )  ;
assign n10941 =  ( n106 ) & ( n9428 )  ;
assign n10942 =  ( n106 ) & ( n9430 )  ;
assign n10943 =  ( n106 ) & ( n9432 )  ;
assign n10944 =  ( n106 ) & ( n9434 )  ;
assign n10945 =  ( n106 ) & ( n9436 )  ;
assign n10946 =  ( n106 ) & ( n9438 )  ;
assign n10947 =  ( n106 ) & ( n9440 )  ;
assign n10948 =  ( n106 ) & ( n9442 )  ;
assign n10949 =  ( n106 ) & ( n9444 )  ;
assign n10950 =  ( n106 ) & ( n9446 )  ;
assign n10951 =  ( n106 ) & ( n9448 )  ;
assign n10952 =  ( n106 ) & ( n9450 )  ;
assign n10953 =  ( n106 ) & ( n9452 )  ;
assign n10954 =  ( n106 ) & ( n9454 )  ;
assign n10955 =  ( n106 ) & ( n9456 )  ;
assign n10956 =  ( n107 ) & ( n9426 )  ;
assign n10957 =  ( n107 ) & ( n9428 )  ;
assign n10958 =  ( n107 ) & ( n9430 )  ;
assign n10959 =  ( n107 ) & ( n9432 )  ;
assign n10960 =  ( n107 ) & ( n9434 )  ;
assign n10961 =  ( n107 ) & ( n9436 )  ;
assign n10962 =  ( n107 ) & ( n9438 )  ;
assign n10963 =  ( n107 ) & ( n9440 )  ;
assign n10964 =  ( n107 ) & ( n9442 )  ;
assign n10965 =  ( n107 ) & ( n9444 )  ;
assign n10966 =  ( n107 ) & ( n9446 )  ;
assign n10967 =  ( n107 ) & ( n9448 )  ;
assign n10968 =  ( n107 ) & ( n9450 )  ;
assign n10969 =  ( n107 ) & ( n9452 )  ;
assign n10970 =  ( n107 ) & ( n9454 )  ;
assign n10971 =  ( n107 ) & ( n9456 )  ;
assign n10972 =  ( n108 ) & ( n9426 )  ;
assign n10973 =  ( n108 ) & ( n9428 )  ;
assign n10974 =  ( n108 ) & ( n9430 )  ;
assign n10975 =  ( n108 ) & ( n9432 )  ;
assign n10976 =  ( n108 ) & ( n9434 )  ;
assign n10977 =  ( n108 ) & ( n9436 )  ;
assign n10978 =  ( n108 ) & ( n9438 )  ;
assign n10979 =  ( n108 ) & ( n9440 )  ;
assign n10980 =  ( n108 ) & ( n9442 )  ;
assign n10981 =  ( n108 ) & ( n9444 )  ;
assign n10982 =  ( n108 ) & ( n9446 )  ;
assign n10983 =  ( n108 ) & ( n9448 )  ;
assign n10984 =  ( n108 ) & ( n9450 )  ;
assign n10985 =  ( n108 ) & ( n9452 )  ;
assign n10986 =  ( n108 ) & ( n9454 )  ;
assign n10987 =  ( n108 ) & ( n9456 )  ;
assign n10988 =  ( n10987 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n10989 =  ( n10986 ) ? ( VREG_0_1 ) : ( n10988 ) ;
assign n10990 =  ( n10985 ) ? ( VREG_0_2 ) : ( n10989 ) ;
assign n10991 =  ( n10984 ) ? ( VREG_0_3 ) : ( n10990 ) ;
assign n10992 =  ( n10983 ) ? ( VREG_0_4 ) : ( n10991 ) ;
assign n10993 =  ( n10982 ) ? ( VREG_0_5 ) : ( n10992 ) ;
assign n10994 =  ( n10981 ) ? ( VREG_0_6 ) : ( n10993 ) ;
assign n10995 =  ( n10980 ) ? ( VREG_0_7 ) : ( n10994 ) ;
assign n10996 =  ( n10979 ) ? ( VREG_0_8 ) : ( n10995 ) ;
assign n10997 =  ( n10978 ) ? ( VREG_0_9 ) : ( n10996 ) ;
assign n10998 =  ( n10977 ) ? ( VREG_0_10 ) : ( n10997 ) ;
assign n10999 =  ( n10976 ) ? ( VREG_0_11 ) : ( n10998 ) ;
assign n11000 =  ( n10975 ) ? ( VREG_0_12 ) : ( n10999 ) ;
assign n11001 =  ( n10974 ) ? ( VREG_0_13 ) : ( n11000 ) ;
assign n11002 =  ( n10973 ) ? ( VREG_0_14 ) : ( n11001 ) ;
assign n11003 =  ( n10972 ) ? ( VREG_0_15 ) : ( n11002 ) ;
assign n11004 =  ( n10971 ) ? ( VREG_1_0 ) : ( n11003 ) ;
assign n11005 =  ( n10970 ) ? ( VREG_1_1 ) : ( n11004 ) ;
assign n11006 =  ( n10969 ) ? ( VREG_1_2 ) : ( n11005 ) ;
assign n11007 =  ( n10968 ) ? ( VREG_1_3 ) : ( n11006 ) ;
assign n11008 =  ( n10967 ) ? ( VREG_1_4 ) : ( n11007 ) ;
assign n11009 =  ( n10966 ) ? ( VREG_1_5 ) : ( n11008 ) ;
assign n11010 =  ( n10965 ) ? ( VREG_1_6 ) : ( n11009 ) ;
assign n11011 =  ( n10964 ) ? ( VREG_1_7 ) : ( n11010 ) ;
assign n11012 =  ( n10963 ) ? ( VREG_1_8 ) : ( n11011 ) ;
assign n11013 =  ( n10962 ) ? ( VREG_1_9 ) : ( n11012 ) ;
assign n11014 =  ( n10961 ) ? ( VREG_1_10 ) : ( n11013 ) ;
assign n11015 =  ( n10960 ) ? ( VREG_1_11 ) : ( n11014 ) ;
assign n11016 =  ( n10959 ) ? ( VREG_1_12 ) : ( n11015 ) ;
assign n11017 =  ( n10958 ) ? ( VREG_1_13 ) : ( n11016 ) ;
assign n11018 =  ( n10957 ) ? ( VREG_1_14 ) : ( n11017 ) ;
assign n11019 =  ( n10956 ) ? ( VREG_1_15 ) : ( n11018 ) ;
assign n11020 =  ( n10955 ) ? ( VREG_2_0 ) : ( n11019 ) ;
assign n11021 =  ( n10954 ) ? ( VREG_2_1 ) : ( n11020 ) ;
assign n11022 =  ( n10953 ) ? ( VREG_2_2 ) : ( n11021 ) ;
assign n11023 =  ( n10952 ) ? ( VREG_2_3 ) : ( n11022 ) ;
assign n11024 =  ( n10951 ) ? ( VREG_2_4 ) : ( n11023 ) ;
assign n11025 =  ( n10950 ) ? ( VREG_2_5 ) : ( n11024 ) ;
assign n11026 =  ( n10949 ) ? ( VREG_2_6 ) : ( n11025 ) ;
assign n11027 =  ( n10948 ) ? ( VREG_2_7 ) : ( n11026 ) ;
assign n11028 =  ( n10947 ) ? ( VREG_2_8 ) : ( n11027 ) ;
assign n11029 =  ( n10946 ) ? ( VREG_2_9 ) : ( n11028 ) ;
assign n11030 =  ( n10945 ) ? ( VREG_2_10 ) : ( n11029 ) ;
assign n11031 =  ( n10944 ) ? ( VREG_2_11 ) : ( n11030 ) ;
assign n11032 =  ( n10943 ) ? ( VREG_2_12 ) : ( n11031 ) ;
assign n11033 =  ( n10942 ) ? ( VREG_2_13 ) : ( n11032 ) ;
assign n11034 =  ( n10941 ) ? ( VREG_2_14 ) : ( n11033 ) ;
assign n11035 =  ( n10940 ) ? ( VREG_2_15 ) : ( n11034 ) ;
assign n11036 =  ( n10939 ) ? ( VREG_3_0 ) : ( n11035 ) ;
assign n11037 =  ( n10938 ) ? ( VREG_3_1 ) : ( n11036 ) ;
assign n11038 =  ( n10937 ) ? ( VREG_3_2 ) : ( n11037 ) ;
assign n11039 =  ( n10936 ) ? ( VREG_3_3 ) : ( n11038 ) ;
assign n11040 =  ( n10935 ) ? ( VREG_3_4 ) : ( n11039 ) ;
assign n11041 =  ( n10934 ) ? ( VREG_3_5 ) : ( n11040 ) ;
assign n11042 =  ( n10933 ) ? ( VREG_3_6 ) : ( n11041 ) ;
assign n11043 =  ( n10932 ) ? ( VREG_3_7 ) : ( n11042 ) ;
assign n11044 =  ( n10931 ) ? ( VREG_3_8 ) : ( n11043 ) ;
assign n11045 =  ( n10930 ) ? ( VREG_3_9 ) : ( n11044 ) ;
assign n11046 =  ( n10929 ) ? ( VREG_3_10 ) : ( n11045 ) ;
assign n11047 =  ( n10928 ) ? ( VREG_3_11 ) : ( n11046 ) ;
assign n11048 =  ( n10927 ) ? ( VREG_3_12 ) : ( n11047 ) ;
assign n11049 =  ( n10926 ) ? ( VREG_3_13 ) : ( n11048 ) ;
assign n11050 =  ( n10925 ) ? ( VREG_3_14 ) : ( n11049 ) ;
assign n11051 =  ( n10924 ) ? ( VREG_3_15 ) : ( n11050 ) ;
assign n11052 =  ( n10923 ) ? ( VREG_4_0 ) : ( n11051 ) ;
assign n11053 =  ( n10922 ) ? ( VREG_4_1 ) : ( n11052 ) ;
assign n11054 =  ( n10921 ) ? ( VREG_4_2 ) : ( n11053 ) ;
assign n11055 =  ( n10920 ) ? ( VREG_4_3 ) : ( n11054 ) ;
assign n11056 =  ( n10919 ) ? ( VREG_4_4 ) : ( n11055 ) ;
assign n11057 =  ( n10918 ) ? ( VREG_4_5 ) : ( n11056 ) ;
assign n11058 =  ( n10917 ) ? ( VREG_4_6 ) : ( n11057 ) ;
assign n11059 =  ( n10916 ) ? ( VREG_4_7 ) : ( n11058 ) ;
assign n11060 =  ( n10915 ) ? ( VREG_4_8 ) : ( n11059 ) ;
assign n11061 =  ( n10914 ) ? ( VREG_4_9 ) : ( n11060 ) ;
assign n11062 =  ( n10913 ) ? ( VREG_4_10 ) : ( n11061 ) ;
assign n11063 =  ( n10912 ) ? ( VREG_4_11 ) : ( n11062 ) ;
assign n11064 =  ( n10911 ) ? ( VREG_4_12 ) : ( n11063 ) ;
assign n11065 =  ( n10910 ) ? ( VREG_4_13 ) : ( n11064 ) ;
assign n11066 =  ( n10909 ) ? ( VREG_4_14 ) : ( n11065 ) ;
assign n11067 =  ( n10908 ) ? ( VREG_4_15 ) : ( n11066 ) ;
assign n11068 =  ( n10907 ) ? ( VREG_5_0 ) : ( n11067 ) ;
assign n11069 =  ( n10906 ) ? ( VREG_5_1 ) : ( n11068 ) ;
assign n11070 =  ( n10905 ) ? ( VREG_5_2 ) : ( n11069 ) ;
assign n11071 =  ( n10904 ) ? ( VREG_5_3 ) : ( n11070 ) ;
assign n11072 =  ( n10903 ) ? ( VREG_5_4 ) : ( n11071 ) ;
assign n11073 =  ( n10902 ) ? ( VREG_5_5 ) : ( n11072 ) ;
assign n11074 =  ( n10901 ) ? ( VREG_5_6 ) : ( n11073 ) ;
assign n11075 =  ( n10900 ) ? ( VREG_5_7 ) : ( n11074 ) ;
assign n11076 =  ( n10899 ) ? ( VREG_5_8 ) : ( n11075 ) ;
assign n11077 =  ( n10898 ) ? ( VREG_5_9 ) : ( n11076 ) ;
assign n11078 =  ( n10897 ) ? ( VREG_5_10 ) : ( n11077 ) ;
assign n11079 =  ( n10896 ) ? ( VREG_5_11 ) : ( n11078 ) ;
assign n11080 =  ( n10895 ) ? ( VREG_5_12 ) : ( n11079 ) ;
assign n11081 =  ( n10894 ) ? ( VREG_5_13 ) : ( n11080 ) ;
assign n11082 =  ( n10893 ) ? ( VREG_5_14 ) : ( n11081 ) ;
assign n11083 =  ( n10892 ) ? ( VREG_5_15 ) : ( n11082 ) ;
assign n11084 =  ( n10891 ) ? ( VREG_6_0 ) : ( n11083 ) ;
assign n11085 =  ( n10890 ) ? ( VREG_6_1 ) : ( n11084 ) ;
assign n11086 =  ( n10889 ) ? ( VREG_6_2 ) : ( n11085 ) ;
assign n11087 =  ( n10888 ) ? ( VREG_6_3 ) : ( n11086 ) ;
assign n11088 =  ( n10887 ) ? ( VREG_6_4 ) : ( n11087 ) ;
assign n11089 =  ( n10886 ) ? ( VREG_6_5 ) : ( n11088 ) ;
assign n11090 =  ( n10885 ) ? ( VREG_6_6 ) : ( n11089 ) ;
assign n11091 =  ( n10884 ) ? ( VREG_6_7 ) : ( n11090 ) ;
assign n11092 =  ( n10883 ) ? ( VREG_6_8 ) : ( n11091 ) ;
assign n11093 =  ( n10882 ) ? ( VREG_6_9 ) : ( n11092 ) ;
assign n11094 =  ( n10881 ) ? ( VREG_6_10 ) : ( n11093 ) ;
assign n11095 =  ( n10880 ) ? ( VREG_6_11 ) : ( n11094 ) ;
assign n11096 =  ( n10879 ) ? ( VREG_6_12 ) : ( n11095 ) ;
assign n11097 =  ( n10878 ) ? ( VREG_6_13 ) : ( n11096 ) ;
assign n11098 =  ( n10877 ) ? ( VREG_6_14 ) : ( n11097 ) ;
assign n11099 =  ( n10876 ) ? ( VREG_6_15 ) : ( n11098 ) ;
assign n11100 =  ( n10875 ) ? ( VREG_7_0 ) : ( n11099 ) ;
assign n11101 =  ( n10874 ) ? ( VREG_7_1 ) : ( n11100 ) ;
assign n11102 =  ( n10873 ) ? ( VREG_7_2 ) : ( n11101 ) ;
assign n11103 =  ( n10872 ) ? ( VREG_7_3 ) : ( n11102 ) ;
assign n11104 =  ( n10871 ) ? ( VREG_7_4 ) : ( n11103 ) ;
assign n11105 =  ( n10870 ) ? ( VREG_7_5 ) : ( n11104 ) ;
assign n11106 =  ( n10869 ) ? ( VREG_7_6 ) : ( n11105 ) ;
assign n11107 =  ( n10868 ) ? ( VREG_7_7 ) : ( n11106 ) ;
assign n11108 =  ( n10867 ) ? ( VREG_7_8 ) : ( n11107 ) ;
assign n11109 =  ( n10866 ) ? ( VREG_7_9 ) : ( n11108 ) ;
assign n11110 =  ( n10865 ) ? ( VREG_7_10 ) : ( n11109 ) ;
assign n11111 =  ( n10864 ) ? ( VREG_7_11 ) : ( n11110 ) ;
assign n11112 =  ( n10863 ) ? ( VREG_7_12 ) : ( n11111 ) ;
assign n11113 =  ( n10862 ) ? ( VREG_7_13 ) : ( n11112 ) ;
assign n11114 =  ( n10861 ) ? ( VREG_7_14 ) : ( n11113 ) ;
assign n11115 =  ( n10860 ) ? ( VREG_7_15 ) : ( n11114 ) ;
assign n11116 =  ( n10859 ) ? ( VREG_8_0 ) : ( n11115 ) ;
assign n11117 =  ( n10858 ) ? ( VREG_8_1 ) : ( n11116 ) ;
assign n11118 =  ( n10857 ) ? ( VREG_8_2 ) : ( n11117 ) ;
assign n11119 =  ( n10856 ) ? ( VREG_8_3 ) : ( n11118 ) ;
assign n11120 =  ( n10855 ) ? ( VREG_8_4 ) : ( n11119 ) ;
assign n11121 =  ( n10854 ) ? ( VREG_8_5 ) : ( n11120 ) ;
assign n11122 =  ( n10853 ) ? ( VREG_8_6 ) : ( n11121 ) ;
assign n11123 =  ( n10852 ) ? ( VREG_8_7 ) : ( n11122 ) ;
assign n11124 =  ( n10851 ) ? ( VREG_8_8 ) : ( n11123 ) ;
assign n11125 =  ( n10850 ) ? ( VREG_8_9 ) : ( n11124 ) ;
assign n11126 =  ( n10849 ) ? ( VREG_8_10 ) : ( n11125 ) ;
assign n11127 =  ( n10848 ) ? ( VREG_8_11 ) : ( n11126 ) ;
assign n11128 =  ( n10847 ) ? ( VREG_8_12 ) : ( n11127 ) ;
assign n11129 =  ( n10846 ) ? ( VREG_8_13 ) : ( n11128 ) ;
assign n11130 =  ( n10845 ) ? ( VREG_8_14 ) : ( n11129 ) ;
assign n11131 =  ( n10844 ) ? ( VREG_8_15 ) : ( n11130 ) ;
assign n11132 =  ( n10843 ) ? ( VREG_9_0 ) : ( n11131 ) ;
assign n11133 =  ( n10842 ) ? ( VREG_9_1 ) : ( n11132 ) ;
assign n11134 =  ( n10841 ) ? ( VREG_9_2 ) : ( n11133 ) ;
assign n11135 =  ( n10840 ) ? ( VREG_9_3 ) : ( n11134 ) ;
assign n11136 =  ( n10839 ) ? ( VREG_9_4 ) : ( n11135 ) ;
assign n11137 =  ( n10838 ) ? ( VREG_9_5 ) : ( n11136 ) ;
assign n11138 =  ( n10837 ) ? ( VREG_9_6 ) : ( n11137 ) ;
assign n11139 =  ( n10836 ) ? ( VREG_9_7 ) : ( n11138 ) ;
assign n11140 =  ( n10835 ) ? ( VREG_9_8 ) : ( n11139 ) ;
assign n11141 =  ( n10834 ) ? ( VREG_9_9 ) : ( n11140 ) ;
assign n11142 =  ( n10833 ) ? ( VREG_9_10 ) : ( n11141 ) ;
assign n11143 =  ( n10832 ) ? ( VREG_9_11 ) : ( n11142 ) ;
assign n11144 =  ( n10831 ) ? ( VREG_9_12 ) : ( n11143 ) ;
assign n11145 =  ( n10830 ) ? ( VREG_9_13 ) : ( n11144 ) ;
assign n11146 =  ( n10829 ) ? ( VREG_9_14 ) : ( n11145 ) ;
assign n11147 =  ( n10828 ) ? ( VREG_9_15 ) : ( n11146 ) ;
assign n11148 =  ( n10827 ) ? ( VREG_10_0 ) : ( n11147 ) ;
assign n11149 =  ( n10826 ) ? ( VREG_10_1 ) : ( n11148 ) ;
assign n11150 =  ( n10825 ) ? ( VREG_10_2 ) : ( n11149 ) ;
assign n11151 =  ( n10824 ) ? ( VREG_10_3 ) : ( n11150 ) ;
assign n11152 =  ( n10823 ) ? ( VREG_10_4 ) : ( n11151 ) ;
assign n11153 =  ( n10822 ) ? ( VREG_10_5 ) : ( n11152 ) ;
assign n11154 =  ( n10821 ) ? ( VREG_10_6 ) : ( n11153 ) ;
assign n11155 =  ( n10820 ) ? ( VREG_10_7 ) : ( n11154 ) ;
assign n11156 =  ( n10819 ) ? ( VREG_10_8 ) : ( n11155 ) ;
assign n11157 =  ( n10818 ) ? ( VREG_10_9 ) : ( n11156 ) ;
assign n11158 =  ( n10817 ) ? ( VREG_10_10 ) : ( n11157 ) ;
assign n11159 =  ( n10816 ) ? ( VREG_10_11 ) : ( n11158 ) ;
assign n11160 =  ( n10815 ) ? ( VREG_10_12 ) : ( n11159 ) ;
assign n11161 =  ( n10814 ) ? ( VREG_10_13 ) : ( n11160 ) ;
assign n11162 =  ( n10813 ) ? ( VREG_10_14 ) : ( n11161 ) ;
assign n11163 =  ( n10812 ) ? ( VREG_10_15 ) : ( n11162 ) ;
assign n11164 =  ( n10811 ) ? ( VREG_11_0 ) : ( n11163 ) ;
assign n11165 =  ( n10810 ) ? ( VREG_11_1 ) : ( n11164 ) ;
assign n11166 =  ( n10809 ) ? ( VREG_11_2 ) : ( n11165 ) ;
assign n11167 =  ( n10808 ) ? ( VREG_11_3 ) : ( n11166 ) ;
assign n11168 =  ( n10807 ) ? ( VREG_11_4 ) : ( n11167 ) ;
assign n11169 =  ( n10806 ) ? ( VREG_11_5 ) : ( n11168 ) ;
assign n11170 =  ( n10805 ) ? ( VREG_11_6 ) : ( n11169 ) ;
assign n11171 =  ( n10804 ) ? ( VREG_11_7 ) : ( n11170 ) ;
assign n11172 =  ( n10803 ) ? ( VREG_11_8 ) : ( n11171 ) ;
assign n11173 =  ( n10802 ) ? ( VREG_11_9 ) : ( n11172 ) ;
assign n11174 =  ( n10801 ) ? ( VREG_11_10 ) : ( n11173 ) ;
assign n11175 =  ( n10800 ) ? ( VREG_11_11 ) : ( n11174 ) ;
assign n11176 =  ( n10799 ) ? ( VREG_11_12 ) : ( n11175 ) ;
assign n11177 =  ( n10798 ) ? ( VREG_11_13 ) : ( n11176 ) ;
assign n11178 =  ( n10797 ) ? ( VREG_11_14 ) : ( n11177 ) ;
assign n11179 =  ( n10796 ) ? ( VREG_11_15 ) : ( n11178 ) ;
assign n11180 =  ( n10795 ) ? ( VREG_12_0 ) : ( n11179 ) ;
assign n11181 =  ( n10794 ) ? ( VREG_12_1 ) : ( n11180 ) ;
assign n11182 =  ( n10793 ) ? ( VREG_12_2 ) : ( n11181 ) ;
assign n11183 =  ( n10792 ) ? ( VREG_12_3 ) : ( n11182 ) ;
assign n11184 =  ( n10791 ) ? ( VREG_12_4 ) : ( n11183 ) ;
assign n11185 =  ( n10790 ) ? ( VREG_12_5 ) : ( n11184 ) ;
assign n11186 =  ( n10789 ) ? ( VREG_12_6 ) : ( n11185 ) ;
assign n11187 =  ( n10788 ) ? ( VREG_12_7 ) : ( n11186 ) ;
assign n11188 =  ( n10787 ) ? ( VREG_12_8 ) : ( n11187 ) ;
assign n11189 =  ( n10786 ) ? ( VREG_12_9 ) : ( n11188 ) ;
assign n11190 =  ( n10785 ) ? ( VREG_12_10 ) : ( n11189 ) ;
assign n11191 =  ( n10784 ) ? ( VREG_12_11 ) : ( n11190 ) ;
assign n11192 =  ( n10783 ) ? ( VREG_12_12 ) : ( n11191 ) ;
assign n11193 =  ( n10782 ) ? ( VREG_12_13 ) : ( n11192 ) ;
assign n11194 =  ( n10781 ) ? ( VREG_12_14 ) : ( n11193 ) ;
assign n11195 =  ( n10780 ) ? ( VREG_12_15 ) : ( n11194 ) ;
assign n11196 =  ( n10779 ) ? ( VREG_13_0 ) : ( n11195 ) ;
assign n11197 =  ( n10778 ) ? ( VREG_13_1 ) : ( n11196 ) ;
assign n11198 =  ( n10777 ) ? ( VREG_13_2 ) : ( n11197 ) ;
assign n11199 =  ( n10776 ) ? ( VREG_13_3 ) : ( n11198 ) ;
assign n11200 =  ( n10775 ) ? ( VREG_13_4 ) : ( n11199 ) ;
assign n11201 =  ( n10774 ) ? ( VREG_13_5 ) : ( n11200 ) ;
assign n11202 =  ( n10773 ) ? ( VREG_13_6 ) : ( n11201 ) ;
assign n11203 =  ( n10772 ) ? ( VREG_13_7 ) : ( n11202 ) ;
assign n11204 =  ( n10771 ) ? ( VREG_13_8 ) : ( n11203 ) ;
assign n11205 =  ( n10770 ) ? ( VREG_13_9 ) : ( n11204 ) ;
assign n11206 =  ( n10769 ) ? ( VREG_13_10 ) : ( n11205 ) ;
assign n11207 =  ( n10768 ) ? ( VREG_13_11 ) : ( n11206 ) ;
assign n11208 =  ( n10767 ) ? ( VREG_13_12 ) : ( n11207 ) ;
assign n11209 =  ( n10766 ) ? ( VREG_13_13 ) : ( n11208 ) ;
assign n11210 =  ( n10765 ) ? ( VREG_13_14 ) : ( n11209 ) ;
assign n11211 =  ( n10764 ) ? ( VREG_13_15 ) : ( n11210 ) ;
assign n11212 =  ( n10763 ) ? ( VREG_14_0 ) : ( n11211 ) ;
assign n11213 =  ( n10762 ) ? ( VREG_14_1 ) : ( n11212 ) ;
assign n11214 =  ( n10761 ) ? ( VREG_14_2 ) : ( n11213 ) ;
assign n11215 =  ( n10760 ) ? ( VREG_14_3 ) : ( n11214 ) ;
assign n11216 =  ( n10759 ) ? ( VREG_14_4 ) : ( n11215 ) ;
assign n11217 =  ( n10758 ) ? ( VREG_14_5 ) : ( n11216 ) ;
assign n11218 =  ( n10757 ) ? ( VREG_14_6 ) : ( n11217 ) ;
assign n11219 =  ( n10756 ) ? ( VREG_14_7 ) : ( n11218 ) ;
assign n11220 =  ( n10755 ) ? ( VREG_14_8 ) : ( n11219 ) ;
assign n11221 =  ( n10754 ) ? ( VREG_14_9 ) : ( n11220 ) ;
assign n11222 =  ( n10753 ) ? ( VREG_14_10 ) : ( n11221 ) ;
assign n11223 =  ( n10752 ) ? ( VREG_14_11 ) : ( n11222 ) ;
assign n11224 =  ( n10751 ) ? ( VREG_14_12 ) : ( n11223 ) ;
assign n11225 =  ( n10750 ) ? ( VREG_14_13 ) : ( n11224 ) ;
assign n11226 =  ( n10749 ) ? ( VREG_14_14 ) : ( n11225 ) ;
assign n11227 =  ( n10748 ) ? ( VREG_14_15 ) : ( n11226 ) ;
assign n11228 =  ( n10747 ) ? ( VREG_15_0 ) : ( n11227 ) ;
assign n11229 =  ( n10746 ) ? ( VREG_15_1 ) : ( n11228 ) ;
assign n11230 =  ( n10745 ) ? ( VREG_15_2 ) : ( n11229 ) ;
assign n11231 =  ( n10744 ) ? ( VREG_15_3 ) : ( n11230 ) ;
assign n11232 =  ( n10743 ) ? ( VREG_15_4 ) : ( n11231 ) ;
assign n11233 =  ( n10742 ) ? ( VREG_15_5 ) : ( n11232 ) ;
assign n11234 =  ( n10741 ) ? ( VREG_15_6 ) : ( n11233 ) ;
assign n11235 =  ( n10740 ) ? ( VREG_15_7 ) : ( n11234 ) ;
assign n11236 =  ( n10739 ) ? ( VREG_15_8 ) : ( n11235 ) ;
assign n11237 =  ( n10738 ) ? ( VREG_15_9 ) : ( n11236 ) ;
assign n11238 =  ( n10737 ) ? ( VREG_15_10 ) : ( n11237 ) ;
assign n11239 =  ( n10736 ) ? ( VREG_15_11 ) : ( n11238 ) ;
assign n11240 =  ( n10735 ) ? ( VREG_15_12 ) : ( n11239 ) ;
assign n11241 =  ( n10734 ) ? ( VREG_15_13 ) : ( n11240 ) ;
assign n11242 =  ( n10733 ) ? ( VREG_15_14 ) : ( n11241 ) ;
assign n11243 =  ( n10732 ) ? ( VREG_15_15 ) : ( n11242 ) ;
assign n11244 =  ( n10731 ) ? ( VREG_16_0 ) : ( n11243 ) ;
assign n11245 =  ( n10730 ) ? ( VREG_16_1 ) : ( n11244 ) ;
assign n11246 =  ( n10729 ) ? ( VREG_16_2 ) : ( n11245 ) ;
assign n11247 =  ( n10728 ) ? ( VREG_16_3 ) : ( n11246 ) ;
assign n11248 =  ( n10727 ) ? ( VREG_16_4 ) : ( n11247 ) ;
assign n11249 =  ( n10726 ) ? ( VREG_16_5 ) : ( n11248 ) ;
assign n11250 =  ( n10725 ) ? ( VREG_16_6 ) : ( n11249 ) ;
assign n11251 =  ( n10724 ) ? ( VREG_16_7 ) : ( n11250 ) ;
assign n11252 =  ( n10723 ) ? ( VREG_16_8 ) : ( n11251 ) ;
assign n11253 =  ( n10722 ) ? ( VREG_16_9 ) : ( n11252 ) ;
assign n11254 =  ( n10721 ) ? ( VREG_16_10 ) : ( n11253 ) ;
assign n11255 =  ( n10720 ) ? ( VREG_16_11 ) : ( n11254 ) ;
assign n11256 =  ( n10719 ) ? ( VREG_16_12 ) : ( n11255 ) ;
assign n11257 =  ( n10718 ) ? ( VREG_16_13 ) : ( n11256 ) ;
assign n11258 =  ( n10717 ) ? ( VREG_16_14 ) : ( n11257 ) ;
assign n11259 =  ( n10716 ) ? ( VREG_16_15 ) : ( n11258 ) ;
assign n11260 =  ( n10715 ) ? ( VREG_17_0 ) : ( n11259 ) ;
assign n11261 =  ( n10714 ) ? ( VREG_17_1 ) : ( n11260 ) ;
assign n11262 =  ( n10713 ) ? ( VREG_17_2 ) : ( n11261 ) ;
assign n11263 =  ( n10712 ) ? ( VREG_17_3 ) : ( n11262 ) ;
assign n11264 =  ( n10711 ) ? ( VREG_17_4 ) : ( n11263 ) ;
assign n11265 =  ( n10710 ) ? ( VREG_17_5 ) : ( n11264 ) ;
assign n11266 =  ( n10709 ) ? ( VREG_17_6 ) : ( n11265 ) ;
assign n11267 =  ( n10708 ) ? ( VREG_17_7 ) : ( n11266 ) ;
assign n11268 =  ( n10707 ) ? ( VREG_17_8 ) : ( n11267 ) ;
assign n11269 =  ( n10706 ) ? ( VREG_17_9 ) : ( n11268 ) ;
assign n11270 =  ( n10705 ) ? ( VREG_17_10 ) : ( n11269 ) ;
assign n11271 =  ( n10704 ) ? ( VREG_17_11 ) : ( n11270 ) ;
assign n11272 =  ( n10703 ) ? ( VREG_17_12 ) : ( n11271 ) ;
assign n11273 =  ( n10702 ) ? ( VREG_17_13 ) : ( n11272 ) ;
assign n11274 =  ( n10701 ) ? ( VREG_17_14 ) : ( n11273 ) ;
assign n11275 =  ( n10700 ) ? ( VREG_17_15 ) : ( n11274 ) ;
assign n11276 =  ( n10699 ) ? ( VREG_18_0 ) : ( n11275 ) ;
assign n11277 =  ( n10698 ) ? ( VREG_18_1 ) : ( n11276 ) ;
assign n11278 =  ( n10697 ) ? ( VREG_18_2 ) : ( n11277 ) ;
assign n11279 =  ( n10696 ) ? ( VREG_18_3 ) : ( n11278 ) ;
assign n11280 =  ( n10695 ) ? ( VREG_18_4 ) : ( n11279 ) ;
assign n11281 =  ( n10694 ) ? ( VREG_18_5 ) : ( n11280 ) ;
assign n11282 =  ( n10693 ) ? ( VREG_18_6 ) : ( n11281 ) ;
assign n11283 =  ( n10692 ) ? ( VREG_18_7 ) : ( n11282 ) ;
assign n11284 =  ( n10691 ) ? ( VREG_18_8 ) : ( n11283 ) ;
assign n11285 =  ( n10690 ) ? ( VREG_18_9 ) : ( n11284 ) ;
assign n11286 =  ( n10689 ) ? ( VREG_18_10 ) : ( n11285 ) ;
assign n11287 =  ( n10688 ) ? ( VREG_18_11 ) : ( n11286 ) ;
assign n11288 =  ( n10687 ) ? ( VREG_18_12 ) : ( n11287 ) ;
assign n11289 =  ( n10686 ) ? ( VREG_18_13 ) : ( n11288 ) ;
assign n11290 =  ( n10685 ) ? ( VREG_18_14 ) : ( n11289 ) ;
assign n11291 =  ( n10684 ) ? ( VREG_18_15 ) : ( n11290 ) ;
assign n11292 =  ( n10683 ) ? ( VREG_19_0 ) : ( n11291 ) ;
assign n11293 =  ( n10682 ) ? ( VREG_19_1 ) : ( n11292 ) ;
assign n11294 =  ( n10681 ) ? ( VREG_19_2 ) : ( n11293 ) ;
assign n11295 =  ( n10680 ) ? ( VREG_19_3 ) : ( n11294 ) ;
assign n11296 =  ( n10679 ) ? ( VREG_19_4 ) : ( n11295 ) ;
assign n11297 =  ( n10678 ) ? ( VREG_19_5 ) : ( n11296 ) ;
assign n11298 =  ( n10677 ) ? ( VREG_19_6 ) : ( n11297 ) ;
assign n11299 =  ( n10676 ) ? ( VREG_19_7 ) : ( n11298 ) ;
assign n11300 =  ( n10675 ) ? ( VREG_19_8 ) : ( n11299 ) ;
assign n11301 =  ( n10674 ) ? ( VREG_19_9 ) : ( n11300 ) ;
assign n11302 =  ( n10673 ) ? ( VREG_19_10 ) : ( n11301 ) ;
assign n11303 =  ( n10672 ) ? ( VREG_19_11 ) : ( n11302 ) ;
assign n11304 =  ( n10671 ) ? ( VREG_19_12 ) : ( n11303 ) ;
assign n11305 =  ( n10670 ) ? ( VREG_19_13 ) : ( n11304 ) ;
assign n11306 =  ( n10669 ) ? ( VREG_19_14 ) : ( n11305 ) ;
assign n11307 =  ( n10668 ) ? ( VREG_19_15 ) : ( n11306 ) ;
assign n11308 =  ( n10667 ) ? ( VREG_20_0 ) : ( n11307 ) ;
assign n11309 =  ( n10666 ) ? ( VREG_20_1 ) : ( n11308 ) ;
assign n11310 =  ( n10665 ) ? ( VREG_20_2 ) : ( n11309 ) ;
assign n11311 =  ( n10664 ) ? ( VREG_20_3 ) : ( n11310 ) ;
assign n11312 =  ( n10663 ) ? ( VREG_20_4 ) : ( n11311 ) ;
assign n11313 =  ( n10662 ) ? ( VREG_20_5 ) : ( n11312 ) ;
assign n11314 =  ( n10661 ) ? ( VREG_20_6 ) : ( n11313 ) ;
assign n11315 =  ( n10660 ) ? ( VREG_20_7 ) : ( n11314 ) ;
assign n11316 =  ( n10659 ) ? ( VREG_20_8 ) : ( n11315 ) ;
assign n11317 =  ( n10658 ) ? ( VREG_20_9 ) : ( n11316 ) ;
assign n11318 =  ( n10657 ) ? ( VREG_20_10 ) : ( n11317 ) ;
assign n11319 =  ( n10656 ) ? ( VREG_20_11 ) : ( n11318 ) ;
assign n11320 =  ( n10655 ) ? ( VREG_20_12 ) : ( n11319 ) ;
assign n11321 =  ( n10654 ) ? ( VREG_20_13 ) : ( n11320 ) ;
assign n11322 =  ( n10653 ) ? ( VREG_20_14 ) : ( n11321 ) ;
assign n11323 =  ( n10652 ) ? ( VREG_20_15 ) : ( n11322 ) ;
assign n11324 =  ( n10651 ) ? ( VREG_21_0 ) : ( n11323 ) ;
assign n11325 =  ( n10650 ) ? ( VREG_21_1 ) : ( n11324 ) ;
assign n11326 =  ( n10649 ) ? ( VREG_21_2 ) : ( n11325 ) ;
assign n11327 =  ( n10648 ) ? ( VREG_21_3 ) : ( n11326 ) ;
assign n11328 =  ( n10647 ) ? ( VREG_21_4 ) : ( n11327 ) ;
assign n11329 =  ( n10646 ) ? ( VREG_21_5 ) : ( n11328 ) ;
assign n11330 =  ( n10645 ) ? ( VREG_21_6 ) : ( n11329 ) ;
assign n11331 =  ( n10644 ) ? ( VREG_21_7 ) : ( n11330 ) ;
assign n11332 =  ( n10643 ) ? ( VREG_21_8 ) : ( n11331 ) ;
assign n11333 =  ( n10642 ) ? ( VREG_21_9 ) : ( n11332 ) ;
assign n11334 =  ( n10641 ) ? ( VREG_21_10 ) : ( n11333 ) ;
assign n11335 =  ( n10640 ) ? ( VREG_21_11 ) : ( n11334 ) ;
assign n11336 =  ( n10639 ) ? ( VREG_21_12 ) : ( n11335 ) ;
assign n11337 =  ( n10638 ) ? ( VREG_21_13 ) : ( n11336 ) ;
assign n11338 =  ( n10637 ) ? ( VREG_21_14 ) : ( n11337 ) ;
assign n11339 =  ( n10636 ) ? ( VREG_21_15 ) : ( n11338 ) ;
assign n11340 =  ( n10635 ) ? ( VREG_22_0 ) : ( n11339 ) ;
assign n11341 =  ( n10634 ) ? ( VREG_22_1 ) : ( n11340 ) ;
assign n11342 =  ( n10633 ) ? ( VREG_22_2 ) : ( n11341 ) ;
assign n11343 =  ( n10632 ) ? ( VREG_22_3 ) : ( n11342 ) ;
assign n11344 =  ( n10631 ) ? ( VREG_22_4 ) : ( n11343 ) ;
assign n11345 =  ( n10630 ) ? ( VREG_22_5 ) : ( n11344 ) ;
assign n11346 =  ( n10629 ) ? ( VREG_22_6 ) : ( n11345 ) ;
assign n11347 =  ( n10628 ) ? ( VREG_22_7 ) : ( n11346 ) ;
assign n11348 =  ( n10627 ) ? ( VREG_22_8 ) : ( n11347 ) ;
assign n11349 =  ( n10626 ) ? ( VREG_22_9 ) : ( n11348 ) ;
assign n11350 =  ( n10625 ) ? ( VREG_22_10 ) : ( n11349 ) ;
assign n11351 =  ( n10624 ) ? ( VREG_22_11 ) : ( n11350 ) ;
assign n11352 =  ( n10623 ) ? ( VREG_22_12 ) : ( n11351 ) ;
assign n11353 =  ( n10622 ) ? ( VREG_22_13 ) : ( n11352 ) ;
assign n11354 =  ( n10621 ) ? ( VREG_22_14 ) : ( n11353 ) ;
assign n11355 =  ( n10620 ) ? ( VREG_22_15 ) : ( n11354 ) ;
assign n11356 =  ( n10619 ) ? ( VREG_23_0 ) : ( n11355 ) ;
assign n11357 =  ( n10618 ) ? ( VREG_23_1 ) : ( n11356 ) ;
assign n11358 =  ( n10617 ) ? ( VREG_23_2 ) : ( n11357 ) ;
assign n11359 =  ( n10616 ) ? ( VREG_23_3 ) : ( n11358 ) ;
assign n11360 =  ( n10615 ) ? ( VREG_23_4 ) : ( n11359 ) ;
assign n11361 =  ( n10614 ) ? ( VREG_23_5 ) : ( n11360 ) ;
assign n11362 =  ( n10613 ) ? ( VREG_23_6 ) : ( n11361 ) ;
assign n11363 =  ( n10612 ) ? ( VREG_23_7 ) : ( n11362 ) ;
assign n11364 =  ( n10611 ) ? ( VREG_23_8 ) : ( n11363 ) ;
assign n11365 =  ( n10610 ) ? ( VREG_23_9 ) : ( n11364 ) ;
assign n11366 =  ( n10609 ) ? ( VREG_23_10 ) : ( n11365 ) ;
assign n11367 =  ( n10608 ) ? ( VREG_23_11 ) : ( n11366 ) ;
assign n11368 =  ( n10607 ) ? ( VREG_23_12 ) : ( n11367 ) ;
assign n11369 =  ( n10606 ) ? ( VREG_23_13 ) : ( n11368 ) ;
assign n11370 =  ( n10605 ) ? ( VREG_23_14 ) : ( n11369 ) ;
assign n11371 =  ( n10604 ) ? ( VREG_23_15 ) : ( n11370 ) ;
assign n11372 =  ( n10603 ) ? ( VREG_24_0 ) : ( n11371 ) ;
assign n11373 =  ( n10602 ) ? ( VREG_24_1 ) : ( n11372 ) ;
assign n11374 =  ( n10601 ) ? ( VREG_24_2 ) : ( n11373 ) ;
assign n11375 =  ( n10600 ) ? ( VREG_24_3 ) : ( n11374 ) ;
assign n11376 =  ( n10599 ) ? ( VREG_24_4 ) : ( n11375 ) ;
assign n11377 =  ( n10598 ) ? ( VREG_24_5 ) : ( n11376 ) ;
assign n11378 =  ( n10597 ) ? ( VREG_24_6 ) : ( n11377 ) ;
assign n11379 =  ( n10596 ) ? ( VREG_24_7 ) : ( n11378 ) ;
assign n11380 =  ( n10595 ) ? ( VREG_24_8 ) : ( n11379 ) ;
assign n11381 =  ( n10594 ) ? ( VREG_24_9 ) : ( n11380 ) ;
assign n11382 =  ( n10593 ) ? ( VREG_24_10 ) : ( n11381 ) ;
assign n11383 =  ( n10592 ) ? ( VREG_24_11 ) : ( n11382 ) ;
assign n11384 =  ( n10591 ) ? ( VREG_24_12 ) : ( n11383 ) ;
assign n11385 =  ( n10590 ) ? ( VREG_24_13 ) : ( n11384 ) ;
assign n11386 =  ( n10589 ) ? ( VREG_24_14 ) : ( n11385 ) ;
assign n11387 =  ( n10588 ) ? ( VREG_24_15 ) : ( n11386 ) ;
assign n11388 =  ( n10587 ) ? ( VREG_25_0 ) : ( n11387 ) ;
assign n11389 =  ( n10586 ) ? ( VREG_25_1 ) : ( n11388 ) ;
assign n11390 =  ( n10585 ) ? ( VREG_25_2 ) : ( n11389 ) ;
assign n11391 =  ( n10584 ) ? ( VREG_25_3 ) : ( n11390 ) ;
assign n11392 =  ( n10583 ) ? ( VREG_25_4 ) : ( n11391 ) ;
assign n11393 =  ( n10582 ) ? ( VREG_25_5 ) : ( n11392 ) ;
assign n11394 =  ( n10581 ) ? ( VREG_25_6 ) : ( n11393 ) ;
assign n11395 =  ( n10580 ) ? ( VREG_25_7 ) : ( n11394 ) ;
assign n11396 =  ( n10579 ) ? ( VREG_25_8 ) : ( n11395 ) ;
assign n11397 =  ( n10578 ) ? ( VREG_25_9 ) : ( n11396 ) ;
assign n11398 =  ( n10577 ) ? ( VREG_25_10 ) : ( n11397 ) ;
assign n11399 =  ( n10576 ) ? ( VREG_25_11 ) : ( n11398 ) ;
assign n11400 =  ( n10575 ) ? ( VREG_25_12 ) : ( n11399 ) ;
assign n11401 =  ( n10574 ) ? ( VREG_25_13 ) : ( n11400 ) ;
assign n11402 =  ( n10573 ) ? ( VREG_25_14 ) : ( n11401 ) ;
assign n11403 =  ( n10572 ) ? ( VREG_25_15 ) : ( n11402 ) ;
assign n11404 =  ( n10571 ) ? ( VREG_26_0 ) : ( n11403 ) ;
assign n11405 =  ( n10570 ) ? ( VREG_26_1 ) : ( n11404 ) ;
assign n11406 =  ( n10569 ) ? ( VREG_26_2 ) : ( n11405 ) ;
assign n11407 =  ( n10568 ) ? ( VREG_26_3 ) : ( n11406 ) ;
assign n11408 =  ( n10567 ) ? ( VREG_26_4 ) : ( n11407 ) ;
assign n11409 =  ( n10566 ) ? ( VREG_26_5 ) : ( n11408 ) ;
assign n11410 =  ( n10565 ) ? ( VREG_26_6 ) : ( n11409 ) ;
assign n11411 =  ( n10564 ) ? ( VREG_26_7 ) : ( n11410 ) ;
assign n11412 =  ( n10563 ) ? ( VREG_26_8 ) : ( n11411 ) ;
assign n11413 =  ( n10562 ) ? ( VREG_26_9 ) : ( n11412 ) ;
assign n11414 =  ( n10561 ) ? ( VREG_26_10 ) : ( n11413 ) ;
assign n11415 =  ( n10560 ) ? ( VREG_26_11 ) : ( n11414 ) ;
assign n11416 =  ( n10559 ) ? ( VREG_26_12 ) : ( n11415 ) ;
assign n11417 =  ( n10558 ) ? ( VREG_26_13 ) : ( n11416 ) ;
assign n11418 =  ( n10557 ) ? ( VREG_26_14 ) : ( n11417 ) ;
assign n11419 =  ( n10556 ) ? ( VREG_26_15 ) : ( n11418 ) ;
assign n11420 =  ( n10555 ) ? ( VREG_27_0 ) : ( n11419 ) ;
assign n11421 =  ( n10554 ) ? ( VREG_27_1 ) : ( n11420 ) ;
assign n11422 =  ( n10553 ) ? ( VREG_27_2 ) : ( n11421 ) ;
assign n11423 =  ( n10552 ) ? ( VREG_27_3 ) : ( n11422 ) ;
assign n11424 =  ( n10551 ) ? ( VREG_27_4 ) : ( n11423 ) ;
assign n11425 =  ( n10550 ) ? ( VREG_27_5 ) : ( n11424 ) ;
assign n11426 =  ( n10549 ) ? ( VREG_27_6 ) : ( n11425 ) ;
assign n11427 =  ( n10548 ) ? ( VREG_27_7 ) : ( n11426 ) ;
assign n11428 =  ( n10547 ) ? ( VREG_27_8 ) : ( n11427 ) ;
assign n11429 =  ( n10546 ) ? ( VREG_27_9 ) : ( n11428 ) ;
assign n11430 =  ( n10545 ) ? ( VREG_27_10 ) : ( n11429 ) ;
assign n11431 =  ( n10544 ) ? ( VREG_27_11 ) : ( n11430 ) ;
assign n11432 =  ( n10543 ) ? ( VREG_27_12 ) : ( n11431 ) ;
assign n11433 =  ( n10542 ) ? ( VREG_27_13 ) : ( n11432 ) ;
assign n11434 =  ( n10541 ) ? ( VREG_27_14 ) : ( n11433 ) ;
assign n11435 =  ( n10540 ) ? ( VREG_27_15 ) : ( n11434 ) ;
assign n11436 =  ( n10539 ) ? ( VREG_28_0 ) : ( n11435 ) ;
assign n11437 =  ( n10538 ) ? ( VREG_28_1 ) : ( n11436 ) ;
assign n11438 =  ( n10537 ) ? ( VREG_28_2 ) : ( n11437 ) ;
assign n11439 =  ( n10536 ) ? ( VREG_28_3 ) : ( n11438 ) ;
assign n11440 =  ( n10535 ) ? ( VREG_28_4 ) : ( n11439 ) ;
assign n11441 =  ( n10534 ) ? ( VREG_28_5 ) : ( n11440 ) ;
assign n11442 =  ( n10533 ) ? ( VREG_28_6 ) : ( n11441 ) ;
assign n11443 =  ( n10532 ) ? ( VREG_28_7 ) : ( n11442 ) ;
assign n11444 =  ( n10531 ) ? ( VREG_28_8 ) : ( n11443 ) ;
assign n11445 =  ( n10530 ) ? ( VREG_28_9 ) : ( n11444 ) ;
assign n11446 =  ( n10529 ) ? ( VREG_28_10 ) : ( n11445 ) ;
assign n11447 =  ( n10528 ) ? ( VREG_28_11 ) : ( n11446 ) ;
assign n11448 =  ( n10527 ) ? ( VREG_28_12 ) : ( n11447 ) ;
assign n11449 =  ( n10526 ) ? ( VREG_28_13 ) : ( n11448 ) ;
assign n11450 =  ( n10525 ) ? ( VREG_28_14 ) : ( n11449 ) ;
assign n11451 =  ( n10524 ) ? ( VREG_28_15 ) : ( n11450 ) ;
assign n11452 =  ( n10523 ) ? ( VREG_29_0 ) : ( n11451 ) ;
assign n11453 =  ( n10522 ) ? ( VREG_29_1 ) : ( n11452 ) ;
assign n11454 =  ( n10521 ) ? ( VREG_29_2 ) : ( n11453 ) ;
assign n11455 =  ( n10520 ) ? ( VREG_29_3 ) : ( n11454 ) ;
assign n11456 =  ( n10519 ) ? ( VREG_29_4 ) : ( n11455 ) ;
assign n11457 =  ( n10518 ) ? ( VREG_29_5 ) : ( n11456 ) ;
assign n11458 =  ( n10517 ) ? ( VREG_29_6 ) : ( n11457 ) ;
assign n11459 =  ( n10516 ) ? ( VREG_29_7 ) : ( n11458 ) ;
assign n11460 =  ( n10515 ) ? ( VREG_29_8 ) : ( n11459 ) ;
assign n11461 =  ( n10514 ) ? ( VREG_29_9 ) : ( n11460 ) ;
assign n11462 =  ( n10513 ) ? ( VREG_29_10 ) : ( n11461 ) ;
assign n11463 =  ( n10512 ) ? ( VREG_29_11 ) : ( n11462 ) ;
assign n11464 =  ( n10511 ) ? ( VREG_29_12 ) : ( n11463 ) ;
assign n11465 =  ( n10510 ) ? ( VREG_29_13 ) : ( n11464 ) ;
assign n11466 =  ( n10509 ) ? ( VREG_29_14 ) : ( n11465 ) ;
assign n11467 =  ( n10508 ) ? ( VREG_29_15 ) : ( n11466 ) ;
assign n11468 =  ( n10507 ) ? ( VREG_30_0 ) : ( n11467 ) ;
assign n11469 =  ( n10506 ) ? ( VREG_30_1 ) : ( n11468 ) ;
assign n11470 =  ( n10505 ) ? ( VREG_30_2 ) : ( n11469 ) ;
assign n11471 =  ( n10504 ) ? ( VREG_30_3 ) : ( n11470 ) ;
assign n11472 =  ( n10503 ) ? ( VREG_30_4 ) : ( n11471 ) ;
assign n11473 =  ( n10502 ) ? ( VREG_30_5 ) : ( n11472 ) ;
assign n11474 =  ( n10501 ) ? ( VREG_30_6 ) : ( n11473 ) ;
assign n11475 =  ( n10500 ) ? ( VREG_30_7 ) : ( n11474 ) ;
assign n11476 =  ( n10499 ) ? ( VREG_30_8 ) : ( n11475 ) ;
assign n11477 =  ( n10498 ) ? ( VREG_30_9 ) : ( n11476 ) ;
assign n11478 =  ( n10497 ) ? ( VREG_30_10 ) : ( n11477 ) ;
assign n11479 =  ( n10496 ) ? ( VREG_30_11 ) : ( n11478 ) ;
assign n11480 =  ( n10495 ) ? ( VREG_30_12 ) : ( n11479 ) ;
assign n11481 =  ( n10494 ) ? ( VREG_30_13 ) : ( n11480 ) ;
assign n11482 =  ( n10493 ) ? ( VREG_30_14 ) : ( n11481 ) ;
assign n11483 =  ( n10492 ) ? ( VREG_30_15 ) : ( n11482 ) ;
assign n11484 =  ( n10491 ) ? ( VREG_31_0 ) : ( n11483 ) ;
assign n11485 =  ( n10490 ) ? ( VREG_31_1 ) : ( n11484 ) ;
assign n11486 =  ( n10489 ) ? ( VREG_31_2 ) : ( n11485 ) ;
assign n11487 =  ( n10488 ) ? ( VREG_31_3 ) : ( n11486 ) ;
assign n11488 =  ( n10487 ) ? ( VREG_31_4 ) : ( n11487 ) ;
assign n11489 =  ( n10486 ) ? ( VREG_31_5 ) : ( n11488 ) ;
assign n11490 =  ( n10485 ) ? ( VREG_31_6 ) : ( n11489 ) ;
assign n11491 =  ( n10484 ) ? ( VREG_31_7 ) : ( n11490 ) ;
assign n11492 =  ( n10483 ) ? ( VREG_31_8 ) : ( n11491 ) ;
assign n11493 =  ( n10482 ) ? ( VREG_31_9 ) : ( n11492 ) ;
assign n11494 =  ( n10481 ) ? ( VREG_31_10 ) : ( n11493 ) ;
assign n11495 =  ( n10480 ) ? ( VREG_31_11 ) : ( n11494 ) ;
assign n11496 =  ( n10479 ) ? ( VREG_31_12 ) : ( n11495 ) ;
assign n11497 =  ( n10478 ) ? ( VREG_31_13 ) : ( n11496 ) ;
assign n11498 =  ( n10477 ) ? ( VREG_31_14 ) : ( n11497 ) ;
assign n11499 =  ( n10476 ) ? ( VREG_31_15 ) : ( n11498 ) ;
assign n11500 =  ( n10465 ) + ( n11499 )  ;
assign n11501 =  ( n10465 ) - ( n11499 )  ;
assign n11502 =  ( n10465 ) & ( n11499 )  ;
assign n11503 =  ( n10465 ) | ( n11499 )  ;
assign n11504 =  ( ( n10465 ) * ( n11499 ))  ;
assign n11505 =  ( n148 ) ? ( n11504 ) : ( VREG_0_12 ) ;
assign n11506 =  ( n146 ) ? ( n11503 ) : ( n11505 ) ;
assign n11507 =  ( n144 ) ? ( n11502 ) : ( n11506 ) ;
assign n11508 =  ( n142 ) ? ( n11501 ) : ( n11507 ) ;
assign n11509 =  ( n10 ) ? ( n11500 ) : ( n11508 ) ;
assign n11510 = n3030[12:12] ;
assign n11511 =  ( n11510 ) == ( 1'd0 )  ;
assign n11512 =  ( n11511 ) ? ( VREG_0_12 ) : ( n10475 ) ;
assign n11513 =  ( n11511 ) ? ( VREG_0_12 ) : ( n11509 ) ;
assign n11514 =  ( n3034 ) ? ( n11513 ) : ( VREG_0_12 ) ;
assign n11515 =  ( n2965 ) ? ( n11512 ) : ( n11514 ) ;
assign n11516 =  ( n1930 ) ? ( n11509 ) : ( n11515 ) ;
assign n11517 =  ( n879 ) ? ( n10475 ) : ( n11516 ) ;
assign n11518 =  ( n10465 ) + ( n164 )  ;
assign n11519 =  ( n10465 ) - ( n164 )  ;
assign n11520 =  ( n10465 ) & ( n164 )  ;
assign n11521 =  ( n10465 ) | ( n164 )  ;
assign n11522 =  ( ( n10465 ) * ( n164 ))  ;
assign n11523 =  ( n172 ) ? ( n11522 ) : ( VREG_0_12 ) ;
assign n11524 =  ( n170 ) ? ( n11521 ) : ( n11523 ) ;
assign n11525 =  ( n168 ) ? ( n11520 ) : ( n11524 ) ;
assign n11526 =  ( n166 ) ? ( n11519 ) : ( n11525 ) ;
assign n11527 =  ( n162 ) ? ( n11518 ) : ( n11526 ) ;
assign n11528 =  ( n10465 ) + ( n180 )  ;
assign n11529 =  ( n10465 ) - ( n180 )  ;
assign n11530 =  ( n10465 ) & ( n180 )  ;
assign n11531 =  ( n10465 ) | ( n180 )  ;
assign n11532 =  ( ( n10465 ) * ( n180 ))  ;
assign n11533 =  ( n172 ) ? ( n11532 ) : ( VREG_0_12 ) ;
assign n11534 =  ( n170 ) ? ( n11531 ) : ( n11533 ) ;
assign n11535 =  ( n168 ) ? ( n11530 ) : ( n11534 ) ;
assign n11536 =  ( n166 ) ? ( n11529 ) : ( n11535 ) ;
assign n11537 =  ( n162 ) ? ( n11528 ) : ( n11536 ) ;
assign n11538 =  ( n11511 ) ? ( VREG_0_12 ) : ( n11537 ) ;
assign n11539 =  ( n3051 ) ? ( n11538 ) : ( VREG_0_12 ) ;
assign n11540 =  ( n3040 ) ? ( n11527 ) : ( n11539 ) ;
assign n11541 =  ( n192 ) ? ( VREG_0_12 ) : ( VREG_0_12 ) ;
assign n11542 =  ( n157 ) ? ( n11540 ) : ( n11541 ) ;
assign n11543 =  ( n6 ) ? ( n11517 ) : ( n11542 ) ;
assign n11544 =  ( n4 ) ? ( n11543 ) : ( VREG_0_12 ) ;
assign n11545 =  ( 32'd13 ) == ( 32'd15 )  ;
assign n11546 =  ( n12 ) & ( n11545 )  ;
assign n11547 =  ( 32'd13 ) == ( 32'd14 )  ;
assign n11548 =  ( n12 ) & ( n11547 )  ;
assign n11549 =  ( 32'd13 ) == ( 32'd13 )  ;
assign n11550 =  ( n12 ) & ( n11549 )  ;
assign n11551 =  ( 32'd13 ) == ( 32'd12 )  ;
assign n11552 =  ( n12 ) & ( n11551 )  ;
assign n11553 =  ( 32'd13 ) == ( 32'd11 )  ;
assign n11554 =  ( n12 ) & ( n11553 )  ;
assign n11555 =  ( 32'd13 ) == ( 32'd10 )  ;
assign n11556 =  ( n12 ) & ( n11555 )  ;
assign n11557 =  ( 32'd13 ) == ( 32'd9 )  ;
assign n11558 =  ( n12 ) & ( n11557 )  ;
assign n11559 =  ( 32'd13 ) == ( 32'd8 )  ;
assign n11560 =  ( n12 ) & ( n11559 )  ;
assign n11561 =  ( 32'd13 ) == ( 32'd7 )  ;
assign n11562 =  ( n12 ) & ( n11561 )  ;
assign n11563 =  ( 32'd13 ) == ( 32'd6 )  ;
assign n11564 =  ( n12 ) & ( n11563 )  ;
assign n11565 =  ( 32'd13 ) == ( 32'd5 )  ;
assign n11566 =  ( n12 ) & ( n11565 )  ;
assign n11567 =  ( 32'd13 ) == ( 32'd4 )  ;
assign n11568 =  ( n12 ) & ( n11567 )  ;
assign n11569 =  ( 32'd13 ) == ( 32'd3 )  ;
assign n11570 =  ( n12 ) & ( n11569 )  ;
assign n11571 =  ( 32'd13 ) == ( 32'd2 )  ;
assign n11572 =  ( n12 ) & ( n11571 )  ;
assign n11573 =  ( 32'd13 ) == ( 32'd1 )  ;
assign n11574 =  ( n12 ) & ( n11573 )  ;
assign n11575 =  ( 32'd13 ) == ( 32'd0 )  ;
assign n11576 =  ( n12 ) & ( n11575 )  ;
assign n11577 =  ( n13 ) & ( n11545 )  ;
assign n11578 =  ( n13 ) & ( n11547 )  ;
assign n11579 =  ( n13 ) & ( n11549 )  ;
assign n11580 =  ( n13 ) & ( n11551 )  ;
assign n11581 =  ( n13 ) & ( n11553 )  ;
assign n11582 =  ( n13 ) & ( n11555 )  ;
assign n11583 =  ( n13 ) & ( n11557 )  ;
assign n11584 =  ( n13 ) & ( n11559 )  ;
assign n11585 =  ( n13 ) & ( n11561 )  ;
assign n11586 =  ( n13 ) & ( n11563 )  ;
assign n11587 =  ( n13 ) & ( n11565 )  ;
assign n11588 =  ( n13 ) & ( n11567 )  ;
assign n11589 =  ( n13 ) & ( n11569 )  ;
assign n11590 =  ( n13 ) & ( n11571 )  ;
assign n11591 =  ( n13 ) & ( n11573 )  ;
assign n11592 =  ( n13 ) & ( n11575 )  ;
assign n11593 =  ( n14 ) & ( n11545 )  ;
assign n11594 =  ( n14 ) & ( n11547 )  ;
assign n11595 =  ( n14 ) & ( n11549 )  ;
assign n11596 =  ( n14 ) & ( n11551 )  ;
assign n11597 =  ( n14 ) & ( n11553 )  ;
assign n11598 =  ( n14 ) & ( n11555 )  ;
assign n11599 =  ( n14 ) & ( n11557 )  ;
assign n11600 =  ( n14 ) & ( n11559 )  ;
assign n11601 =  ( n14 ) & ( n11561 )  ;
assign n11602 =  ( n14 ) & ( n11563 )  ;
assign n11603 =  ( n14 ) & ( n11565 )  ;
assign n11604 =  ( n14 ) & ( n11567 )  ;
assign n11605 =  ( n14 ) & ( n11569 )  ;
assign n11606 =  ( n14 ) & ( n11571 )  ;
assign n11607 =  ( n14 ) & ( n11573 )  ;
assign n11608 =  ( n14 ) & ( n11575 )  ;
assign n11609 =  ( n15 ) & ( n11545 )  ;
assign n11610 =  ( n15 ) & ( n11547 )  ;
assign n11611 =  ( n15 ) & ( n11549 )  ;
assign n11612 =  ( n15 ) & ( n11551 )  ;
assign n11613 =  ( n15 ) & ( n11553 )  ;
assign n11614 =  ( n15 ) & ( n11555 )  ;
assign n11615 =  ( n15 ) & ( n11557 )  ;
assign n11616 =  ( n15 ) & ( n11559 )  ;
assign n11617 =  ( n15 ) & ( n11561 )  ;
assign n11618 =  ( n15 ) & ( n11563 )  ;
assign n11619 =  ( n15 ) & ( n11565 )  ;
assign n11620 =  ( n15 ) & ( n11567 )  ;
assign n11621 =  ( n15 ) & ( n11569 )  ;
assign n11622 =  ( n15 ) & ( n11571 )  ;
assign n11623 =  ( n15 ) & ( n11573 )  ;
assign n11624 =  ( n15 ) & ( n11575 )  ;
assign n11625 =  ( n16 ) & ( n11545 )  ;
assign n11626 =  ( n16 ) & ( n11547 )  ;
assign n11627 =  ( n16 ) & ( n11549 )  ;
assign n11628 =  ( n16 ) & ( n11551 )  ;
assign n11629 =  ( n16 ) & ( n11553 )  ;
assign n11630 =  ( n16 ) & ( n11555 )  ;
assign n11631 =  ( n16 ) & ( n11557 )  ;
assign n11632 =  ( n16 ) & ( n11559 )  ;
assign n11633 =  ( n16 ) & ( n11561 )  ;
assign n11634 =  ( n16 ) & ( n11563 )  ;
assign n11635 =  ( n16 ) & ( n11565 )  ;
assign n11636 =  ( n16 ) & ( n11567 )  ;
assign n11637 =  ( n16 ) & ( n11569 )  ;
assign n11638 =  ( n16 ) & ( n11571 )  ;
assign n11639 =  ( n16 ) & ( n11573 )  ;
assign n11640 =  ( n16 ) & ( n11575 )  ;
assign n11641 =  ( n17 ) & ( n11545 )  ;
assign n11642 =  ( n17 ) & ( n11547 )  ;
assign n11643 =  ( n17 ) & ( n11549 )  ;
assign n11644 =  ( n17 ) & ( n11551 )  ;
assign n11645 =  ( n17 ) & ( n11553 )  ;
assign n11646 =  ( n17 ) & ( n11555 )  ;
assign n11647 =  ( n17 ) & ( n11557 )  ;
assign n11648 =  ( n17 ) & ( n11559 )  ;
assign n11649 =  ( n17 ) & ( n11561 )  ;
assign n11650 =  ( n17 ) & ( n11563 )  ;
assign n11651 =  ( n17 ) & ( n11565 )  ;
assign n11652 =  ( n17 ) & ( n11567 )  ;
assign n11653 =  ( n17 ) & ( n11569 )  ;
assign n11654 =  ( n17 ) & ( n11571 )  ;
assign n11655 =  ( n17 ) & ( n11573 )  ;
assign n11656 =  ( n17 ) & ( n11575 )  ;
assign n11657 =  ( n18 ) & ( n11545 )  ;
assign n11658 =  ( n18 ) & ( n11547 )  ;
assign n11659 =  ( n18 ) & ( n11549 )  ;
assign n11660 =  ( n18 ) & ( n11551 )  ;
assign n11661 =  ( n18 ) & ( n11553 )  ;
assign n11662 =  ( n18 ) & ( n11555 )  ;
assign n11663 =  ( n18 ) & ( n11557 )  ;
assign n11664 =  ( n18 ) & ( n11559 )  ;
assign n11665 =  ( n18 ) & ( n11561 )  ;
assign n11666 =  ( n18 ) & ( n11563 )  ;
assign n11667 =  ( n18 ) & ( n11565 )  ;
assign n11668 =  ( n18 ) & ( n11567 )  ;
assign n11669 =  ( n18 ) & ( n11569 )  ;
assign n11670 =  ( n18 ) & ( n11571 )  ;
assign n11671 =  ( n18 ) & ( n11573 )  ;
assign n11672 =  ( n18 ) & ( n11575 )  ;
assign n11673 =  ( n19 ) & ( n11545 )  ;
assign n11674 =  ( n19 ) & ( n11547 )  ;
assign n11675 =  ( n19 ) & ( n11549 )  ;
assign n11676 =  ( n19 ) & ( n11551 )  ;
assign n11677 =  ( n19 ) & ( n11553 )  ;
assign n11678 =  ( n19 ) & ( n11555 )  ;
assign n11679 =  ( n19 ) & ( n11557 )  ;
assign n11680 =  ( n19 ) & ( n11559 )  ;
assign n11681 =  ( n19 ) & ( n11561 )  ;
assign n11682 =  ( n19 ) & ( n11563 )  ;
assign n11683 =  ( n19 ) & ( n11565 )  ;
assign n11684 =  ( n19 ) & ( n11567 )  ;
assign n11685 =  ( n19 ) & ( n11569 )  ;
assign n11686 =  ( n19 ) & ( n11571 )  ;
assign n11687 =  ( n19 ) & ( n11573 )  ;
assign n11688 =  ( n19 ) & ( n11575 )  ;
assign n11689 =  ( n20 ) & ( n11545 )  ;
assign n11690 =  ( n20 ) & ( n11547 )  ;
assign n11691 =  ( n20 ) & ( n11549 )  ;
assign n11692 =  ( n20 ) & ( n11551 )  ;
assign n11693 =  ( n20 ) & ( n11553 )  ;
assign n11694 =  ( n20 ) & ( n11555 )  ;
assign n11695 =  ( n20 ) & ( n11557 )  ;
assign n11696 =  ( n20 ) & ( n11559 )  ;
assign n11697 =  ( n20 ) & ( n11561 )  ;
assign n11698 =  ( n20 ) & ( n11563 )  ;
assign n11699 =  ( n20 ) & ( n11565 )  ;
assign n11700 =  ( n20 ) & ( n11567 )  ;
assign n11701 =  ( n20 ) & ( n11569 )  ;
assign n11702 =  ( n20 ) & ( n11571 )  ;
assign n11703 =  ( n20 ) & ( n11573 )  ;
assign n11704 =  ( n20 ) & ( n11575 )  ;
assign n11705 =  ( n21 ) & ( n11545 )  ;
assign n11706 =  ( n21 ) & ( n11547 )  ;
assign n11707 =  ( n21 ) & ( n11549 )  ;
assign n11708 =  ( n21 ) & ( n11551 )  ;
assign n11709 =  ( n21 ) & ( n11553 )  ;
assign n11710 =  ( n21 ) & ( n11555 )  ;
assign n11711 =  ( n21 ) & ( n11557 )  ;
assign n11712 =  ( n21 ) & ( n11559 )  ;
assign n11713 =  ( n21 ) & ( n11561 )  ;
assign n11714 =  ( n21 ) & ( n11563 )  ;
assign n11715 =  ( n21 ) & ( n11565 )  ;
assign n11716 =  ( n21 ) & ( n11567 )  ;
assign n11717 =  ( n21 ) & ( n11569 )  ;
assign n11718 =  ( n21 ) & ( n11571 )  ;
assign n11719 =  ( n21 ) & ( n11573 )  ;
assign n11720 =  ( n21 ) & ( n11575 )  ;
assign n11721 =  ( n22 ) & ( n11545 )  ;
assign n11722 =  ( n22 ) & ( n11547 )  ;
assign n11723 =  ( n22 ) & ( n11549 )  ;
assign n11724 =  ( n22 ) & ( n11551 )  ;
assign n11725 =  ( n22 ) & ( n11553 )  ;
assign n11726 =  ( n22 ) & ( n11555 )  ;
assign n11727 =  ( n22 ) & ( n11557 )  ;
assign n11728 =  ( n22 ) & ( n11559 )  ;
assign n11729 =  ( n22 ) & ( n11561 )  ;
assign n11730 =  ( n22 ) & ( n11563 )  ;
assign n11731 =  ( n22 ) & ( n11565 )  ;
assign n11732 =  ( n22 ) & ( n11567 )  ;
assign n11733 =  ( n22 ) & ( n11569 )  ;
assign n11734 =  ( n22 ) & ( n11571 )  ;
assign n11735 =  ( n22 ) & ( n11573 )  ;
assign n11736 =  ( n22 ) & ( n11575 )  ;
assign n11737 =  ( n23 ) & ( n11545 )  ;
assign n11738 =  ( n23 ) & ( n11547 )  ;
assign n11739 =  ( n23 ) & ( n11549 )  ;
assign n11740 =  ( n23 ) & ( n11551 )  ;
assign n11741 =  ( n23 ) & ( n11553 )  ;
assign n11742 =  ( n23 ) & ( n11555 )  ;
assign n11743 =  ( n23 ) & ( n11557 )  ;
assign n11744 =  ( n23 ) & ( n11559 )  ;
assign n11745 =  ( n23 ) & ( n11561 )  ;
assign n11746 =  ( n23 ) & ( n11563 )  ;
assign n11747 =  ( n23 ) & ( n11565 )  ;
assign n11748 =  ( n23 ) & ( n11567 )  ;
assign n11749 =  ( n23 ) & ( n11569 )  ;
assign n11750 =  ( n23 ) & ( n11571 )  ;
assign n11751 =  ( n23 ) & ( n11573 )  ;
assign n11752 =  ( n23 ) & ( n11575 )  ;
assign n11753 =  ( n24 ) & ( n11545 )  ;
assign n11754 =  ( n24 ) & ( n11547 )  ;
assign n11755 =  ( n24 ) & ( n11549 )  ;
assign n11756 =  ( n24 ) & ( n11551 )  ;
assign n11757 =  ( n24 ) & ( n11553 )  ;
assign n11758 =  ( n24 ) & ( n11555 )  ;
assign n11759 =  ( n24 ) & ( n11557 )  ;
assign n11760 =  ( n24 ) & ( n11559 )  ;
assign n11761 =  ( n24 ) & ( n11561 )  ;
assign n11762 =  ( n24 ) & ( n11563 )  ;
assign n11763 =  ( n24 ) & ( n11565 )  ;
assign n11764 =  ( n24 ) & ( n11567 )  ;
assign n11765 =  ( n24 ) & ( n11569 )  ;
assign n11766 =  ( n24 ) & ( n11571 )  ;
assign n11767 =  ( n24 ) & ( n11573 )  ;
assign n11768 =  ( n24 ) & ( n11575 )  ;
assign n11769 =  ( n25 ) & ( n11545 )  ;
assign n11770 =  ( n25 ) & ( n11547 )  ;
assign n11771 =  ( n25 ) & ( n11549 )  ;
assign n11772 =  ( n25 ) & ( n11551 )  ;
assign n11773 =  ( n25 ) & ( n11553 )  ;
assign n11774 =  ( n25 ) & ( n11555 )  ;
assign n11775 =  ( n25 ) & ( n11557 )  ;
assign n11776 =  ( n25 ) & ( n11559 )  ;
assign n11777 =  ( n25 ) & ( n11561 )  ;
assign n11778 =  ( n25 ) & ( n11563 )  ;
assign n11779 =  ( n25 ) & ( n11565 )  ;
assign n11780 =  ( n25 ) & ( n11567 )  ;
assign n11781 =  ( n25 ) & ( n11569 )  ;
assign n11782 =  ( n25 ) & ( n11571 )  ;
assign n11783 =  ( n25 ) & ( n11573 )  ;
assign n11784 =  ( n25 ) & ( n11575 )  ;
assign n11785 =  ( n26 ) & ( n11545 )  ;
assign n11786 =  ( n26 ) & ( n11547 )  ;
assign n11787 =  ( n26 ) & ( n11549 )  ;
assign n11788 =  ( n26 ) & ( n11551 )  ;
assign n11789 =  ( n26 ) & ( n11553 )  ;
assign n11790 =  ( n26 ) & ( n11555 )  ;
assign n11791 =  ( n26 ) & ( n11557 )  ;
assign n11792 =  ( n26 ) & ( n11559 )  ;
assign n11793 =  ( n26 ) & ( n11561 )  ;
assign n11794 =  ( n26 ) & ( n11563 )  ;
assign n11795 =  ( n26 ) & ( n11565 )  ;
assign n11796 =  ( n26 ) & ( n11567 )  ;
assign n11797 =  ( n26 ) & ( n11569 )  ;
assign n11798 =  ( n26 ) & ( n11571 )  ;
assign n11799 =  ( n26 ) & ( n11573 )  ;
assign n11800 =  ( n26 ) & ( n11575 )  ;
assign n11801 =  ( n27 ) & ( n11545 )  ;
assign n11802 =  ( n27 ) & ( n11547 )  ;
assign n11803 =  ( n27 ) & ( n11549 )  ;
assign n11804 =  ( n27 ) & ( n11551 )  ;
assign n11805 =  ( n27 ) & ( n11553 )  ;
assign n11806 =  ( n27 ) & ( n11555 )  ;
assign n11807 =  ( n27 ) & ( n11557 )  ;
assign n11808 =  ( n27 ) & ( n11559 )  ;
assign n11809 =  ( n27 ) & ( n11561 )  ;
assign n11810 =  ( n27 ) & ( n11563 )  ;
assign n11811 =  ( n27 ) & ( n11565 )  ;
assign n11812 =  ( n27 ) & ( n11567 )  ;
assign n11813 =  ( n27 ) & ( n11569 )  ;
assign n11814 =  ( n27 ) & ( n11571 )  ;
assign n11815 =  ( n27 ) & ( n11573 )  ;
assign n11816 =  ( n27 ) & ( n11575 )  ;
assign n11817 =  ( n28 ) & ( n11545 )  ;
assign n11818 =  ( n28 ) & ( n11547 )  ;
assign n11819 =  ( n28 ) & ( n11549 )  ;
assign n11820 =  ( n28 ) & ( n11551 )  ;
assign n11821 =  ( n28 ) & ( n11553 )  ;
assign n11822 =  ( n28 ) & ( n11555 )  ;
assign n11823 =  ( n28 ) & ( n11557 )  ;
assign n11824 =  ( n28 ) & ( n11559 )  ;
assign n11825 =  ( n28 ) & ( n11561 )  ;
assign n11826 =  ( n28 ) & ( n11563 )  ;
assign n11827 =  ( n28 ) & ( n11565 )  ;
assign n11828 =  ( n28 ) & ( n11567 )  ;
assign n11829 =  ( n28 ) & ( n11569 )  ;
assign n11830 =  ( n28 ) & ( n11571 )  ;
assign n11831 =  ( n28 ) & ( n11573 )  ;
assign n11832 =  ( n28 ) & ( n11575 )  ;
assign n11833 =  ( n29 ) & ( n11545 )  ;
assign n11834 =  ( n29 ) & ( n11547 )  ;
assign n11835 =  ( n29 ) & ( n11549 )  ;
assign n11836 =  ( n29 ) & ( n11551 )  ;
assign n11837 =  ( n29 ) & ( n11553 )  ;
assign n11838 =  ( n29 ) & ( n11555 )  ;
assign n11839 =  ( n29 ) & ( n11557 )  ;
assign n11840 =  ( n29 ) & ( n11559 )  ;
assign n11841 =  ( n29 ) & ( n11561 )  ;
assign n11842 =  ( n29 ) & ( n11563 )  ;
assign n11843 =  ( n29 ) & ( n11565 )  ;
assign n11844 =  ( n29 ) & ( n11567 )  ;
assign n11845 =  ( n29 ) & ( n11569 )  ;
assign n11846 =  ( n29 ) & ( n11571 )  ;
assign n11847 =  ( n29 ) & ( n11573 )  ;
assign n11848 =  ( n29 ) & ( n11575 )  ;
assign n11849 =  ( n30 ) & ( n11545 )  ;
assign n11850 =  ( n30 ) & ( n11547 )  ;
assign n11851 =  ( n30 ) & ( n11549 )  ;
assign n11852 =  ( n30 ) & ( n11551 )  ;
assign n11853 =  ( n30 ) & ( n11553 )  ;
assign n11854 =  ( n30 ) & ( n11555 )  ;
assign n11855 =  ( n30 ) & ( n11557 )  ;
assign n11856 =  ( n30 ) & ( n11559 )  ;
assign n11857 =  ( n30 ) & ( n11561 )  ;
assign n11858 =  ( n30 ) & ( n11563 )  ;
assign n11859 =  ( n30 ) & ( n11565 )  ;
assign n11860 =  ( n30 ) & ( n11567 )  ;
assign n11861 =  ( n30 ) & ( n11569 )  ;
assign n11862 =  ( n30 ) & ( n11571 )  ;
assign n11863 =  ( n30 ) & ( n11573 )  ;
assign n11864 =  ( n30 ) & ( n11575 )  ;
assign n11865 =  ( n31 ) & ( n11545 )  ;
assign n11866 =  ( n31 ) & ( n11547 )  ;
assign n11867 =  ( n31 ) & ( n11549 )  ;
assign n11868 =  ( n31 ) & ( n11551 )  ;
assign n11869 =  ( n31 ) & ( n11553 )  ;
assign n11870 =  ( n31 ) & ( n11555 )  ;
assign n11871 =  ( n31 ) & ( n11557 )  ;
assign n11872 =  ( n31 ) & ( n11559 )  ;
assign n11873 =  ( n31 ) & ( n11561 )  ;
assign n11874 =  ( n31 ) & ( n11563 )  ;
assign n11875 =  ( n31 ) & ( n11565 )  ;
assign n11876 =  ( n31 ) & ( n11567 )  ;
assign n11877 =  ( n31 ) & ( n11569 )  ;
assign n11878 =  ( n31 ) & ( n11571 )  ;
assign n11879 =  ( n31 ) & ( n11573 )  ;
assign n11880 =  ( n31 ) & ( n11575 )  ;
assign n11881 =  ( n32 ) & ( n11545 )  ;
assign n11882 =  ( n32 ) & ( n11547 )  ;
assign n11883 =  ( n32 ) & ( n11549 )  ;
assign n11884 =  ( n32 ) & ( n11551 )  ;
assign n11885 =  ( n32 ) & ( n11553 )  ;
assign n11886 =  ( n32 ) & ( n11555 )  ;
assign n11887 =  ( n32 ) & ( n11557 )  ;
assign n11888 =  ( n32 ) & ( n11559 )  ;
assign n11889 =  ( n32 ) & ( n11561 )  ;
assign n11890 =  ( n32 ) & ( n11563 )  ;
assign n11891 =  ( n32 ) & ( n11565 )  ;
assign n11892 =  ( n32 ) & ( n11567 )  ;
assign n11893 =  ( n32 ) & ( n11569 )  ;
assign n11894 =  ( n32 ) & ( n11571 )  ;
assign n11895 =  ( n32 ) & ( n11573 )  ;
assign n11896 =  ( n32 ) & ( n11575 )  ;
assign n11897 =  ( n33 ) & ( n11545 )  ;
assign n11898 =  ( n33 ) & ( n11547 )  ;
assign n11899 =  ( n33 ) & ( n11549 )  ;
assign n11900 =  ( n33 ) & ( n11551 )  ;
assign n11901 =  ( n33 ) & ( n11553 )  ;
assign n11902 =  ( n33 ) & ( n11555 )  ;
assign n11903 =  ( n33 ) & ( n11557 )  ;
assign n11904 =  ( n33 ) & ( n11559 )  ;
assign n11905 =  ( n33 ) & ( n11561 )  ;
assign n11906 =  ( n33 ) & ( n11563 )  ;
assign n11907 =  ( n33 ) & ( n11565 )  ;
assign n11908 =  ( n33 ) & ( n11567 )  ;
assign n11909 =  ( n33 ) & ( n11569 )  ;
assign n11910 =  ( n33 ) & ( n11571 )  ;
assign n11911 =  ( n33 ) & ( n11573 )  ;
assign n11912 =  ( n33 ) & ( n11575 )  ;
assign n11913 =  ( n34 ) & ( n11545 )  ;
assign n11914 =  ( n34 ) & ( n11547 )  ;
assign n11915 =  ( n34 ) & ( n11549 )  ;
assign n11916 =  ( n34 ) & ( n11551 )  ;
assign n11917 =  ( n34 ) & ( n11553 )  ;
assign n11918 =  ( n34 ) & ( n11555 )  ;
assign n11919 =  ( n34 ) & ( n11557 )  ;
assign n11920 =  ( n34 ) & ( n11559 )  ;
assign n11921 =  ( n34 ) & ( n11561 )  ;
assign n11922 =  ( n34 ) & ( n11563 )  ;
assign n11923 =  ( n34 ) & ( n11565 )  ;
assign n11924 =  ( n34 ) & ( n11567 )  ;
assign n11925 =  ( n34 ) & ( n11569 )  ;
assign n11926 =  ( n34 ) & ( n11571 )  ;
assign n11927 =  ( n34 ) & ( n11573 )  ;
assign n11928 =  ( n34 ) & ( n11575 )  ;
assign n11929 =  ( n35 ) & ( n11545 )  ;
assign n11930 =  ( n35 ) & ( n11547 )  ;
assign n11931 =  ( n35 ) & ( n11549 )  ;
assign n11932 =  ( n35 ) & ( n11551 )  ;
assign n11933 =  ( n35 ) & ( n11553 )  ;
assign n11934 =  ( n35 ) & ( n11555 )  ;
assign n11935 =  ( n35 ) & ( n11557 )  ;
assign n11936 =  ( n35 ) & ( n11559 )  ;
assign n11937 =  ( n35 ) & ( n11561 )  ;
assign n11938 =  ( n35 ) & ( n11563 )  ;
assign n11939 =  ( n35 ) & ( n11565 )  ;
assign n11940 =  ( n35 ) & ( n11567 )  ;
assign n11941 =  ( n35 ) & ( n11569 )  ;
assign n11942 =  ( n35 ) & ( n11571 )  ;
assign n11943 =  ( n35 ) & ( n11573 )  ;
assign n11944 =  ( n35 ) & ( n11575 )  ;
assign n11945 =  ( n36 ) & ( n11545 )  ;
assign n11946 =  ( n36 ) & ( n11547 )  ;
assign n11947 =  ( n36 ) & ( n11549 )  ;
assign n11948 =  ( n36 ) & ( n11551 )  ;
assign n11949 =  ( n36 ) & ( n11553 )  ;
assign n11950 =  ( n36 ) & ( n11555 )  ;
assign n11951 =  ( n36 ) & ( n11557 )  ;
assign n11952 =  ( n36 ) & ( n11559 )  ;
assign n11953 =  ( n36 ) & ( n11561 )  ;
assign n11954 =  ( n36 ) & ( n11563 )  ;
assign n11955 =  ( n36 ) & ( n11565 )  ;
assign n11956 =  ( n36 ) & ( n11567 )  ;
assign n11957 =  ( n36 ) & ( n11569 )  ;
assign n11958 =  ( n36 ) & ( n11571 )  ;
assign n11959 =  ( n36 ) & ( n11573 )  ;
assign n11960 =  ( n36 ) & ( n11575 )  ;
assign n11961 =  ( n37 ) & ( n11545 )  ;
assign n11962 =  ( n37 ) & ( n11547 )  ;
assign n11963 =  ( n37 ) & ( n11549 )  ;
assign n11964 =  ( n37 ) & ( n11551 )  ;
assign n11965 =  ( n37 ) & ( n11553 )  ;
assign n11966 =  ( n37 ) & ( n11555 )  ;
assign n11967 =  ( n37 ) & ( n11557 )  ;
assign n11968 =  ( n37 ) & ( n11559 )  ;
assign n11969 =  ( n37 ) & ( n11561 )  ;
assign n11970 =  ( n37 ) & ( n11563 )  ;
assign n11971 =  ( n37 ) & ( n11565 )  ;
assign n11972 =  ( n37 ) & ( n11567 )  ;
assign n11973 =  ( n37 ) & ( n11569 )  ;
assign n11974 =  ( n37 ) & ( n11571 )  ;
assign n11975 =  ( n37 ) & ( n11573 )  ;
assign n11976 =  ( n37 ) & ( n11575 )  ;
assign n11977 =  ( n38 ) & ( n11545 )  ;
assign n11978 =  ( n38 ) & ( n11547 )  ;
assign n11979 =  ( n38 ) & ( n11549 )  ;
assign n11980 =  ( n38 ) & ( n11551 )  ;
assign n11981 =  ( n38 ) & ( n11553 )  ;
assign n11982 =  ( n38 ) & ( n11555 )  ;
assign n11983 =  ( n38 ) & ( n11557 )  ;
assign n11984 =  ( n38 ) & ( n11559 )  ;
assign n11985 =  ( n38 ) & ( n11561 )  ;
assign n11986 =  ( n38 ) & ( n11563 )  ;
assign n11987 =  ( n38 ) & ( n11565 )  ;
assign n11988 =  ( n38 ) & ( n11567 )  ;
assign n11989 =  ( n38 ) & ( n11569 )  ;
assign n11990 =  ( n38 ) & ( n11571 )  ;
assign n11991 =  ( n38 ) & ( n11573 )  ;
assign n11992 =  ( n38 ) & ( n11575 )  ;
assign n11993 =  ( n39 ) & ( n11545 )  ;
assign n11994 =  ( n39 ) & ( n11547 )  ;
assign n11995 =  ( n39 ) & ( n11549 )  ;
assign n11996 =  ( n39 ) & ( n11551 )  ;
assign n11997 =  ( n39 ) & ( n11553 )  ;
assign n11998 =  ( n39 ) & ( n11555 )  ;
assign n11999 =  ( n39 ) & ( n11557 )  ;
assign n12000 =  ( n39 ) & ( n11559 )  ;
assign n12001 =  ( n39 ) & ( n11561 )  ;
assign n12002 =  ( n39 ) & ( n11563 )  ;
assign n12003 =  ( n39 ) & ( n11565 )  ;
assign n12004 =  ( n39 ) & ( n11567 )  ;
assign n12005 =  ( n39 ) & ( n11569 )  ;
assign n12006 =  ( n39 ) & ( n11571 )  ;
assign n12007 =  ( n39 ) & ( n11573 )  ;
assign n12008 =  ( n39 ) & ( n11575 )  ;
assign n12009 =  ( n40 ) & ( n11545 )  ;
assign n12010 =  ( n40 ) & ( n11547 )  ;
assign n12011 =  ( n40 ) & ( n11549 )  ;
assign n12012 =  ( n40 ) & ( n11551 )  ;
assign n12013 =  ( n40 ) & ( n11553 )  ;
assign n12014 =  ( n40 ) & ( n11555 )  ;
assign n12015 =  ( n40 ) & ( n11557 )  ;
assign n12016 =  ( n40 ) & ( n11559 )  ;
assign n12017 =  ( n40 ) & ( n11561 )  ;
assign n12018 =  ( n40 ) & ( n11563 )  ;
assign n12019 =  ( n40 ) & ( n11565 )  ;
assign n12020 =  ( n40 ) & ( n11567 )  ;
assign n12021 =  ( n40 ) & ( n11569 )  ;
assign n12022 =  ( n40 ) & ( n11571 )  ;
assign n12023 =  ( n40 ) & ( n11573 )  ;
assign n12024 =  ( n40 ) & ( n11575 )  ;
assign n12025 =  ( n41 ) & ( n11545 )  ;
assign n12026 =  ( n41 ) & ( n11547 )  ;
assign n12027 =  ( n41 ) & ( n11549 )  ;
assign n12028 =  ( n41 ) & ( n11551 )  ;
assign n12029 =  ( n41 ) & ( n11553 )  ;
assign n12030 =  ( n41 ) & ( n11555 )  ;
assign n12031 =  ( n41 ) & ( n11557 )  ;
assign n12032 =  ( n41 ) & ( n11559 )  ;
assign n12033 =  ( n41 ) & ( n11561 )  ;
assign n12034 =  ( n41 ) & ( n11563 )  ;
assign n12035 =  ( n41 ) & ( n11565 )  ;
assign n12036 =  ( n41 ) & ( n11567 )  ;
assign n12037 =  ( n41 ) & ( n11569 )  ;
assign n12038 =  ( n41 ) & ( n11571 )  ;
assign n12039 =  ( n41 ) & ( n11573 )  ;
assign n12040 =  ( n41 ) & ( n11575 )  ;
assign n12041 =  ( n42 ) & ( n11545 )  ;
assign n12042 =  ( n42 ) & ( n11547 )  ;
assign n12043 =  ( n42 ) & ( n11549 )  ;
assign n12044 =  ( n42 ) & ( n11551 )  ;
assign n12045 =  ( n42 ) & ( n11553 )  ;
assign n12046 =  ( n42 ) & ( n11555 )  ;
assign n12047 =  ( n42 ) & ( n11557 )  ;
assign n12048 =  ( n42 ) & ( n11559 )  ;
assign n12049 =  ( n42 ) & ( n11561 )  ;
assign n12050 =  ( n42 ) & ( n11563 )  ;
assign n12051 =  ( n42 ) & ( n11565 )  ;
assign n12052 =  ( n42 ) & ( n11567 )  ;
assign n12053 =  ( n42 ) & ( n11569 )  ;
assign n12054 =  ( n42 ) & ( n11571 )  ;
assign n12055 =  ( n42 ) & ( n11573 )  ;
assign n12056 =  ( n42 ) & ( n11575 )  ;
assign n12057 =  ( n43 ) & ( n11545 )  ;
assign n12058 =  ( n43 ) & ( n11547 )  ;
assign n12059 =  ( n43 ) & ( n11549 )  ;
assign n12060 =  ( n43 ) & ( n11551 )  ;
assign n12061 =  ( n43 ) & ( n11553 )  ;
assign n12062 =  ( n43 ) & ( n11555 )  ;
assign n12063 =  ( n43 ) & ( n11557 )  ;
assign n12064 =  ( n43 ) & ( n11559 )  ;
assign n12065 =  ( n43 ) & ( n11561 )  ;
assign n12066 =  ( n43 ) & ( n11563 )  ;
assign n12067 =  ( n43 ) & ( n11565 )  ;
assign n12068 =  ( n43 ) & ( n11567 )  ;
assign n12069 =  ( n43 ) & ( n11569 )  ;
assign n12070 =  ( n43 ) & ( n11571 )  ;
assign n12071 =  ( n43 ) & ( n11573 )  ;
assign n12072 =  ( n43 ) & ( n11575 )  ;
assign n12073 =  ( n12072 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n12074 =  ( n12071 ) ? ( VREG_0_1 ) : ( n12073 ) ;
assign n12075 =  ( n12070 ) ? ( VREG_0_2 ) : ( n12074 ) ;
assign n12076 =  ( n12069 ) ? ( VREG_0_3 ) : ( n12075 ) ;
assign n12077 =  ( n12068 ) ? ( VREG_0_4 ) : ( n12076 ) ;
assign n12078 =  ( n12067 ) ? ( VREG_0_5 ) : ( n12077 ) ;
assign n12079 =  ( n12066 ) ? ( VREG_0_6 ) : ( n12078 ) ;
assign n12080 =  ( n12065 ) ? ( VREG_0_7 ) : ( n12079 ) ;
assign n12081 =  ( n12064 ) ? ( VREG_0_8 ) : ( n12080 ) ;
assign n12082 =  ( n12063 ) ? ( VREG_0_9 ) : ( n12081 ) ;
assign n12083 =  ( n12062 ) ? ( VREG_0_10 ) : ( n12082 ) ;
assign n12084 =  ( n12061 ) ? ( VREG_0_11 ) : ( n12083 ) ;
assign n12085 =  ( n12060 ) ? ( VREG_0_12 ) : ( n12084 ) ;
assign n12086 =  ( n12059 ) ? ( VREG_0_13 ) : ( n12085 ) ;
assign n12087 =  ( n12058 ) ? ( VREG_0_14 ) : ( n12086 ) ;
assign n12088 =  ( n12057 ) ? ( VREG_0_15 ) : ( n12087 ) ;
assign n12089 =  ( n12056 ) ? ( VREG_1_0 ) : ( n12088 ) ;
assign n12090 =  ( n12055 ) ? ( VREG_1_1 ) : ( n12089 ) ;
assign n12091 =  ( n12054 ) ? ( VREG_1_2 ) : ( n12090 ) ;
assign n12092 =  ( n12053 ) ? ( VREG_1_3 ) : ( n12091 ) ;
assign n12093 =  ( n12052 ) ? ( VREG_1_4 ) : ( n12092 ) ;
assign n12094 =  ( n12051 ) ? ( VREG_1_5 ) : ( n12093 ) ;
assign n12095 =  ( n12050 ) ? ( VREG_1_6 ) : ( n12094 ) ;
assign n12096 =  ( n12049 ) ? ( VREG_1_7 ) : ( n12095 ) ;
assign n12097 =  ( n12048 ) ? ( VREG_1_8 ) : ( n12096 ) ;
assign n12098 =  ( n12047 ) ? ( VREG_1_9 ) : ( n12097 ) ;
assign n12099 =  ( n12046 ) ? ( VREG_1_10 ) : ( n12098 ) ;
assign n12100 =  ( n12045 ) ? ( VREG_1_11 ) : ( n12099 ) ;
assign n12101 =  ( n12044 ) ? ( VREG_1_12 ) : ( n12100 ) ;
assign n12102 =  ( n12043 ) ? ( VREG_1_13 ) : ( n12101 ) ;
assign n12103 =  ( n12042 ) ? ( VREG_1_14 ) : ( n12102 ) ;
assign n12104 =  ( n12041 ) ? ( VREG_1_15 ) : ( n12103 ) ;
assign n12105 =  ( n12040 ) ? ( VREG_2_0 ) : ( n12104 ) ;
assign n12106 =  ( n12039 ) ? ( VREG_2_1 ) : ( n12105 ) ;
assign n12107 =  ( n12038 ) ? ( VREG_2_2 ) : ( n12106 ) ;
assign n12108 =  ( n12037 ) ? ( VREG_2_3 ) : ( n12107 ) ;
assign n12109 =  ( n12036 ) ? ( VREG_2_4 ) : ( n12108 ) ;
assign n12110 =  ( n12035 ) ? ( VREG_2_5 ) : ( n12109 ) ;
assign n12111 =  ( n12034 ) ? ( VREG_2_6 ) : ( n12110 ) ;
assign n12112 =  ( n12033 ) ? ( VREG_2_7 ) : ( n12111 ) ;
assign n12113 =  ( n12032 ) ? ( VREG_2_8 ) : ( n12112 ) ;
assign n12114 =  ( n12031 ) ? ( VREG_2_9 ) : ( n12113 ) ;
assign n12115 =  ( n12030 ) ? ( VREG_2_10 ) : ( n12114 ) ;
assign n12116 =  ( n12029 ) ? ( VREG_2_11 ) : ( n12115 ) ;
assign n12117 =  ( n12028 ) ? ( VREG_2_12 ) : ( n12116 ) ;
assign n12118 =  ( n12027 ) ? ( VREG_2_13 ) : ( n12117 ) ;
assign n12119 =  ( n12026 ) ? ( VREG_2_14 ) : ( n12118 ) ;
assign n12120 =  ( n12025 ) ? ( VREG_2_15 ) : ( n12119 ) ;
assign n12121 =  ( n12024 ) ? ( VREG_3_0 ) : ( n12120 ) ;
assign n12122 =  ( n12023 ) ? ( VREG_3_1 ) : ( n12121 ) ;
assign n12123 =  ( n12022 ) ? ( VREG_3_2 ) : ( n12122 ) ;
assign n12124 =  ( n12021 ) ? ( VREG_3_3 ) : ( n12123 ) ;
assign n12125 =  ( n12020 ) ? ( VREG_3_4 ) : ( n12124 ) ;
assign n12126 =  ( n12019 ) ? ( VREG_3_5 ) : ( n12125 ) ;
assign n12127 =  ( n12018 ) ? ( VREG_3_6 ) : ( n12126 ) ;
assign n12128 =  ( n12017 ) ? ( VREG_3_7 ) : ( n12127 ) ;
assign n12129 =  ( n12016 ) ? ( VREG_3_8 ) : ( n12128 ) ;
assign n12130 =  ( n12015 ) ? ( VREG_3_9 ) : ( n12129 ) ;
assign n12131 =  ( n12014 ) ? ( VREG_3_10 ) : ( n12130 ) ;
assign n12132 =  ( n12013 ) ? ( VREG_3_11 ) : ( n12131 ) ;
assign n12133 =  ( n12012 ) ? ( VREG_3_12 ) : ( n12132 ) ;
assign n12134 =  ( n12011 ) ? ( VREG_3_13 ) : ( n12133 ) ;
assign n12135 =  ( n12010 ) ? ( VREG_3_14 ) : ( n12134 ) ;
assign n12136 =  ( n12009 ) ? ( VREG_3_15 ) : ( n12135 ) ;
assign n12137 =  ( n12008 ) ? ( VREG_4_0 ) : ( n12136 ) ;
assign n12138 =  ( n12007 ) ? ( VREG_4_1 ) : ( n12137 ) ;
assign n12139 =  ( n12006 ) ? ( VREG_4_2 ) : ( n12138 ) ;
assign n12140 =  ( n12005 ) ? ( VREG_4_3 ) : ( n12139 ) ;
assign n12141 =  ( n12004 ) ? ( VREG_4_4 ) : ( n12140 ) ;
assign n12142 =  ( n12003 ) ? ( VREG_4_5 ) : ( n12141 ) ;
assign n12143 =  ( n12002 ) ? ( VREG_4_6 ) : ( n12142 ) ;
assign n12144 =  ( n12001 ) ? ( VREG_4_7 ) : ( n12143 ) ;
assign n12145 =  ( n12000 ) ? ( VREG_4_8 ) : ( n12144 ) ;
assign n12146 =  ( n11999 ) ? ( VREG_4_9 ) : ( n12145 ) ;
assign n12147 =  ( n11998 ) ? ( VREG_4_10 ) : ( n12146 ) ;
assign n12148 =  ( n11997 ) ? ( VREG_4_11 ) : ( n12147 ) ;
assign n12149 =  ( n11996 ) ? ( VREG_4_12 ) : ( n12148 ) ;
assign n12150 =  ( n11995 ) ? ( VREG_4_13 ) : ( n12149 ) ;
assign n12151 =  ( n11994 ) ? ( VREG_4_14 ) : ( n12150 ) ;
assign n12152 =  ( n11993 ) ? ( VREG_4_15 ) : ( n12151 ) ;
assign n12153 =  ( n11992 ) ? ( VREG_5_0 ) : ( n12152 ) ;
assign n12154 =  ( n11991 ) ? ( VREG_5_1 ) : ( n12153 ) ;
assign n12155 =  ( n11990 ) ? ( VREG_5_2 ) : ( n12154 ) ;
assign n12156 =  ( n11989 ) ? ( VREG_5_3 ) : ( n12155 ) ;
assign n12157 =  ( n11988 ) ? ( VREG_5_4 ) : ( n12156 ) ;
assign n12158 =  ( n11987 ) ? ( VREG_5_5 ) : ( n12157 ) ;
assign n12159 =  ( n11986 ) ? ( VREG_5_6 ) : ( n12158 ) ;
assign n12160 =  ( n11985 ) ? ( VREG_5_7 ) : ( n12159 ) ;
assign n12161 =  ( n11984 ) ? ( VREG_5_8 ) : ( n12160 ) ;
assign n12162 =  ( n11983 ) ? ( VREG_5_9 ) : ( n12161 ) ;
assign n12163 =  ( n11982 ) ? ( VREG_5_10 ) : ( n12162 ) ;
assign n12164 =  ( n11981 ) ? ( VREG_5_11 ) : ( n12163 ) ;
assign n12165 =  ( n11980 ) ? ( VREG_5_12 ) : ( n12164 ) ;
assign n12166 =  ( n11979 ) ? ( VREG_5_13 ) : ( n12165 ) ;
assign n12167 =  ( n11978 ) ? ( VREG_5_14 ) : ( n12166 ) ;
assign n12168 =  ( n11977 ) ? ( VREG_5_15 ) : ( n12167 ) ;
assign n12169 =  ( n11976 ) ? ( VREG_6_0 ) : ( n12168 ) ;
assign n12170 =  ( n11975 ) ? ( VREG_6_1 ) : ( n12169 ) ;
assign n12171 =  ( n11974 ) ? ( VREG_6_2 ) : ( n12170 ) ;
assign n12172 =  ( n11973 ) ? ( VREG_6_3 ) : ( n12171 ) ;
assign n12173 =  ( n11972 ) ? ( VREG_6_4 ) : ( n12172 ) ;
assign n12174 =  ( n11971 ) ? ( VREG_6_5 ) : ( n12173 ) ;
assign n12175 =  ( n11970 ) ? ( VREG_6_6 ) : ( n12174 ) ;
assign n12176 =  ( n11969 ) ? ( VREG_6_7 ) : ( n12175 ) ;
assign n12177 =  ( n11968 ) ? ( VREG_6_8 ) : ( n12176 ) ;
assign n12178 =  ( n11967 ) ? ( VREG_6_9 ) : ( n12177 ) ;
assign n12179 =  ( n11966 ) ? ( VREG_6_10 ) : ( n12178 ) ;
assign n12180 =  ( n11965 ) ? ( VREG_6_11 ) : ( n12179 ) ;
assign n12181 =  ( n11964 ) ? ( VREG_6_12 ) : ( n12180 ) ;
assign n12182 =  ( n11963 ) ? ( VREG_6_13 ) : ( n12181 ) ;
assign n12183 =  ( n11962 ) ? ( VREG_6_14 ) : ( n12182 ) ;
assign n12184 =  ( n11961 ) ? ( VREG_6_15 ) : ( n12183 ) ;
assign n12185 =  ( n11960 ) ? ( VREG_7_0 ) : ( n12184 ) ;
assign n12186 =  ( n11959 ) ? ( VREG_7_1 ) : ( n12185 ) ;
assign n12187 =  ( n11958 ) ? ( VREG_7_2 ) : ( n12186 ) ;
assign n12188 =  ( n11957 ) ? ( VREG_7_3 ) : ( n12187 ) ;
assign n12189 =  ( n11956 ) ? ( VREG_7_4 ) : ( n12188 ) ;
assign n12190 =  ( n11955 ) ? ( VREG_7_5 ) : ( n12189 ) ;
assign n12191 =  ( n11954 ) ? ( VREG_7_6 ) : ( n12190 ) ;
assign n12192 =  ( n11953 ) ? ( VREG_7_7 ) : ( n12191 ) ;
assign n12193 =  ( n11952 ) ? ( VREG_7_8 ) : ( n12192 ) ;
assign n12194 =  ( n11951 ) ? ( VREG_7_9 ) : ( n12193 ) ;
assign n12195 =  ( n11950 ) ? ( VREG_7_10 ) : ( n12194 ) ;
assign n12196 =  ( n11949 ) ? ( VREG_7_11 ) : ( n12195 ) ;
assign n12197 =  ( n11948 ) ? ( VREG_7_12 ) : ( n12196 ) ;
assign n12198 =  ( n11947 ) ? ( VREG_7_13 ) : ( n12197 ) ;
assign n12199 =  ( n11946 ) ? ( VREG_7_14 ) : ( n12198 ) ;
assign n12200 =  ( n11945 ) ? ( VREG_7_15 ) : ( n12199 ) ;
assign n12201 =  ( n11944 ) ? ( VREG_8_0 ) : ( n12200 ) ;
assign n12202 =  ( n11943 ) ? ( VREG_8_1 ) : ( n12201 ) ;
assign n12203 =  ( n11942 ) ? ( VREG_8_2 ) : ( n12202 ) ;
assign n12204 =  ( n11941 ) ? ( VREG_8_3 ) : ( n12203 ) ;
assign n12205 =  ( n11940 ) ? ( VREG_8_4 ) : ( n12204 ) ;
assign n12206 =  ( n11939 ) ? ( VREG_8_5 ) : ( n12205 ) ;
assign n12207 =  ( n11938 ) ? ( VREG_8_6 ) : ( n12206 ) ;
assign n12208 =  ( n11937 ) ? ( VREG_8_7 ) : ( n12207 ) ;
assign n12209 =  ( n11936 ) ? ( VREG_8_8 ) : ( n12208 ) ;
assign n12210 =  ( n11935 ) ? ( VREG_8_9 ) : ( n12209 ) ;
assign n12211 =  ( n11934 ) ? ( VREG_8_10 ) : ( n12210 ) ;
assign n12212 =  ( n11933 ) ? ( VREG_8_11 ) : ( n12211 ) ;
assign n12213 =  ( n11932 ) ? ( VREG_8_12 ) : ( n12212 ) ;
assign n12214 =  ( n11931 ) ? ( VREG_8_13 ) : ( n12213 ) ;
assign n12215 =  ( n11930 ) ? ( VREG_8_14 ) : ( n12214 ) ;
assign n12216 =  ( n11929 ) ? ( VREG_8_15 ) : ( n12215 ) ;
assign n12217 =  ( n11928 ) ? ( VREG_9_0 ) : ( n12216 ) ;
assign n12218 =  ( n11927 ) ? ( VREG_9_1 ) : ( n12217 ) ;
assign n12219 =  ( n11926 ) ? ( VREG_9_2 ) : ( n12218 ) ;
assign n12220 =  ( n11925 ) ? ( VREG_9_3 ) : ( n12219 ) ;
assign n12221 =  ( n11924 ) ? ( VREG_9_4 ) : ( n12220 ) ;
assign n12222 =  ( n11923 ) ? ( VREG_9_5 ) : ( n12221 ) ;
assign n12223 =  ( n11922 ) ? ( VREG_9_6 ) : ( n12222 ) ;
assign n12224 =  ( n11921 ) ? ( VREG_9_7 ) : ( n12223 ) ;
assign n12225 =  ( n11920 ) ? ( VREG_9_8 ) : ( n12224 ) ;
assign n12226 =  ( n11919 ) ? ( VREG_9_9 ) : ( n12225 ) ;
assign n12227 =  ( n11918 ) ? ( VREG_9_10 ) : ( n12226 ) ;
assign n12228 =  ( n11917 ) ? ( VREG_9_11 ) : ( n12227 ) ;
assign n12229 =  ( n11916 ) ? ( VREG_9_12 ) : ( n12228 ) ;
assign n12230 =  ( n11915 ) ? ( VREG_9_13 ) : ( n12229 ) ;
assign n12231 =  ( n11914 ) ? ( VREG_9_14 ) : ( n12230 ) ;
assign n12232 =  ( n11913 ) ? ( VREG_9_15 ) : ( n12231 ) ;
assign n12233 =  ( n11912 ) ? ( VREG_10_0 ) : ( n12232 ) ;
assign n12234 =  ( n11911 ) ? ( VREG_10_1 ) : ( n12233 ) ;
assign n12235 =  ( n11910 ) ? ( VREG_10_2 ) : ( n12234 ) ;
assign n12236 =  ( n11909 ) ? ( VREG_10_3 ) : ( n12235 ) ;
assign n12237 =  ( n11908 ) ? ( VREG_10_4 ) : ( n12236 ) ;
assign n12238 =  ( n11907 ) ? ( VREG_10_5 ) : ( n12237 ) ;
assign n12239 =  ( n11906 ) ? ( VREG_10_6 ) : ( n12238 ) ;
assign n12240 =  ( n11905 ) ? ( VREG_10_7 ) : ( n12239 ) ;
assign n12241 =  ( n11904 ) ? ( VREG_10_8 ) : ( n12240 ) ;
assign n12242 =  ( n11903 ) ? ( VREG_10_9 ) : ( n12241 ) ;
assign n12243 =  ( n11902 ) ? ( VREG_10_10 ) : ( n12242 ) ;
assign n12244 =  ( n11901 ) ? ( VREG_10_11 ) : ( n12243 ) ;
assign n12245 =  ( n11900 ) ? ( VREG_10_12 ) : ( n12244 ) ;
assign n12246 =  ( n11899 ) ? ( VREG_10_13 ) : ( n12245 ) ;
assign n12247 =  ( n11898 ) ? ( VREG_10_14 ) : ( n12246 ) ;
assign n12248 =  ( n11897 ) ? ( VREG_10_15 ) : ( n12247 ) ;
assign n12249 =  ( n11896 ) ? ( VREG_11_0 ) : ( n12248 ) ;
assign n12250 =  ( n11895 ) ? ( VREG_11_1 ) : ( n12249 ) ;
assign n12251 =  ( n11894 ) ? ( VREG_11_2 ) : ( n12250 ) ;
assign n12252 =  ( n11893 ) ? ( VREG_11_3 ) : ( n12251 ) ;
assign n12253 =  ( n11892 ) ? ( VREG_11_4 ) : ( n12252 ) ;
assign n12254 =  ( n11891 ) ? ( VREG_11_5 ) : ( n12253 ) ;
assign n12255 =  ( n11890 ) ? ( VREG_11_6 ) : ( n12254 ) ;
assign n12256 =  ( n11889 ) ? ( VREG_11_7 ) : ( n12255 ) ;
assign n12257 =  ( n11888 ) ? ( VREG_11_8 ) : ( n12256 ) ;
assign n12258 =  ( n11887 ) ? ( VREG_11_9 ) : ( n12257 ) ;
assign n12259 =  ( n11886 ) ? ( VREG_11_10 ) : ( n12258 ) ;
assign n12260 =  ( n11885 ) ? ( VREG_11_11 ) : ( n12259 ) ;
assign n12261 =  ( n11884 ) ? ( VREG_11_12 ) : ( n12260 ) ;
assign n12262 =  ( n11883 ) ? ( VREG_11_13 ) : ( n12261 ) ;
assign n12263 =  ( n11882 ) ? ( VREG_11_14 ) : ( n12262 ) ;
assign n12264 =  ( n11881 ) ? ( VREG_11_15 ) : ( n12263 ) ;
assign n12265 =  ( n11880 ) ? ( VREG_12_0 ) : ( n12264 ) ;
assign n12266 =  ( n11879 ) ? ( VREG_12_1 ) : ( n12265 ) ;
assign n12267 =  ( n11878 ) ? ( VREG_12_2 ) : ( n12266 ) ;
assign n12268 =  ( n11877 ) ? ( VREG_12_3 ) : ( n12267 ) ;
assign n12269 =  ( n11876 ) ? ( VREG_12_4 ) : ( n12268 ) ;
assign n12270 =  ( n11875 ) ? ( VREG_12_5 ) : ( n12269 ) ;
assign n12271 =  ( n11874 ) ? ( VREG_12_6 ) : ( n12270 ) ;
assign n12272 =  ( n11873 ) ? ( VREG_12_7 ) : ( n12271 ) ;
assign n12273 =  ( n11872 ) ? ( VREG_12_8 ) : ( n12272 ) ;
assign n12274 =  ( n11871 ) ? ( VREG_12_9 ) : ( n12273 ) ;
assign n12275 =  ( n11870 ) ? ( VREG_12_10 ) : ( n12274 ) ;
assign n12276 =  ( n11869 ) ? ( VREG_12_11 ) : ( n12275 ) ;
assign n12277 =  ( n11868 ) ? ( VREG_12_12 ) : ( n12276 ) ;
assign n12278 =  ( n11867 ) ? ( VREG_12_13 ) : ( n12277 ) ;
assign n12279 =  ( n11866 ) ? ( VREG_12_14 ) : ( n12278 ) ;
assign n12280 =  ( n11865 ) ? ( VREG_12_15 ) : ( n12279 ) ;
assign n12281 =  ( n11864 ) ? ( VREG_13_0 ) : ( n12280 ) ;
assign n12282 =  ( n11863 ) ? ( VREG_13_1 ) : ( n12281 ) ;
assign n12283 =  ( n11862 ) ? ( VREG_13_2 ) : ( n12282 ) ;
assign n12284 =  ( n11861 ) ? ( VREG_13_3 ) : ( n12283 ) ;
assign n12285 =  ( n11860 ) ? ( VREG_13_4 ) : ( n12284 ) ;
assign n12286 =  ( n11859 ) ? ( VREG_13_5 ) : ( n12285 ) ;
assign n12287 =  ( n11858 ) ? ( VREG_13_6 ) : ( n12286 ) ;
assign n12288 =  ( n11857 ) ? ( VREG_13_7 ) : ( n12287 ) ;
assign n12289 =  ( n11856 ) ? ( VREG_13_8 ) : ( n12288 ) ;
assign n12290 =  ( n11855 ) ? ( VREG_13_9 ) : ( n12289 ) ;
assign n12291 =  ( n11854 ) ? ( VREG_13_10 ) : ( n12290 ) ;
assign n12292 =  ( n11853 ) ? ( VREG_13_11 ) : ( n12291 ) ;
assign n12293 =  ( n11852 ) ? ( VREG_13_12 ) : ( n12292 ) ;
assign n12294 =  ( n11851 ) ? ( VREG_13_13 ) : ( n12293 ) ;
assign n12295 =  ( n11850 ) ? ( VREG_13_14 ) : ( n12294 ) ;
assign n12296 =  ( n11849 ) ? ( VREG_13_15 ) : ( n12295 ) ;
assign n12297 =  ( n11848 ) ? ( VREG_14_0 ) : ( n12296 ) ;
assign n12298 =  ( n11847 ) ? ( VREG_14_1 ) : ( n12297 ) ;
assign n12299 =  ( n11846 ) ? ( VREG_14_2 ) : ( n12298 ) ;
assign n12300 =  ( n11845 ) ? ( VREG_14_3 ) : ( n12299 ) ;
assign n12301 =  ( n11844 ) ? ( VREG_14_4 ) : ( n12300 ) ;
assign n12302 =  ( n11843 ) ? ( VREG_14_5 ) : ( n12301 ) ;
assign n12303 =  ( n11842 ) ? ( VREG_14_6 ) : ( n12302 ) ;
assign n12304 =  ( n11841 ) ? ( VREG_14_7 ) : ( n12303 ) ;
assign n12305 =  ( n11840 ) ? ( VREG_14_8 ) : ( n12304 ) ;
assign n12306 =  ( n11839 ) ? ( VREG_14_9 ) : ( n12305 ) ;
assign n12307 =  ( n11838 ) ? ( VREG_14_10 ) : ( n12306 ) ;
assign n12308 =  ( n11837 ) ? ( VREG_14_11 ) : ( n12307 ) ;
assign n12309 =  ( n11836 ) ? ( VREG_14_12 ) : ( n12308 ) ;
assign n12310 =  ( n11835 ) ? ( VREG_14_13 ) : ( n12309 ) ;
assign n12311 =  ( n11834 ) ? ( VREG_14_14 ) : ( n12310 ) ;
assign n12312 =  ( n11833 ) ? ( VREG_14_15 ) : ( n12311 ) ;
assign n12313 =  ( n11832 ) ? ( VREG_15_0 ) : ( n12312 ) ;
assign n12314 =  ( n11831 ) ? ( VREG_15_1 ) : ( n12313 ) ;
assign n12315 =  ( n11830 ) ? ( VREG_15_2 ) : ( n12314 ) ;
assign n12316 =  ( n11829 ) ? ( VREG_15_3 ) : ( n12315 ) ;
assign n12317 =  ( n11828 ) ? ( VREG_15_4 ) : ( n12316 ) ;
assign n12318 =  ( n11827 ) ? ( VREG_15_5 ) : ( n12317 ) ;
assign n12319 =  ( n11826 ) ? ( VREG_15_6 ) : ( n12318 ) ;
assign n12320 =  ( n11825 ) ? ( VREG_15_7 ) : ( n12319 ) ;
assign n12321 =  ( n11824 ) ? ( VREG_15_8 ) : ( n12320 ) ;
assign n12322 =  ( n11823 ) ? ( VREG_15_9 ) : ( n12321 ) ;
assign n12323 =  ( n11822 ) ? ( VREG_15_10 ) : ( n12322 ) ;
assign n12324 =  ( n11821 ) ? ( VREG_15_11 ) : ( n12323 ) ;
assign n12325 =  ( n11820 ) ? ( VREG_15_12 ) : ( n12324 ) ;
assign n12326 =  ( n11819 ) ? ( VREG_15_13 ) : ( n12325 ) ;
assign n12327 =  ( n11818 ) ? ( VREG_15_14 ) : ( n12326 ) ;
assign n12328 =  ( n11817 ) ? ( VREG_15_15 ) : ( n12327 ) ;
assign n12329 =  ( n11816 ) ? ( VREG_16_0 ) : ( n12328 ) ;
assign n12330 =  ( n11815 ) ? ( VREG_16_1 ) : ( n12329 ) ;
assign n12331 =  ( n11814 ) ? ( VREG_16_2 ) : ( n12330 ) ;
assign n12332 =  ( n11813 ) ? ( VREG_16_3 ) : ( n12331 ) ;
assign n12333 =  ( n11812 ) ? ( VREG_16_4 ) : ( n12332 ) ;
assign n12334 =  ( n11811 ) ? ( VREG_16_5 ) : ( n12333 ) ;
assign n12335 =  ( n11810 ) ? ( VREG_16_6 ) : ( n12334 ) ;
assign n12336 =  ( n11809 ) ? ( VREG_16_7 ) : ( n12335 ) ;
assign n12337 =  ( n11808 ) ? ( VREG_16_8 ) : ( n12336 ) ;
assign n12338 =  ( n11807 ) ? ( VREG_16_9 ) : ( n12337 ) ;
assign n12339 =  ( n11806 ) ? ( VREG_16_10 ) : ( n12338 ) ;
assign n12340 =  ( n11805 ) ? ( VREG_16_11 ) : ( n12339 ) ;
assign n12341 =  ( n11804 ) ? ( VREG_16_12 ) : ( n12340 ) ;
assign n12342 =  ( n11803 ) ? ( VREG_16_13 ) : ( n12341 ) ;
assign n12343 =  ( n11802 ) ? ( VREG_16_14 ) : ( n12342 ) ;
assign n12344 =  ( n11801 ) ? ( VREG_16_15 ) : ( n12343 ) ;
assign n12345 =  ( n11800 ) ? ( VREG_17_0 ) : ( n12344 ) ;
assign n12346 =  ( n11799 ) ? ( VREG_17_1 ) : ( n12345 ) ;
assign n12347 =  ( n11798 ) ? ( VREG_17_2 ) : ( n12346 ) ;
assign n12348 =  ( n11797 ) ? ( VREG_17_3 ) : ( n12347 ) ;
assign n12349 =  ( n11796 ) ? ( VREG_17_4 ) : ( n12348 ) ;
assign n12350 =  ( n11795 ) ? ( VREG_17_5 ) : ( n12349 ) ;
assign n12351 =  ( n11794 ) ? ( VREG_17_6 ) : ( n12350 ) ;
assign n12352 =  ( n11793 ) ? ( VREG_17_7 ) : ( n12351 ) ;
assign n12353 =  ( n11792 ) ? ( VREG_17_8 ) : ( n12352 ) ;
assign n12354 =  ( n11791 ) ? ( VREG_17_9 ) : ( n12353 ) ;
assign n12355 =  ( n11790 ) ? ( VREG_17_10 ) : ( n12354 ) ;
assign n12356 =  ( n11789 ) ? ( VREG_17_11 ) : ( n12355 ) ;
assign n12357 =  ( n11788 ) ? ( VREG_17_12 ) : ( n12356 ) ;
assign n12358 =  ( n11787 ) ? ( VREG_17_13 ) : ( n12357 ) ;
assign n12359 =  ( n11786 ) ? ( VREG_17_14 ) : ( n12358 ) ;
assign n12360 =  ( n11785 ) ? ( VREG_17_15 ) : ( n12359 ) ;
assign n12361 =  ( n11784 ) ? ( VREG_18_0 ) : ( n12360 ) ;
assign n12362 =  ( n11783 ) ? ( VREG_18_1 ) : ( n12361 ) ;
assign n12363 =  ( n11782 ) ? ( VREG_18_2 ) : ( n12362 ) ;
assign n12364 =  ( n11781 ) ? ( VREG_18_3 ) : ( n12363 ) ;
assign n12365 =  ( n11780 ) ? ( VREG_18_4 ) : ( n12364 ) ;
assign n12366 =  ( n11779 ) ? ( VREG_18_5 ) : ( n12365 ) ;
assign n12367 =  ( n11778 ) ? ( VREG_18_6 ) : ( n12366 ) ;
assign n12368 =  ( n11777 ) ? ( VREG_18_7 ) : ( n12367 ) ;
assign n12369 =  ( n11776 ) ? ( VREG_18_8 ) : ( n12368 ) ;
assign n12370 =  ( n11775 ) ? ( VREG_18_9 ) : ( n12369 ) ;
assign n12371 =  ( n11774 ) ? ( VREG_18_10 ) : ( n12370 ) ;
assign n12372 =  ( n11773 ) ? ( VREG_18_11 ) : ( n12371 ) ;
assign n12373 =  ( n11772 ) ? ( VREG_18_12 ) : ( n12372 ) ;
assign n12374 =  ( n11771 ) ? ( VREG_18_13 ) : ( n12373 ) ;
assign n12375 =  ( n11770 ) ? ( VREG_18_14 ) : ( n12374 ) ;
assign n12376 =  ( n11769 ) ? ( VREG_18_15 ) : ( n12375 ) ;
assign n12377 =  ( n11768 ) ? ( VREG_19_0 ) : ( n12376 ) ;
assign n12378 =  ( n11767 ) ? ( VREG_19_1 ) : ( n12377 ) ;
assign n12379 =  ( n11766 ) ? ( VREG_19_2 ) : ( n12378 ) ;
assign n12380 =  ( n11765 ) ? ( VREG_19_3 ) : ( n12379 ) ;
assign n12381 =  ( n11764 ) ? ( VREG_19_4 ) : ( n12380 ) ;
assign n12382 =  ( n11763 ) ? ( VREG_19_5 ) : ( n12381 ) ;
assign n12383 =  ( n11762 ) ? ( VREG_19_6 ) : ( n12382 ) ;
assign n12384 =  ( n11761 ) ? ( VREG_19_7 ) : ( n12383 ) ;
assign n12385 =  ( n11760 ) ? ( VREG_19_8 ) : ( n12384 ) ;
assign n12386 =  ( n11759 ) ? ( VREG_19_9 ) : ( n12385 ) ;
assign n12387 =  ( n11758 ) ? ( VREG_19_10 ) : ( n12386 ) ;
assign n12388 =  ( n11757 ) ? ( VREG_19_11 ) : ( n12387 ) ;
assign n12389 =  ( n11756 ) ? ( VREG_19_12 ) : ( n12388 ) ;
assign n12390 =  ( n11755 ) ? ( VREG_19_13 ) : ( n12389 ) ;
assign n12391 =  ( n11754 ) ? ( VREG_19_14 ) : ( n12390 ) ;
assign n12392 =  ( n11753 ) ? ( VREG_19_15 ) : ( n12391 ) ;
assign n12393 =  ( n11752 ) ? ( VREG_20_0 ) : ( n12392 ) ;
assign n12394 =  ( n11751 ) ? ( VREG_20_1 ) : ( n12393 ) ;
assign n12395 =  ( n11750 ) ? ( VREG_20_2 ) : ( n12394 ) ;
assign n12396 =  ( n11749 ) ? ( VREG_20_3 ) : ( n12395 ) ;
assign n12397 =  ( n11748 ) ? ( VREG_20_4 ) : ( n12396 ) ;
assign n12398 =  ( n11747 ) ? ( VREG_20_5 ) : ( n12397 ) ;
assign n12399 =  ( n11746 ) ? ( VREG_20_6 ) : ( n12398 ) ;
assign n12400 =  ( n11745 ) ? ( VREG_20_7 ) : ( n12399 ) ;
assign n12401 =  ( n11744 ) ? ( VREG_20_8 ) : ( n12400 ) ;
assign n12402 =  ( n11743 ) ? ( VREG_20_9 ) : ( n12401 ) ;
assign n12403 =  ( n11742 ) ? ( VREG_20_10 ) : ( n12402 ) ;
assign n12404 =  ( n11741 ) ? ( VREG_20_11 ) : ( n12403 ) ;
assign n12405 =  ( n11740 ) ? ( VREG_20_12 ) : ( n12404 ) ;
assign n12406 =  ( n11739 ) ? ( VREG_20_13 ) : ( n12405 ) ;
assign n12407 =  ( n11738 ) ? ( VREG_20_14 ) : ( n12406 ) ;
assign n12408 =  ( n11737 ) ? ( VREG_20_15 ) : ( n12407 ) ;
assign n12409 =  ( n11736 ) ? ( VREG_21_0 ) : ( n12408 ) ;
assign n12410 =  ( n11735 ) ? ( VREG_21_1 ) : ( n12409 ) ;
assign n12411 =  ( n11734 ) ? ( VREG_21_2 ) : ( n12410 ) ;
assign n12412 =  ( n11733 ) ? ( VREG_21_3 ) : ( n12411 ) ;
assign n12413 =  ( n11732 ) ? ( VREG_21_4 ) : ( n12412 ) ;
assign n12414 =  ( n11731 ) ? ( VREG_21_5 ) : ( n12413 ) ;
assign n12415 =  ( n11730 ) ? ( VREG_21_6 ) : ( n12414 ) ;
assign n12416 =  ( n11729 ) ? ( VREG_21_7 ) : ( n12415 ) ;
assign n12417 =  ( n11728 ) ? ( VREG_21_8 ) : ( n12416 ) ;
assign n12418 =  ( n11727 ) ? ( VREG_21_9 ) : ( n12417 ) ;
assign n12419 =  ( n11726 ) ? ( VREG_21_10 ) : ( n12418 ) ;
assign n12420 =  ( n11725 ) ? ( VREG_21_11 ) : ( n12419 ) ;
assign n12421 =  ( n11724 ) ? ( VREG_21_12 ) : ( n12420 ) ;
assign n12422 =  ( n11723 ) ? ( VREG_21_13 ) : ( n12421 ) ;
assign n12423 =  ( n11722 ) ? ( VREG_21_14 ) : ( n12422 ) ;
assign n12424 =  ( n11721 ) ? ( VREG_21_15 ) : ( n12423 ) ;
assign n12425 =  ( n11720 ) ? ( VREG_22_0 ) : ( n12424 ) ;
assign n12426 =  ( n11719 ) ? ( VREG_22_1 ) : ( n12425 ) ;
assign n12427 =  ( n11718 ) ? ( VREG_22_2 ) : ( n12426 ) ;
assign n12428 =  ( n11717 ) ? ( VREG_22_3 ) : ( n12427 ) ;
assign n12429 =  ( n11716 ) ? ( VREG_22_4 ) : ( n12428 ) ;
assign n12430 =  ( n11715 ) ? ( VREG_22_5 ) : ( n12429 ) ;
assign n12431 =  ( n11714 ) ? ( VREG_22_6 ) : ( n12430 ) ;
assign n12432 =  ( n11713 ) ? ( VREG_22_7 ) : ( n12431 ) ;
assign n12433 =  ( n11712 ) ? ( VREG_22_8 ) : ( n12432 ) ;
assign n12434 =  ( n11711 ) ? ( VREG_22_9 ) : ( n12433 ) ;
assign n12435 =  ( n11710 ) ? ( VREG_22_10 ) : ( n12434 ) ;
assign n12436 =  ( n11709 ) ? ( VREG_22_11 ) : ( n12435 ) ;
assign n12437 =  ( n11708 ) ? ( VREG_22_12 ) : ( n12436 ) ;
assign n12438 =  ( n11707 ) ? ( VREG_22_13 ) : ( n12437 ) ;
assign n12439 =  ( n11706 ) ? ( VREG_22_14 ) : ( n12438 ) ;
assign n12440 =  ( n11705 ) ? ( VREG_22_15 ) : ( n12439 ) ;
assign n12441 =  ( n11704 ) ? ( VREG_23_0 ) : ( n12440 ) ;
assign n12442 =  ( n11703 ) ? ( VREG_23_1 ) : ( n12441 ) ;
assign n12443 =  ( n11702 ) ? ( VREG_23_2 ) : ( n12442 ) ;
assign n12444 =  ( n11701 ) ? ( VREG_23_3 ) : ( n12443 ) ;
assign n12445 =  ( n11700 ) ? ( VREG_23_4 ) : ( n12444 ) ;
assign n12446 =  ( n11699 ) ? ( VREG_23_5 ) : ( n12445 ) ;
assign n12447 =  ( n11698 ) ? ( VREG_23_6 ) : ( n12446 ) ;
assign n12448 =  ( n11697 ) ? ( VREG_23_7 ) : ( n12447 ) ;
assign n12449 =  ( n11696 ) ? ( VREG_23_8 ) : ( n12448 ) ;
assign n12450 =  ( n11695 ) ? ( VREG_23_9 ) : ( n12449 ) ;
assign n12451 =  ( n11694 ) ? ( VREG_23_10 ) : ( n12450 ) ;
assign n12452 =  ( n11693 ) ? ( VREG_23_11 ) : ( n12451 ) ;
assign n12453 =  ( n11692 ) ? ( VREG_23_12 ) : ( n12452 ) ;
assign n12454 =  ( n11691 ) ? ( VREG_23_13 ) : ( n12453 ) ;
assign n12455 =  ( n11690 ) ? ( VREG_23_14 ) : ( n12454 ) ;
assign n12456 =  ( n11689 ) ? ( VREG_23_15 ) : ( n12455 ) ;
assign n12457 =  ( n11688 ) ? ( VREG_24_0 ) : ( n12456 ) ;
assign n12458 =  ( n11687 ) ? ( VREG_24_1 ) : ( n12457 ) ;
assign n12459 =  ( n11686 ) ? ( VREG_24_2 ) : ( n12458 ) ;
assign n12460 =  ( n11685 ) ? ( VREG_24_3 ) : ( n12459 ) ;
assign n12461 =  ( n11684 ) ? ( VREG_24_4 ) : ( n12460 ) ;
assign n12462 =  ( n11683 ) ? ( VREG_24_5 ) : ( n12461 ) ;
assign n12463 =  ( n11682 ) ? ( VREG_24_6 ) : ( n12462 ) ;
assign n12464 =  ( n11681 ) ? ( VREG_24_7 ) : ( n12463 ) ;
assign n12465 =  ( n11680 ) ? ( VREG_24_8 ) : ( n12464 ) ;
assign n12466 =  ( n11679 ) ? ( VREG_24_9 ) : ( n12465 ) ;
assign n12467 =  ( n11678 ) ? ( VREG_24_10 ) : ( n12466 ) ;
assign n12468 =  ( n11677 ) ? ( VREG_24_11 ) : ( n12467 ) ;
assign n12469 =  ( n11676 ) ? ( VREG_24_12 ) : ( n12468 ) ;
assign n12470 =  ( n11675 ) ? ( VREG_24_13 ) : ( n12469 ) ;
assign n12471 =  ( n11674 ) ? ( VREG_24_14 ) : ( n12470 ) ;
assign n12472 =  ( n11673 ) ? ( VREG_24_15 ) : ( n12471 ) ;
assign n12473 =  ( n11672 ) ? ( VREG_25_0 ) : ( n12472 ) ;
assign n12474 =  ( n11671 ) ? ( VREG_25_1 ) : ( n12473 ) ;
assign n12475 =  ( n11670 ) ? ( VREG_25_2 ) : ( n12474 ) ;
assign n12476 =  ( n11669 ) ? ( VREG_25_3 ) : ( n12475 ) ;
assign n12477 =  ( n11668 ) ? ( VREG_25_4 ) : ( n12476 ) ;
assign n12478 =  ( n11667 ) ? ( VREG_25_5 ) : ( n12477 ) ;
assign n12479 =  ( n11666 ) ? ( VREG_25_6 ) : ( n12478 ) ;
assign n12480 =  ( n11665 ) ? ( VREG_25_7 ) : ( n12479 ) ;
assign n12481 =  ( n11664 ) ? ( VREG_25_8 ) : ( n12480 ) ;
assign n12482 =  ( n11663 ) ? ( VREG_25_9 ) : ( n12481 ) ;
assign n12483 =  ( n11662 ) ? ( VREG_25_10 ) : ( n12482 ) ;
assign n12484 =  ( n11661 ) ? ( VREG_25_11 ) : ( n12483 ) ;
assign n12485 =  ( n11660 ) ? ( VREG_25_12 ) : ( n12484 ) ;
assign n12486 =  ( n11659 ) ? ( VREG_25_13 ) : ( n12485 ) ;
assign n12487 =  ( n11658 ) ? ( VREG_25_14 ) : ( n12486 ) ;
assign n12488 =  ( n11657 ) ? ( VREG_25_15 ) : ( n12487 ) ;
assign n12489 =  ( n11656 ) ? ( VREG_26_0 ) : ( n12488 ) ;
assign n12490 =  ( n11655 ) ? ( VREG_26_1 ) : ( n12489 ) ;
assign n12491 =  ( n11654 ) ? ( VREG_26_2 ) : ( n12490 ) ;
assign n12492 =  ( n11653 ) ? ( VREG_26_3 ) : ( n12491 ) ;
assign n12493 =  ( n11652 ) ? ( VREG_26_4 ) : ( n12492 ) ;
assign n12494 =  ( n11651 ) ? ( VREG_26_5 ) : ( n12493 ) ;
assign n12495 =  ( n11650 ) ? ( VREG_26_6 ) : ( n12494 ) ;
assign n12496 =  ( n11649 ) ? ( VREG_26_7 ) : ( n12495 ) ;
assign n12497 =  ( n11648 ) ? ( VREG_26_8 ) : ( n12496 ) ;
assign n12498 =  ( n11647 ) ? ( VREG_26_9 ) : ( n12497 ) ;
assign n12499 =  ( n11646 ) ? ( VREG_26_10 ) : ( n12498 ) ;
assign n12500 =  ( n11645 ) ? ( VREG_26_11 ) : ( n12499 ) ;
assign n12501 =  ( n11644 ) ? ( VREG_26_12 ) : ( n12500 ) ;
assign n12502 =  ( n11643 ) ? ( VREG_26_13 ) : ( n12501 ) ;
assign n12503 =  ( n11642 ) ? ( VREG_26_14 ) : ( n12502 ) ;
assign n12504 =  ( n11641 ) ? ( VREG_26_15 ) : ( n12503 ) ;
assign n12505 =  ( n11640 ) ? ( VREG_27_0 ) : ( n12504 ) ;
assign n12506 =  ( n11639 ) ? ( VREG_27_1 ) : ( n12505 ) ;
assign n12507 =  ( n11638 ) ? ( VREG_27_2 ) : ( n12506 ) ;
assign n12508 =  ( n11637 ) ? ( VREG_27_3 ) : ( n12507 ) ;
assign n12509 =  ( n11636 ) ? ( VREG_27_4 ) : ( n12508 ) ;
assign n12510 =  ( n11635 ) ? ( VREG_27_5 ) : ( n12509 ) ;
assign n12511 =  ( n11634 ) ? ( VREG_27_6 ) : ( n12510 ) ;
assign n12512 =  ( n11633 ) ? ( VREG_27_7 ) : ( n12511 ) ;
assign n12513 =  ( n11632 ) ? ( VREG_27_8 ) : ( n12512 ) ;
assign n12514 =  ( n11631 ) ? ( VREG_27_9 ) : ( n12513 ) ;
assign n12515 =  ( n11630 ) ? ( VREG_27_10 ) : ( n12514 ) ;
assign n12516 =  ( n11629 ) ? ( VREG_27_11 ) : ( n12515 ) ;
assign n12517 =  ( n11628 ) ? ( VREG_27_12 ) : ( n12516 ) ;
assign n12518 =  ( n11627 ) ? ( VREG_27_13 ) : ( n12517 ) ;
assign n12519 =  ( n11626 ) ? ( VREG_27_14 ) : ( n12518 ) ;
assign n12520 =  ( n11625 ) ? ( VREG_27_15 ) : ( n12519 ) ;
assign n12521 =  ( n11624 ) ? ( VREG_28_0 ) : ( n12520 ) ;
assign n12522 =  ( n11623 ) ? ( VREG_28_1 ) : ( n12521 ) ;
assign n12523 =  ( n11622 ) ? ( VREG_28_2 ) : ( n12522 ) ;
assign n12524 =  ( n11621 ) ? ( VREG_28_3 ) : ( n12523 ) ;
assign n12525 =  ( n11620 ) ? ( VREG_28_4 ) : ( n12524 ) ;
assign n12526 =  ( n11619 ) ? ( VREG_28_5 ) : ( n12525 ) ;
assign n12527 =  ( n11618 ) ? ( VREG_28_6 ) : ( n12526 ) ;
assign n12528 =  ( n11617 ) ? ( VREG_28_7 ) : ( n12527 ) ;
assign n12529 =  ( n11616 ) ? ( VREG_28_8 ) : ( n12528 ) ;
assign n12530 =  ( n11615 ) ? ( VREG_28_9 ) : ( n12529 ) ;
assign n12531 =  ( n11614 ) ? ( VREG_28_10 ) : ( n12530 ) ;
assign n12532 =  ( n11613 ) ? ( VREG_28_11 ) : ( n12531 ) ;
assign n12533 =  ( n11612 ) ? ( VREG_28_12 ) : ( n12532 ) ;
assign n12534 =  ( n11611 ) ? ( VREG_28_13 ) : ( n12533 ) ;
assign n12535 =  ( n11610 ) ? ( VREG_28_14 ) : ( n12534 ) ;
assign n12536 =  ( n11609 ) ? ( VREG_28_15 ) : ( n12535 ) ;
assign n12537 =  ( n11608 ) ? ( VREG_29_0 ) : ( n12536 ) ;
assign n12538 =  ( n11607 ) ? ( VREG_29_1 ) : ( n12537 ) ;
assign n12539 =  ( n11606 ) ? ( VREG_29_2 ) : ( n12538 ) ;
assign n12540 =  ( n11605 ) ? ( VREG_29_3 ) : ( n12539 ) ;
assign n12541 =  ( n11604 ) ? ( VREG_29_4 ) : ( n12540 ) ;
assign n12542 =  ( n11603 ) ? ( VREG_29_5 ) : ( n12541 ) ;
assign n12543 =  ( n11602 ) ? ( VREG_29_6 ) : ( n12542 ) ;
assign n12544 =  ( n11601 ) ? ( VREG_29_7 ) : ( n12543 ) ;
assign n12545 =  ( n11600 ) ? ( VREG_29_8 ) : ( n12544 ) ;
assign n12546 =  ( n11599 ) ? ( VREG_29_9 ) : ( n12545 ) ;
assign n12547 =  ( n11598 ) ? ( VREG_29_10 ) : ( n12546 ) ;
assign n12548 =  ( n11597 ) ? ( VREG_29_11 ) : ( n12547 ) ;
assign n12549 =  ( n11596 ) ? ( VREG_29_12 ) : ( n12548 ) ;
assign n12550 =  ( n11595 ) ? ( VREG_29_13 ) : ( n12549 ) ;
assign n12551 =  ( n11594 ) ? ( VREG_29_14 ) : ( n12550 ) ;
assign n12552 =  ( n11593 ) ? ( VREG_29_15 ) : ( n12551 ) ;
assign n12553 =  ( n11592 ) ? ( VREG_30_0 ) : ( n12552 ) ;
assign n12554 =  ( n11591 ) ? ( VREG_30_1 ) : ( n12553 ) ;
assign n12555 =  ( n11590 ) ? ( VREG_30_2 ) : ( n12554 ) ;
assign n12556 =  ( n11589 ) ? ( VREG_30_3 ) : ( n12555 ) ;
assign n12557 =  ( n11588 ) ? ( VREG_30_4 ) : ( n12556 ) ;
assign n12558 =  ( n11587 ) ? ( VREG_30_5 ) : ( n12557 ) ;
assign n12559 =  ( n11586 ) ? ( VREG_30_6 ) : ( n12558 ) ;
assign n12560 =  ( n11585 ) ? ( VREG_30_7 ) : ( n12559 ) ;
assign n12561 =  ( n11584 ) ? ( VREG_30_8 ) : ( n12560 ) ;
assign n12562 =  ( n11583 ) ? ( VREG_30_9 ) : ( n12561 ) ;
assign n12563 =  ( n11582 ) ? ( VREG_30_10 ) : ( n12562 ) ;
assign n12564 =  ( n11581 ) ? ( VREG_30_11 ) : ( n12563 ) ;
assign n12565 =  ( n11580 ) ? ( VREG_30_12 ) : ( n12564 ) ;
assign n12566 =  ( n11579 ) ? ( VREG_30_13 ) : ( n12565 ) ;
assign n12567 =  ( n11578 ) ? ( VREG_30_14 ) : ( n12566 ) ;
assign n12568 =  ( n11577 ) ? ( VREG_30_15 ) : ( n12567 ) ;
assign n12569 =  ( n11576 ) ? ( VREG_31_0 ) : ( n12568 ) ;
assign n12570 =  ( n11574 ) ? ( VREG_31_1 ) : ( n12569 ) ;
assign n12571 =  ( n11572 ) ? ( VREG_31_2 ) : ( n12570 ) ;
assign n12572 =  ( n11570 ) ? ( VREG_31_3 ) : ( n12571 ) ;
assign n12573 =  ( n11568 ) ? ( VREG_31_4 ) : ( n12572 ) ;
assign n12574 =  ( n11566 ) ? ( VREG_31_5 ) : ( n12573 ) ;
assign n12575 =  ( n11564 ) ? ( VREG_31_6 ) : ( n12574 ) ;
assign n12576 =  ( n11562 ) ? ( VREG_31_7 ) : ( n12575 ) ;
assign n12577 =  ( n11560 ) ? ( VREG_31_8 ) : ( n12576 ) ;
assign n12578 =  ( n11558 ) ? ( VREG_31_9 ) : ( n12577 ) ;
assign n12579 =  ( n11556 ) ? ( VREG_31_10 ) : ( n12578 ) ;
assign n12580 =  ( n11554 ) ? ( VREG_31_11 ) : ( n12579 ) ;
assign n12581 =  ( n11552 ) ? ( VREG_31_12 ) : ( n12580 ) ;
assign n12582 =  ( n11550 ) ? ( VREG_31_13 ) : ( n12581 ) ;
assign n12583 =  ( n11548 ) ? ( VREG_31_14 ) : ( n12582 ) ;
assign n12584 =  ( n11546 ) ? ( VREG_31_15 ) : ( n12583 ) ;
assign n12585 =  ( n12584 ) + ( n140 )  ;
assign n12586 =  ( n12584 ) - ( n140 )  ;
assign n12587 =  ( n12584 ) & ( n140 )  ;
assign n12588 =  ( n12584 ) | ( n140 )  ;
assign n12589 =  ( ( n12584 ) * ( n140 ))  ;
assign n12590 =  ( n148 ) ? ( n12589 ) : ( VREG_0_13 ) ;
assign n12591 =  ( n146 ) ? ( n12588 ) : ( n12590 ) ;
assign n12592 =  ( n144 ) ? ( n12587 ) : ( n12591 ) ;
assign n12593 =  ( n142 ) ? ( n12586 ) : ( n12592 ) ;
assign n12594 =  ( n10 ) ? ( n12585 ) : ( n12593 ) ;
assign n12595 =  ( n77 ) & ( n11545 )  ;
assign n12596 =  ( n77 ) & ( n11547 )  ;
assign n12597 =  ( n77 ) & ( n11549 )  ;
assign n12598 =  ( n77 ) & ( n11551 )  ;
assign n12599 =  ( n77 ) & ( n11553 )  ;
assign n12600 =  ( n77 ) & ( n11555 )  ;
assign n12601 =  ( n77 ) & ( n11557 )  ;
assign n12602 =  ( n77 ) & ( n11559 )  ;
assign n12603 =  ( n77 ) & ( n11561 )  ;
assign n12604 =  ( n77 ) & ( n11563 )  ;
assign n12605 =  ( n77 ) & ( n11565 )  ;
assign n12606 =  ( n77 ) & ( n11567 )  ;
assign n12607 =  ( n77 ) & ( n11569 )  ;
assign n12608 =  ( n77 ) & ( n11571 )  ;
assign n12609 =  ( n77 ) & ( n11573 )  ;
assign n12610 =  ( n77 ) & ( n11575 )  ;
assign n12611 =  ( n78 ) & ( n11545 )  ;
assign n12612 =  ( n78 ) & ( n11547 )  ;
assign n12613 =  ( n78 ) & ( n11549 )  ;
assign n12614 =  ( n78 ) & ( n11551 )  ;
assign n12615 =  ( n78 ) & ( n11553 )  ;
assign n12616 =  ( n78 ) & ( n11555 )  ;
assign n12617 =  ( n78 ) & ( n11557 )  ;
assign n12618 =  ( n78 ) & ( n11559 )  ;
assign n12619 =  ( n78 ) & ( n11561 )  ;
assign n12620 =  ( n78 ) & ( n11563 )  ;
assign n12621 =  ( n78 ) & ( n11565 )  ;
assign n12622 =  ( n78 ) & ( n11567 )  ;
assign n12623 =  ( n78 ) & ( n11569 )  ;
assign n12624 =  ( n78 ) & ( n11571 )  ;
assign n12625 =  ( n78 ) & ( n11573 )  ;
assign n12626 =  ( n78 ) & ( n11575 )  ;
assign n12627 =  ( n79 ) & ( n11545 )  ;
assign n12628 =  ( n79 ) & ( n11547 )  ;
assign n12629 =  ( n79 ) & ( n11549 )  ;
assign n12630 =  ( n79 ) & ( n11551 )  ;
assign n12631 =  ( n79 ) & ( n11553 )  ;
assign n12632 =  ( n79 ) & ( n11555 )  ;
assign n12633 =  ( n79 ) & ( n11557 )  ;
assign n12634 =  ( n79 ) & ( n11559 )  ;
assign n12635 =  ( n79 ) & ( n11561 )  ;
assign n12636 =  ( n79 ) & ( n11563 )  ;
assign n12637 =  ( n79 ) & ( n11565 )  ;
assign n12638 =  ( n79 ) & ( n11567 )  ;
assign n12639 =  ( n79 ) & ( n11569 )  ;
assign n12640 =  ( n79 ) & ( n11571 )  ;
assign n12641 =  ( n79 ) & ( n11573 )  ;
assign n12642 =  ( n79 ) & ( n11575 )  ;
assign n12643 =  ( n80 ) & ( n11545 )  ;
assign n12644 =  ( n80 ) & ( n11547 )  ;
assign n12645 =  ( n80 ) & ( n11549 )  ;
assign n12646 =  ( n80 ) & ( n11551 )  ;
assign n12647 =  ( n80 ) & ( n11553 )  ;
assign n12648 =  ( n80 ) & ( n11555 )  ;
assign n12649 =  ( n80 ) & ( n11557 )  ;
assign n12650 =  ( n80 ) & ( n11559 )  ;
assign n12651 =  ( n80 ) & ( n11561 )  ;
assign n12652 =  ( n80 ) & ( n11563 )  ;
assign n12653 =  ( n80 ) & ( n11565 )  ;
assign n12654 =  ( n80 ) & ( n11567 )  ;
assign n12655 =  ( n80 ) & ( n11569 )  ;
assign n12656 =  ( n80 ) & ( n11571 )  ;
assign n12657 =  ( n80 ) & ( n11573 )  ;
assign n12658 =  ( n80 ) & ( n11575 )  ;
assign n12659 =  ( n81 ) & ( n11545 )  ;
assign n12660 =  ( n81 ) & ( n11547 )  ;
assign n12661 =  ( n81 ) & ( n11549 )  ;
assign n12662 =  ( n81 ) & ( n11551 )  ;
assign n12663 =  ( n81 ) & ( n11553 )  ;
assign n12664 =  ( n81 ) & ( n11555 )  ;
assign n12665 =  ( n81 ) & ( n11557 )  ;
assign n12666 =  ( n81 ) & ( n11559 )  ;
assign n12667 =  ( n81 ) & ( n11561 )  ;
assign n12668 =  ( n81 ) & ( n11563 )  ;
assign n12669 =  ( n81 ) & ( n11565 )  ;
assign n12670 =  ( n81 ) & ( n11567 )  ;
assign n12671 =  ( n81 ) & ( n11569 )  ;
assign n12672 =  ( n81 ) & ( n11571 )  ;
assign n12673 =  ( n81 ) & ( n11573 )  ;
assign n12674 =  ( n81 ) & ( n11575 )  ;
assign n12675 =  ( n82 ) & ( n11545 )  ;
assign n12676 =  ( n82 ) & ( n11547 )  ;
assign n12677 =  ( n82 ) & ( n11549 )  ;
assign n12678 =  ( n82 ) & ( n11551 )  ;
assign n12679 =  ( n82 ) & ( n11553 )  ;
assign n12680 =  ( n82 ) & ( n11555 )  ;
assign n12681 =  ( n82 ) & ( n11557 )  ;
assign n12682 =  ( n82 ) & ( n11559 )  ;
assign n12683 =  ( n82 ) & ( n11561 )  ;
assign n12684 =  ( n82 ) & ( n11563 )  ;
assign n12685 =  ( n82 ) & ( n11565 )  ;
assign n12686 =  ( n82 ) & ( n11567 )  ;
assign n12687 =  ( n82 ) & ( n11569 )  ;
assign n12688 =  ( n82 ) & ( n11571 )  ;
assign n12689 =  ( n82 ) & ( n11573 )  ;
assign n12690 =  ( n82 ) & ( n11575 )  ;
assign n12691 =  ( n83 ) & ( n11545 )  ;
assign n12692 =  ( n83 ) & ( n11547 )  ;
assign n12693 =  ( n83 ) & ( n11549 )  ;
assign n12694 =  ( n83 ) & ( n11551 )  ;
assign n12695 =  ( n83 ) & ( n11553 )  ;
assign n12696 =  ( n83 ) & ( n11555 )  ;
assign n12697 =  ( n83 ) & ( n11557 )  ;
assign n12698 =  ( n83 ) & ( n11559 )  ;
assign n12699 =  ( n83 ) & ( n11561 )  ;
assign n12700 =  ( n83 ) & ( n11563 )  ;
assign n12701 =  ( n83 ) & ( n11565 )  ;
assign n12702 =  ( n83 ) & ( n11567 )  ;
assign n12703 =  ( n83 ) & ( n11569 )  ;
assign n12704 =  ( n83 ) & ( n11571 )  ;
assign n12705 =  ( n83 ) & ( n11573 )  ;
assign n12706 =  ( n83 ) & ( n11575 )  ;
assign n12707 =  ( n84 ) & ( n11545 )  ;
assign n12708 =  ( n84 ) & ( n11547 )  ;
assign n12709 =  ( n84 ) & ( n11549 )  ;
assign n12710 =  ( n84 ) & ( n11551 )  ;
assign n12711 =  ( n84 ) & ( n11553 )  ;
assign n12712 =  ( n84 ) & ( n11555 )  ;
assign n12713 =  ( n84 ) & ( n11557 )  ;
assign n12714 =  ( n84 ) & ( n11559 )  ;
assign n12715 =  ( n84 ) & ( n11561 )  ;
assign n12716 =  ( n84 ) & ( n11563 )  ;
assign n12717 =  ( n84 ) & ( n11565 )  ;
assign n12718 =  ( n84 ) & ( n11567 )  ;
assign n12719 =  ( n84 ) & ( n11569 )  ;
assign n12720 =  ( n84 ) & ( n11571 )  ;
assign n12721 =  ( n84 ) & ( n11573 )  ;
assign n12722 =  ( n84 ) & ( n11575 )  ;
assign n12723 =  ( n85 ) & ( n11545 )  ;
assign n12724 =  ( n85 ) & ( n11547 )  ;
assign n12725 =  ( n85 ) & ( n11549 )  ;
assign n12726 =  ( n85 ) & ( n11551 )  ;
assign n12727 =  ( n85 ) & ( n11553 )  ;
assign n12728 =  ( n85 ) & ( n11555 )  ;
assign n12729 =  ( n85 ) & ( n11557 )  ;
assign n12730 =  ( n85 ) & ( n11559 )  ;
assign n12731 =  ( n85 ) & ( n11561 )  ;
assign n12732 =  ( n85 ) & ( n11563 )  ;
assign n12733 =  ( n85 ) & ( n11565 )  ;
assign n12734 =  ( n85 ) & ( n11567 )  ;
assign n12735 =  ( n85 ) & ( n11569 )  ;
assign n12736 =  ( n85 ) & ( n11571 )  ;
assign n12737 =  ( n85 ) & ( n11573 )  ;
assign n12738 =  ( n85 ) & ( n11575 )  ;
assign n12739 =  ( n86 ) & ( n11545 )  ;
assign n12740 =  ( n86 ) & ( n11547 )  ;
assign n12741 =  ( n86 ) & ( n11549 )  ;
assign n12742 =  ( n86 ) & ( n11551 )  ;
assign n12743 =  ( n86 ) & ( n11553 )  ;
assign n12744 =  ( n86 ) & ( n11555 )  ;
assign n12745 =  ( n86 ) & ( n11557 )  ;
assign n12746 =  ( n86 ) & ( n11559 )  ;
assign n12747 =  ( n86 ) & ( n11561 )  ;
assign n12748 =  ( n86 ) & ( n11563 )  ;
assign n12749 =  ( n86 ) & ( n11565 )  ;
assign n12750 =  ( n86 ) & ( n11567 )  ;
assign n12751 =  ( n86 ) & ( n11569 )  ;
assign n12752 =  ( n86 ) & ( n11571 )  ;
assign n12753 =  ( n86 ) & ( n11573 )  ;
assign n12754 =  ( n86 ) & ( n11575 )  ;
assign n12755 =  ( n87 ) & ( n11545 )  ;
assign n12756 =  ( n87 ) & ( n11547 )  ;
assign n12757 =  ( n87 ) & ( n11549 )  ;
assign n12758 =  ( n87 ) & ( n11551 )  ;
assign n12759 =  ( n87 ) & ( n11553 )  ;
assign n12760 =  ( n87 ) & ( n11555 )  ;
assign n12761 =  ( n87 ) & ( n11557 )  ;
assign n12762 =  ( n87 ) & ( n11559 )  ;
assign n12763 =  ( n87 ) & ( n11561 )  ;
assign n12764 =  ( n87 ) & ( n11563 )  ;
assign n12765 =  ( n87 ) & ( n11565 )  ;
assign n12766 =  ( n87 ) & ( n11567 )  ;
assign n12767 =  ( n87 ) & ( n11569 )  ;
assign n12768 =  ( n87 ) & ( n11571 )  ;
assign n12769 =  ( n87 ) & ( n11573 )  ;
assign n12770 =  ( n87 ) & ( n11575 )  ;
assign n12771 =  ( n88 ) & ( n11545 )  ;
assign n12772 =  ( n88 ) & ( n11547 )  ;
assign n12773 =  ( n88 ) & ( n11549 )  ;
assign n12774 =  ( n88 ) & ( n11551 )  ;
assign n12775 =  ( n88 ) & ( n11553 )  ;
assign n12776 =  ( n88 ) & ( n11555 )  ;
assign n12777 =  ( n88 ) & ( n11557 )  ;
assign n12778 =  ( n88 ) & ( n11559 )  ;
assign n12779 =  ( n88 ) & ( n11561 )  ;
assign n12780 =  ( n88 ) & ( n11563 )  ;
assign n12781 =  ( n88 ) & ( n11565 )  ;
assign n12782 =  ( n88 ) & ( n11567 )  ;
assign n12783 =  ( n88 ) & ( n11569 )  ;
assign n12784 =  ( n88 ) & ( n11571 )  ;
assign n12785 =  ( n88 ) & ( n11573 )  ;
assign n12786 =  ( n88 ) & ( n11575 )  ;
assign n12787 =  ( n89 ) & ( n11545 )  ;
assign n12788 =  ( n89 ) & ( n11547 )  ;
assign n12789 =  ( n89 ) & ( n11549 )  ;
assign n12790 =  ( n89 ) & ( n11551 )  ;
assign n12791 =  ( n89 ) & ( n11553 )  ;
assign n12792 =  ( n89 ) & ( n11555 )  ;
assign n12793 =  ( n89 ) & ( n11557 )  ;
assign n12794 =  ( n89 ) & ( n11559 )  ;
assign n12795 =  ( n89 ) & ( n11561 )  ;
assign n12796 =  ( n89 ) & ( n11563 )  ;
assign n12797 =  ( n89 ) & ( n11565 )  ;
assign n12798 =  ( n89 ) & ( n11567 )  ;
assign n12799 =  ( n89 ) & ( n11569 )  ;
assign n12800 =  ( n89 ) & ( n11571 )  ;
assign n12801 =  ( n89 ) & ( n11573 )  ;
assign n12802 =  ( n89 ) & ( n11575 )  ;
assign n12803 =  ( n90 ) & ( n11545 )  ;
assign n12804 =  ( n90 ) & ( n11547 )  ;
assign n12805 =  ( n90 ) & ( n11549 )  ;
assign n12806 =  ( n90 ) & ( n11551 )  ;
assign n12807 =  ( n90 ) & ( n11553 )  ;
assign n12808 =  ( n90 ) & ( n11555 )  ;
assign n12809 =  ( n90 ) & ( n11557 )  ;
assign n12810 =  ( n90 ) & ( n11559 )  ;
assign n12811 =  ( n90 ) & ( n11561 )  ;
assign n12812 =  ( n90 ) & ( n11563 )  ;
assign n12813 =  ( n90 ) & ( n11565 )  ;
assign n12814 =  ( n90 ) & ( n11567 )  ;
assign n12815 =  ( n90 ) & ( n11569 )  ;
assign n12816 =  ( n90 ) & ( n11571 )  ;
assign n12817 =  ( n90 ) & ( n11573 )  ;
assign n12818 =  ( n90 ) & ( n11575 )  ;
assign n12819 =  ( n91 ) & ( n11545 )  ;
assign n12820 =  ( n91 ) & ( n11547 )  ;
assign n12821 =  ( n91 ) & ( n11549 )  ;
assign n12822 =  ( n91 ) & ( n11551 )  ;
assign n12823 =  ( n91 ) & ( n11553 )  ;
assign n12824 =  ( n91 ) & ( n11555 )  ;
assign n12825 =  ( n91 ) & ( n11557 )  ;
assign n12826 =  ( n91 ) & ( n11559 )  ;
assign n12827 =  ( n91 ) & ( n11561 )  ;
assign n12828 =  ( n91 ) & ( n11563 )  ;
assign n12829 =  ( n91 ) & ( n11565 )  ;
assign n12830 =  ( n91 ) & ( n11567 )  ;
assign n12831 =  ( n91 ) & ( n11569 )  ;
assign n12832 =  ( n91 ) & ( n11571 )  ;
assign n12833 =  ( n91 ) & ( n11573 )  ;
assign n12834 =  ( n91 ) & ( n11575 )  ;
assign n12835 =  ( n92 ) & ( n11545 )  ;
assign n12836 =  ( n92 ) & ( n11547 )  ;
assign n12837 =  ( n92 ) & ( n11549 )  ;
assign n12838 =  ( n92 ) & ( n11551 )  ;
assign n12839 =  ( n92 ) & ( n11553 )  ;
assign n12840 =  ( n92 ) & ( n11555 )  ;
assign n12841 =  ( n92 ) & ( n11557 )  ;
assign n12842 =  ( n92 ) & ( n11559 )  ;
assign n12843 =  ( n92 ) & ( n11561 )  ;
assign n12844 =  ( n92 ) & ( n11563 )  ;
assign n12845 =  ( n92 ) & ( n11565 )  ;
assign n12846 =  ( n92 ) & ( n11567 )  ;
assign n12847 =  ( n92 ) & ( n11569 )  ;
assign n12848 =  ( n92 ) & ( n11571 )  ;
assign n12849 =  ( n92 ) & ( n11573 )  ;
assign n12850 =  ( n92 ) & ( n11575 )  ;
assign n12851 =  ( n93 ) & ( n11545 )  ;
assign n12852 =  ( n93 ) & ( n11547 )  ;
assign n12853 =  ( n93 ) & ( n11549 )  ;
assign n12854 =  ( n93 ) & ( n11551 )  ;
assign n12855 =  ( n93 ) & ( n11553 )  ;
assign n12856 =  ( n93 ) & ( n11555 )  ;
assign n12857 =  ( n93 ) & ( n11557 )  ;
assign n12858 =  ( n93 ) & ( n11559 )  ;
assign n12859 =  ( n93 ) & ( n11561 )  ;
assign n12860 =  ( n93 ) & ( n11563 )  ;
assign n12861 =  ( n93 ) & ( n11565 )  ;
assign n12862 =  ( n93 ) & ( n11567 )  ;
assign n12863 =  ( n93 ) & ( n11569 )  ;
assign n12864 =  ( n93 ) & ( n11571 )  ;
assign n12865 =  ( n93 ) & ( n11573 )  ;
assign n12866 =  ( n93 ) & ( n11575 )  ;
assign n12867 =  ( n94 ) & ( n11545 )  ;
assign n12868 =  ( n94 ) & ( n11547 )  ;
assign n12869 =  ( n94 ) & ( n11549 )  ;
assign n12870 =  ( n94 ) & ( n11551 )  ;
assign n12871 =  ( n94 ) & ( n11553 )  ;
assign n12872 =  ( n94 ) & ( n11555 )  ;
assign n12873 =  ( n94 ) & ( n11557 )  ;
assign n12874 =  ( n94 ) & ( n11559 )  ;
assign n12875 =  ( n94 ) & ( n11561 )  ;
assign n12876 =  ( n94 ) & ( n11563 )  ;
assign n12877 =  ( n94 ) & ( n11565 )  ;
assign n12878 =  ( n94 ) & ( n11567 )  ;
assign n12879 =  ( n94 ) & ( n11569 )  ;
assign n12880 =  ( n94 ) & ( n11571 )  ;
assign n12881 =  ( n94 ) & ( n11573 )  ;
assign n12882 =  ( n94 ) & ( n11575 )  ;
assign n12883 =  ( n95 ) & ( n11545 )  ;
assign n12884 =  ( n95 ) & ( n11547 )  ;
assign n12885 =  ( n95 ) & ( n11549 )  ;
assign n12886 =  ( n95 ) & ( n11551 )  ;
assign n12887 =  ( n95 ) & ( n11553 )  ;
assign n12888 =  ( n95 ) & ( n11555 )  ;
assign n12889 =  ( n95 ) & ( n11557 )  ;
assign n12890 =  ( n95 ) & ( n11559 )  ;
assign n12891 =  ( n95 ) & ( n11561 )  ;
assign n12892 =  ( n95 ) & ( n11563 )  ;
assign n12893 =  ( n95 ) & ( n11565 )  ;
assign n12894 =  ( n95 ) & ( n11567 )  ;
assign n12895 =  ( n95 ) & ( n11569 )  ;
assign n12896 =  ( n95 ) & ( n11571 )  ;
assign n12897 =  ( n95 ) & ( n11573 )  ;
assign n12898 =  ( n95 ) & ( n11575 )  ;
assign n12899 =  ( n96 ) & ( n11545 )  ;
assign n12900 =  ( n96 ) & ( n11547 )  ;
assign n12901 =  ( n96 ) & ( n11549 )  ;
assign n12902 =  ( n96 ) & ( n11551 )  ;
assign n12903 =  ( n96 ) & ( n11553 )  ;
assign n12904 =  ( n96 ) & ( n11555 )  ;
assign n12905 =  ( n96 ) & ( n11557 )  ;
assign n12906 =  ( n96 ) & ( n11559 )  ;
assign n12907 =  ( n96 ) & ( n11561 )  ;
assign n12908 =  ( n96 ) & ( n11563 )  ;
assign n12909 =  ( n96 ) & ( n11565 )  ;
assign n12910 =  ( n96 ) & ( n11567 )  ;
assign n12911 =  ( n96 ) & ( n11569 )  ;
assign n12912 =  ( n96 ) & ( n11571 )  ;
assign n12913 =  ( n96 ) & ( n11573 )  ;
assign n12914 =  ( n96 ) & ( n11575 )  ;
assign n12915 =  ( n97 ) & ( n11545 )  ;
assign n12916 =  ( n97 ) & ( n11547 )  ;
assign n12917 =  ( n97 ) & ( n11549 )  ;
assign n12918 =  ( n97 ) & ( n11551 )  ;
assign n12919 =  ( n97 ) & ( n11553 )  ;
assign n12920 =  ( n97 ) & ( n11555 )  ;
assign n12921 =  ( n97 ) & ( n11557 )  ;
assign n12922 =  ( n97 ) & ( n11559 )  ;
assign n12923 =  ( n97 ) & ( n11561 )  ;
assign n12924 =  ( n97 ) & ( n11563 )  ;
assign n12925 =  ( n97 ) & ( n11565 )  ;
assign n12926 =  ( n97 ) & ( n11567 )  ;
assign n12927 =  ( n97 ) & ( n11569 )  ;
assign n12928 =  ( n97 ) & ( n11571 )  ;
assign n12929 =  ( n97 ) & ( n11573 )  ;
assign n12930 =  ( n97 ) & ( n11575 )  ;
assign n12931 =  ( n98 ) & ( n11545 )  ;
assign n12932 =  ( n98 ) & ( n11547 )  ;
assign n12933 =  ( n98 ) & ( n11549 )  ;
assign n12934 =  ( n98 ) & ( n11551 )  ;
assign n12935 =  ( n98 ) & ( n11553 )  ;
assign n12936 =  ( n98 ) & ( n11555 )  ;
assign n12937 =  ( n98 ) & ( n11557 )  ;
assign n12938 =  ( n98 ) & ( n11559 )  ;
assign n12939 =  ( n98 ) & ( n11561 )  ;
assign n12940 =  ( n98 ) & ( n11563 )  ;
assign n12941 =  ( n98 ) & ( n11565 )  ;
assign n12942 =  ( n98 ) & ( n11567 )  ;
assign n12943 =  ( n98 ) & ( n11569 )  ;
assign n12944 =  ( n98 ) & ( n11571 )  ;
assign n12945 =  ( n98 ) & ( n11573 )  ;
assign n12946 =  ( n98 ) & ( n11575 )  ;
assign n12947 =  ( n99 ) & ( n11545 )  ;
assign n12948 =  ( n99 ) & ( n11547 )  ;
assign n12949 =  ( n99 ) & ( n11549 )  ;
assign n12950 =  ( n99 ) & ( n11551 )  ;
assign n12951 =  ( n99 ) & ( n11553 )  ;
assign n12952 =  ( n99 ) & ( n11555 )  ;
assign n12953 =  ( n99 ) & ( n11557 )  ;
assign n12954 =  ( n99 ) & ( n11559 )  ;
assign n12955 =  ( n99 ) & ( n11561 )  ;
assign n12956 =  ( n99 ) & ( n11563 )  ;
assign n12957 =  ( n99 ) & ( n11565 )  ;
assign n12958 =  ( n99 ) & ( n11567 )  ;
assign n12959 =  ( n99 ) & ( n11569 )  ;
assign n12960 =  ( n99 ) & ( n11571 )  ;
assign n12961 =  ( n99 ) & ( n11573 )  ;
assign n12962 =  ( n99 ) & ( n11575 )  ;
assign n12963 =  ( n100 ) & ( n11545 )  ;
assign n12964 =  ( n100 ) & ( n11547 )  ;
assign n12965 =  ( n100 ) & ( n11549 )  ;
assign n12966 =  ( n100 ) & ( n11551 )  ;
assign n12967 =  ( n100 ) & ( n11553 )  ;
assign n12968 =  ( n100 ) & ( n11555 )  ;
assign n12969 =  ( n100 ) & ( n11557 )  ;
assign n12970 =  ( n100 ) & ( n11559 )  ;
assign n12971 =  ( n100 ) & ( n11561 )  ;
assign n12972 =  ( n100 ) & ( n11563 )  ;
assign n12973 =  ( n100 ) & ( n11565 )  ;
assign n12974 =  ( n100 ) & ( n11567 )  ;
assign n12975 =  ( n100 ) & ( n11569 )  ;
assign n12976 =  ( n100 ) & ( n11571 )  ;
assign n12977 =  ( n100 ) & ( n11573 )  ;
assign n12978 =  ( n100 ) & ( n11575 )  ;
assign n12979 =  ( n101 ) & ( n11545 )  ;
assign n12980 =  ( n101 ) & ( n11547 )  ;
assign n12981 =  ( n101 ) & ( n11549 )  ;
assign n12982 =  ( n101 ) & ( n11551 )  ;
assign n12983 =  ( n101 ) & ( n11553 )  ;
assign n12984 =  ( n101 ) & ( n11555 )  ;
assign n12985 =  ( n101 ) & ( n11557 )  ;
assign n12986 =  ( n101 ) & ( n11559 )  ;
assign n12987 =  ( n101 ) & ( n11561 )  ;
assign n12988 =  ( n101 ) & ( n11563 )  ;
assign n12989 =  ( n101 ) & ( n11565 )  ;
assign n12990 =  ( n101 ) & ( n11567 )  ;
assign n12991 =  ( n101 ) & ( n11569 )  ;
assign n12992 =  ( n101 ) & ( n11571 )  ;
assign n12993 =  ( n101 ) & ( n11573 )  ;
assign n12994 =  ( n101 ) & ( n11575 )  ;
assign n12995 =  ( n102 ) & ( n11545 )  ;
assign n12996 =  ( n102 ) & ( n11547 )  ;
assign n12997 =  ( n102 ) & ( n11549 )  ;
assign n12998 =  ( n102 ) & ( n11551 )  ;
assign n12999 =  ( n102 ) & ( n11553 )  ;
assign n13000 =  ( n102 ) & ( n11555 )  ;
assign n13001 =  ( n102 ) & ( n11557 )  ;
assign n13002 =  ( n102 ) & ( n11559 )  ;
assign n13003 =  ( n102 ) & ( n11561 )  ;
assign n13004 =  ( n102 ) & ( n11563 )  ;
assign n13005 =  ( n102 ) & ( n11565 )  ;
assign n13006 =  ( n102 ) & ( n11567 )  ;
assign n13007 =  ( n102 ) & ( n11569 )  ;
assign n13008 =  ( n102 ) & ( n11571 )  ;
assign n13009 =  ( n102 ) & ( n11573 )  ;
assign n13010 =  ( n102 ) & ( n11575 )  ;
assign n13011 =  ( n103 ) & ( n11545 )  ;
assign n13012 =  ( n103 ) & ( n11547 )  ;
assign n13013 =  ( n103 ) & ( n11549 )  ;
assign n13014 =  ( n103 ) & ( n11551 )  ;
assign n13015 =  ( n103 ) & ( n11553 )  ;
assign n13016 =  ( n103 ) & ( n11555 )  ;
assign n13017 =  ( n103 ) & ( n11557 )  ;
assign n13018 =  ( n103 ) & ( n11559 )  ;
assign n13019 =  ( n103 ) & ( n11561 )  ;
assign n13020 =  ( n103 ) & ( n11563 )  ;
assign n13021 =  ( n103 ) & ( n11565 )  ;
assign n13022 =  ( n103 ) & ( n11567 )  ;
assign n13023 =  ( n103 ) & ( n11569 )  ;
assign n13024 =  ( n103 ) & ( n11571 )  ;
assign n13025 =  ( n103 ) & ( n11573 )  ;
assign n13026 =  ( n103 ) & ( n11575 )  ;
assign n13027 =  ( n104 ) & ( n11545 )  ;
assign n13028 =  ( n104 ) & ( n11547 )  ;
assign n13029 =  ( n104 ) & ( n11549 )  ;
assign n13030 =  ( n104 ) & ( n11551 )  ;
assign n13031 =  ( n104 ) & ( n11553 )  ;
assign n13032 =  ( n104 ) & ( n11555 )  ;
assign n13033 =  ( n104 ) & ( n11557 )  ;
assign n13034 =  ( n104 ) & ( n11559 )  ;
assign n13035 =  ( n104 ) & ( n11561 )  ;
assign n13036 =  ( n104 ) & ( n11563 )  ;
assign n13037 =  ( n104 ) & ( n11565 )  ;
assign n13038 =  ( n104 ) & ( n11567 )  ;
assign n13039 =  ( n104 ) & ( n11569 )  ;
assign n13040 =  ( n104 ) & ( n11571 )  ;
assign n13041 =  ( n104 ) & ( n11573 )  ;
assign n13042 =  ( n104 ) & ( n11575 )  ;
assign n13043 =  ( n105 ) & ( n11545 )  ;
assign n13044 =  ( n105 ) & ( n11547 )  ;
assign n13045 =  ( n105 ) & ( n11549 )  ;
assign n13046 =  ( n105 ) & ( n11551 )  ;
assign n13047 =  ( n105 ) & ( n11553 )  ;
assign n13048 =  ( n105 ) & ( n11555 )  ;
assign n13049 =  ( n105 ) & ( n11557 )  ;
assign n13050 =  ( n105 ) & ( n11559 )  ;
assign n13051 =  ( n105 ) & ( n11561 )  ;
assign n13052 =  ( n105 ) & ( n11563 )  ;
assign n13053 =  ( n105 ) & ( n11565 )  ;
assign n13054 =  ( n105 ) & ( n11567 )  ;
assign n13055 =  ( n105 ) & ( n11569 )  ;
assign n13056 =  ( n105 ) & ( n11571 )  ;
assign n13057 =  ( n105 ) & ( n11573 )  ;
assign n13058 =  ( n105 ) & ( n11575 )  ;
assign n13059 =  ( n106 ) & ( n11545 )  ;
assign n13060 =  ( n106 ) & ( n11547 )  ;
assign n13061 =  ( n106 ) & ( n11549 )  ;
assign n13062 =  ( n106 ) & ( n11551 )  ;
assign n13063 =  ( n106 ) & ( n11553 )  ;
assign n13064 =  ( n106 ) & ( n11555 )  ;
assign n13065 =  ( n106 ) & ( n11557 )  ;
assign n13066 =  ( n106 ) & ( n11559 )  ;
assign n13067 =  ( n106 ) & ( n11561 )  ;
assign n13068 =  ( n106 ) & ( n11563 )  ;
assign n13069 =  ( n106 ) & ( n11565 )  ;
assign n13070 =  ( n106 ) & ( n11567 )  ;
assign n13071 =  ( n106 ) & ( n11569 )  ;
assign n13072 =  ( n106 ) & ( n11571 )  ;
assign n13073 =  ( n106 ) & ( n11573 )  ;
assign n13074 =  ( n106 ) & ( n11575 )  ;
assign n13075 =  ( n107 ) & ( n11545 )  ;
assign n13076 =  ( n107 ) & ( n11547 )  ;
assign n13077 =  ( n107 ) & ( n11549 )  ;
assign n13078 =  ( n107 ) & ( n11551 )  ;
assign n13079 =  ( n107 ) & ( n11553 )  ;
assign n13080 =  ( n107 ) & ( n11555 )  ;
assign n13081 =  ( n107 ) & ( n11557 )  ;
assign n13082 =  ( n107 ) & ( n11559 )  ;
assign n13083 =  ( n107 ) & ( n11561 )  ;
assign n13084 =  ( n107 ) & ( n11563 )  ;
assign n13085 =  ( n107 ) & ( n11565 )  ;
assign n13086 =  ( n107 ) & ( n11567 )  ;
assign n13087 =  ( n107 ) & ( n11569 )  ;
assign n13088 =  ( n107 ) & ( n11571 )  ;
assign n13089 =  ( n107 ) & ( n11573 )  ;
assign n13090 =  ( n107 ) & ( n11575 )  ;
assign n13091 =  ( n108 ) & ( n11545 )  ;
assign n13092 =  ( n108 ) & ( n11547 )  ;
assign n13093 =  ( n108 ) & ( n11549 )  ;
assign n13094 =  ( n108 ) & ( n11551 )  ;
assign n13095 =  ( n108 ) & ( n11553 )  ;
assign n13096 =  ( n108 ) & ( n11555 )  ;
assign n13097 =  ( n108 ) & ( n11557 )  ;
assign n13098 =  ( n108 ) & ( n11559 )  ;
assign n13099 =  ( n108 ) & ( n11561 )  ;
assign n13100 =  ( n108 ) & ( n11563 )  ;
assign n13101 =  ( n108 ) & ( n11565 )  ;
assign n13102 =  ( n108 ) & ( n11567 )  ;
assign n13103 =  ( n108 ) & ( n11569 )  ;
assign n13104 =  ( n108 ) & ( n11571 )  ;
assign n13105 =  ( n108 ) & ( n11573 )  ;
assign n13106 =  ( n108 ) & ( n11575 )  ;
assign n13107 =  ( n13106 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n13108 =  ( n13105 ) ? ( VREG_0_1 ) : ( n13107 ) ;
assign n13109 =  ( n13104 ) ? ( VREG_0_2 ) : ( n13108 ) ;
assign n13110 =  ( n13103 ) ? ( VREG_0_3 ) : ( n13109 ) ;
assign n13111 =  ( n13102 ) ? ( VREG_0_4 ) : ( n13110 ) ;
assign n13112 =  ( n13101 ) ? ( VREG_0_5 ) : ( n13111 ) ;
assign n13113 =  ( n13100 ) ? ( VREG_0_6 ) : ( n13112 ) ;
assign n13114 =  ( n13099 ) ? ( VREG_0_7 ) : ( n13113 ) ;
assign n13115 =  ( n13098 ) ? ( VREG_0_8 ) : ( n13114 ) ;
assign n13116 =  ( n13097 ) ? ( VREG_0_9 ) : ( n13115 ) ;
assign n13117 =  ( n13096 ) ? ( VREG_0_10 ) : ( n13116 ) ;
assign n13118 =  ( n13095 ) ? ( VREG_0_11 ) : ( n13117 ) ;
assign n13119 =  ( n13094 ) ? ( VREG_0_12 ) : ( n13118 ) ;
assign n13120 =  ( n13093 ) ? ( VREG_0_13 ) : ( n13119 ) ;
assign n13121 =  ( n13092 ) ? ( VREG_0_14 ) : ( n13120 ) ;
assign n13122 =  ( n13091 ) ? ( VREG_0_15 ) : ( n13121 ) ;
assign n13123 =  ( n13090 ) ? ( VREG_1_0 ) : ( n13122 ) ;
assign n13124 =  ( n13089 ) ? ( VREG_1_1 ) : ( n13123 ) ;
assign n13125 =  ( n13088 ) ? ( VREG_1_2 ) : ( n13124 ) ;
assign n13126 =  ( n13087 ) ? ( VREG_1_3 ) : ( n13125 ) ;
assign n13127 =  ( n13086 ) ? ( VREG_1_4 ) : ( n13126 ) ;
assign n13128 =  ( n13085 ) ? ( VREG_1_5 ) : ( n13127 ) ;
assign n13129 =  ( n13084 ) ? ( VREG_1_6 ) : ( n13128 ) ;
assign n13130 =  ( n13083 ) ? ( VREG_1_7 ) : ( n13129 ) ;
assign n13131 =  ( n13082 ) ? ( VREG_1_8 ) : ( n13130 ) ;
assign n13132 =  ( n13081 ) ? ( VREG_1_9 ) : ( n13131 ) ;
assign n13133 =  ( n13080 ) ? ( VREG_1_10 ) : ( n13132 ) ;
assign n13134 =  ( n13079 ) ? ( VREG_1_11 ) : ( n13133 ) ;
assign n13135 =  ( n13078 ) ? ( VREG_1_12 ) : ( n13134 ) ;
assign n13136 =  ( n13077 ) ? ( VREG_1_13 ) : ( n13135 ) ;
assign n13137 =  ( n13076 ) ? ( VREG_1_14 ) : ( n13136 ) ;
assign n13138 =  ( n13075 ) ? ( VREG_1_15 ) : ( n13137 ) ;
assign n13139 =  ( n13074 ) ? ( VREG_2_0 ) : ( n13138 ) ;
assign n13140 =  ( n13073 ) ? ( VREG_2_1 ) : ( n13139 ) ;
assign n13141 =  ( n13072 ) ? ( VREG_2_2 ) : ( n13140 ) ;
assign n13142 =  ( n13071 ) ? ( VREG_2_3 ) : ( n13141 ) ;
assign n13143 =  ( n13070 ) ? ( VREG_2_4 ) : ( n13142 ) ;
assign n13144 =  ( n13069 ) ? ( VREG_2_5 ) : ( n13143 ) ;
assign n13145 =  ( n13068 ) ? ( VREG_2_6 ) : ( n13144 ) ;
assign n13146 =  ( n13067 ) ? ( VREG_2_7 ) : ( n13145 ) ;
assign n13147 =  ( n13066 ) ? ( VREG_2_8 ) : ( n13146 ) ;
assign n13148 =  ( n13065 ) ? ( VREG_2_9 ) : ( n13147 ) ;
assign n13149 =  ( n13064 ) ? ( VREG_2_10 ) : ( n13148 ) ;
assign n13150 =  ( n13063 ) ? ( VREG_2_11 ) : ( n13149 ) ;
assign n13151 =  ( n13062 ) ? ( VREG_2_12 ) : ( n13150 ) ;
assign n13152 =  ( n13061 ) ? ( VREG_2_13 ) : ( n13151 ) ;
assign n13153 =  ( n13060 ) ? ( VREG_2_14 ) : ( n13152 ) ;
assign n13154 =  ( n13059 ) ? ( VREG_2_15 ) : ( n13153 ) ;
assign n13155 =  ( n13058 ) ? ( VREG_3_0 ) : ( n13154 ) ;
assign n13156 =  ( n13057 ) ? ( VREG_3_1 ) : ( n13155 ) ;
assign n13157 =  ( n13056 ) ? ( VREG_3_2 ) : ( n13156 ) ;
assign n13158 =  ( n13055 ) ? ( VREG_3_3 ) : ( n13157 ) ;
assign n13159 =  ( n13054 ) ? ( VREG_3_4 ) : ( n13158 ) ;
assign n13160 =  ( n13053 ) ? ( VREG_3_5 ) : ( n13159 ) ;
assign n13161 =  ( n13052 ) ? ( VREG_3_6 ) : ( n13160 ) ;
assign n13162 =  ( n13051 ) ? ( VREG_3_7 ) : ( n13161 ) ;
assign n13163 =  ( n13050 ) ? ( VREG_3_8 ) : ( n13162 ) ;
assign n13164 =  ( n13049 ) ? ( VREG_3_9 ) : ( n13163 ) ;
assign n13165 =  ( n13048 ) ? ( VREG_3_10 ) : ( n13164 ) ;
assign n13166 =  ( n13047 ) ? ( VREG_3_11 ) : ( n13165 ) ;
assign n13167 =  ( n13046 ) ? ( VREG_3_12 ) : ( n13166 ) ;
assign n13168 =  ( n13045 ) ? ( VREG_3_13 ) : ( n13167 ) ;
assign n13169 =  ( n13044 ) ? ( VREG_3_14 ) : ( n13168 ) ;
assign n13170 =  ( n13043 ) ? ( VREG_3_15 ) : ( n13169 ) ;
assign n13171 =  ( n13042 ) ? ( VREG_4_0 ) : ( n13170 ) ;
assign n13172 =  ( n13041 ) ? ( VREG_4_1 ) : ( n13171 ) ;
assign n13173 =  ( n13040 ) ? ( VREG_4_2 ) : ( n13172 ) ;
assign n13174 =  ( n13039 ) ? ( VREG_4_3 ) : ( n13173 ) ;
assign n13175 =  ( n13038 ) ? ( VREG_4_4 ) : ( n13174 ) ;
assign n13176 =  ( n13037 ) ? ( VREG_4_5 ) : ( n13175 ) ;
assign n13177 =  ( n13036 ) ? ( VREG_4_6 ) : ( n13176 ) ;
assign n13178 =  ( n13035 ) ? ( VREG_4_7 ) : ( n13177 ) ;
assign n13179 =  ( n13034 ) ? ( VREG_4_8 ) : ( n13178 ) ;
assign n13180 =  ( n13033 ) ? ( VREG_4_9 ) : ( n13179 ) ;
assign n13181 =  ( n13032 ) ? ( VREG_4_10 ) : ( n13180 ) ;
assign n13182 =  ( n13031 ) ? ( VREG_4_11 ) : ( n13181 ) ;
assign n13183 =  ( n13030 ) ? ( VREG_4_12 ) : ( n13182 ) ;
assign n13184 =  ( n13029 ) ? ( VREG_4_13 ) : ( n13183 ) ;
assign n13185 =  ( n13028 ) ? ( VREG_4_14 ) : ( n13184 ) ;
assign n13186 =  ( n13027 ) ? ( VREG_4_15 ) : ( n13185 ) ;
assign n13187 =  ( n13026 ) ? ( VREG_5_0 ) : ( n13186 ) ;
assign n13188 =  ( n13025 ) ? ( VREG_5_1 ) : ( n13187 ) ;
assign n13189 =  ( n13024 ) ? ( VREG_5_2 ) : ( n13188 ) ;
assign n13190 =  ( n13023 ) ? ( VREG_5_3 ) : ( n13189 ) ;
assign n13191 =  ( n13022 ) ? ( VREG_5_4 ) : ( n13190 ) ;
assign n13192 =  ( n13021 ) ? ( VREG_5_5 ) : ( n13191 ) ;
assign n13193 =  ( n13020 ) ? ( VREG_5_6 ) : ( n13192 ) ;
assign n13194 =  ( n13019 ) ? ( VREG_5_7 ) : ( n13193 ) ;
assign n13195 =  ( n13018 ) ? ( VREG_5_8 ) : ( n13194 ) ;
assign n13196 =  ( n13017 ) ? ( VREG_5_9 ) : ( n13195 ) ;
assign n13197 =  ( n13016 ) ? ( VREG_5_10 ) : ( n13196 ) ;
assign n13198 =  ( n13015 ) ? ( VREG_5_11 ) : ( n13197 ) ;
assign n13199 =  ( n13014 ) ? ( VREG_5_12 ) : ( n13198 ) ;
assign n13200 =  ( n13013 ) ? ( VREG_5_13 ) : ( n13199 ) ;
assign n13201 =  ( n13012 ) ? ( VREG_5_14 ) : ( n13200 ) ;
assign n13202 =  ( n13011 ) ? ( VREG_5_15 ) : ( n13201 ) ;
assign n13203 =  ( n13010 ) ? ( VREG_6_0 ) : ( n13202 ) ;
assign n13204 =  ( n13009 ) ? ( VREG_6_1 ) : ( n13203 ) ;
assign n13205 =  ( n13008 ) ? ( VREG_6_2 ) : ( n13204 ) ;
assign n13206 =  ( n13007 ) ? ( VREG_6_3 ) : ( n13205 ) ;
assign n13207 =  ( n13006 ) ? ( VREG_6_4 ) : ( n13206 ) ;
assign n13208 =  ( n13005 ) ? ( VREG_6_5 ) : ( n13207 ) ;
assign n13209 =  ( n13004 ) ? ( VREG_6_6 ) : ( n13208 ) ;
assign n13210 =  ( n13003 ) ? ( VREG_6_7 ) : ( n13209 ) ;
assign n13211 =  ( n13002 ) ? ( VREG_6_8 ) : ( n13210 ) ;
assign n13212 =  ( n13001 ) ? ( VREG_6_9 ) : ( n13211 ) ;
assign n13213 =  ( n13000 ) ? ( VREG_6_10 ) : ( n13212 ) ;
assign n13214 =  ( n12999 ) ? ( VREG_6_11 ) : ( n13213 ) ;
assign n13215 =  ( n12998 ) ? ( VREG_6_12 ) : ( n13214 ) ;
assign n13216 =  ( n12997 ) ? ( VREG_6_13 ) : ( n13215 ) ;
assign n13217 =  ( n12996 ) ? ( VREG_6_14 ) : ( n13216 ) ;
assign n13218 =  ( n12995 ) ? ( VREG_6_15 ) : ( n13217 ) ;
assign n13219 =  ( n12994 ) ? ( VREG_7_0 ) : ( n13218 ) ;
assign n13220 =  ( n12993 ) ? ( VREG_7_1 ) : ( n13219 ) ;
assign n13221 =  ( n12992 ) ? ( VREG_7_2 ) : ( n13220 ) ;
assign n13222 =  ( n12991 ) ? ( VREG_7_3 ) : ( n13221 ) ;
assign n13223 =  ( n12990 ) ? ( VREG_7_4 ) : ( n13222 ) ;
assign n13224 =  ( n12989 ) ? ( VREG_7_5 ) : ( n13223 ) ;
assign n13225 =  ( n12988 ) ? ( VREG_7_6 ) : ( n13224 ) ;
assign n13226 =  ( n12987 ) ? ( VREG_7_7 ) : ( n13225 ) ;
assign n13227 =  ( n12986 ) ? ( VREG_7_8 ) : ( n13226 ) ;
assign n13228 =  ( n12985 ) ? ( VREG_7_9 ) : ( n13227 ) ;
assign n13229 =  ( n12984 ) ? ( VREG_7_10 ) : ( n13228 ) ;
assign n13230 =  ( n12983 ) ? ( VREG_7_11 ) : ( n13229 ) ;
assign n13231 =  ( n12982 ) ? ( VREG_7_12 ) : ( n13230 ) ;
assign n13232 =  ( n12981 ) ? ( VREG_7_13 ) : ( n13231 ) ;
assign n13233 =  ( n12980 ) ? ( VREG_7_14 ) : ( n13232 ) ;
assign n13234 =  ( n12979 ) ? ( VREG_7_15 ) : ( n13233 ) ;
assign n13235 =  ( n12978 ) ? ( VREG_8_0 ) : ( n13234 ) ;
assign n13236 =  ( n12977 ) ? ( VREG_8_1 ) : ( n13235 ) ;
assign n13237 =  ( n12976 ) ? ( VREG_8_2 ) : ( n13236 ) ;
assign n13238 =  ( n12975 ) ? ( VREG_8_3 ) : ( n13237 ) ;
assign n13239 =  ( n12974 ) ? ( VREG_8_4 ) : ( n13238 ) ;
assign n13240 =  ( n12973 ) ? ( VREG_8_5 ) : ( n13239 ) ;
assign n13241 =  ( n12972 ) ? ( VREG_8_6 ) : ( n13240 ) ;
assign n13242 =  ( n12971 ) ? ( VREG_8_7 ) : ( n13241 ) ;
assign n13243 =  ( n12970 ) ? ( VREG_8_8 ) : ( n13242 ) ;
assign n13244 =  ( n12969 ) ? ( VREG_8_9 ) : ( n13243 ) ;
assign n13245 =  ( n12968 ) ? ( VREG_8_10 ) : ( n13244 ) ;
assign n13246 =  ( n12967 ) ? ( VREG_8_11 ) : ( n13245 ) ;
assign n13247 =  ( n12966 ) ? ( VREG_8_12 ) : ( n13246 ) ;
assign n13248 =  ( n12965 ) ? ( VREG_8_13 ) : ( n13247 ) ;
assign n13249 =  ( n12964 ) ? ( VREG_8_14 ) : ( n13248 ) ;
assign n13250 =  ( n12963 ) ? ( VREG_8_15 ) : ( n13249 ) ;
assign n13251 =  ( n12962 ) ? ( VREG_9_0 ) : ( n13250 ) ;
assign n13252 =  ( n12961 ) ? ( VREG_9_1 ) : ( n13251 ) ;
assign n13253 =  ( n12960 ) ? ( VREG_9_2 ) : ( n13252 ) ;
assign n13254 =  ( n12959 ) ? ( VREG_9_3 ) : ( n13253 ) ;
assign n13255 =  ( n12958 ) ? ( VREG_9_4 ) : ( n13254 ) ;
assign n13256 =  ( n12957 ) ? ( VREG_9_5 ) : ( n13255 ) ;
assign n13257 =  ( n12956 ) ? ( VREG_9_6 ) : ( n13256 ) ;
assign n13258 =  ( n12955 ) ? ( VREG_9_7 ) : ( n13257 ) ;
assign n13259 =  ( n12954 ) ? ( VREG_9_8 ) : ( n13258 ) ;
assign n13260 =  ( n12953 ) ? ( VREG_9_9 ) : ( n13259 ) ;
assign n13261 =  ( n12952 ) ? ( VREG_9_10 ) : ( n13260 ) ;
assign n13262 =  ( n12951 ) ? ( VREG_9_11 ) : ( n13261 ) ;
assign n13263 =  ( n12950 ) ? ( VREG_9_12 ) : ( n13262 ) ;
assign n13264 =  ( n12949 ) ? ( VREG_9_13 ) : ( n13263 ) ;
assign n13265 =  ( n12948 ) ? ( VREG_9_14 ) : ( n13264 ) ;
assign n13266 =  ( n12947 ) ? ( VREG_9_15 ) : ( n13265 ) ;
assign n13267 =  ( n12946 ) ? ( VREG_10_0 ) : ( n13266 ) ;
assign n13268 =  ( n12945 ) ? ( VREG_10_1 ) : ( n13267 ) ;
assign n13269 =  ( n12944 ) ? ( VREG_10_2 ) : ( n13268 ) ;
assign n13270 =  ( n12943 ) ? ( VREG_10_3 ) : ( n13269 ) ;
assign n13271 =  ( n12942 ) ? ( VREG_10_4 ) : ( n13270 ) ;
assign n13272 =  ( n12941 ) ? ( VREG_10_5 ) : ( n13271 ) ;
assign n13273 =  ( n12940 ) ? ( VREG_10_6 ) : ( n13272 ) ;
assign n13274 =  ( n12939 ) ? ( VREG_10_7 ) : ( n13273 ) ;
assign n13275 =  ( n12938 ) ? ( VREG_10_8 ) : ( n13274 ) ;
assign n13276 =  ( n12937 ) ? ( VREG_10_9 ) : ( n13275 ) ;
assign n13277 =  ( n12936 ) ? ( VREG_10_10 ) : ( n13276 ) ;
assign n13278 =  ( n12935 ) ? ( VREG_10_11 ) : ( n13277 ) ;
assign n13279 =  ( n12934 ) ? ( VREG_10_12 ) : ( n13278 ) ;
assign n13280 =  ( n12933 ) ? ( VREG_10_13 ) : ( n13279 ) ;
assign n13281 =  ( n12932 ) ? ( VREG_10_14 ) : ( n13280 ) ;
assign n13282 =  ( n12931 ) ? ( VREG_10_15 ) : ( n13281 ) ;
assign n13283 =  ( n12930 ) ? ( VREG_11_0 ) : ( n13282 ) ;
assign n13284 =  ( n12929 ) ? ( VREG_11_1 ) : ( n13283 ) ;
assign n13285 =  ( n12928 ) ? ( VREG_11_2 ) : ( n13284 ) ;
assign n13286 =  ( n12927 ) ? ( VREG_11_3 ) : ( n13285 ) ;
assign n13287 =  ( n12926 ) ? ( VREG_11_4 ) : ( n13286 ) ;
assign n13288 =  ( n12925 ) ? ( VREG_11_5 ) : ( n13287 ) ;
assign n13289 =  ( n12924 ) ? ( VREG_11_6 ) : ( n13288 ) ;
assign n13290 =  ( n12923 ) ? ( VREG_11_7 ) : ( n13289 ) ;
assign n13291 =  ( n12922 ) ? ( VREG_11_8 ) : ( n13290 ) ;
assign n13292 =  ( n12921 ) ? ( VREG_11_9 ) : ( n13291 ) ;
assign n13293 =  ( n12920 ) ? ( VREG_11_10 ) : ( n13292 ) ;
assign n13294 =  ( n12919 ) ? ( VREG_11_11 ) : ( n13293 ) ;
assign n13295 =  ( n12918 ) ? ( VREG_11_12 ) : ( n13294 ) ;
assign n13296 =  ( n12917 ) ? ( VREG_11_13 ) : ( n13295 ) ;
assign n13297 =  ( n12916 ) ? ( VREG_11_14 ) : ( n13296 ) ;
assign n13298 =  ( n12915 ) ? ( VREG_11_15 ) : ( n13297 ) ;
assign n13299 =  ( n12914 ) ? ( VREG_12_0 ) : ( n13298 ) ;
assign n13300 =  ( n12913 ) ? ( VREG_12_1 ) : ( n13299 ) ;
assign n13301 =  ( n12912 ) ? ( VREG_12_2 ) : ( n13300 ) ;
assign n13302 =  ( n12911 ) ? ( VREG_12_3 ) : ( n13301 ) ;
assign n13303 =  ( n12910 ) ? ( VREG_12_4 ) : ( n13302 ) ;
assign n13304 =  ( n12909 ) ? ( VREG_12_5 ) : ( n13303 ) ;
assign n13305 =  ( n12908 ) ? ( VREG_12_6 ) : ( n13304 ) ;
assign n13306 =  ( n12907 ) ? ( VREG_12_7 ) : ( n13305 ) ;
assign n13307 =  ( n12906 ) ? ( VREG_12_8 ) : ( n13306 ) ;
assign n13308 =  ( n12905 ) ? ( VREG_12_9 ) : ( n13307 ) ;
assign n13309 =  ( n12904 ) ? ( VREG_12_10 ) : ( n13308 ) ;
assign n13310 =  ( n12903 ) ? ( VREG_12_11 ) : ( n13309 ) ;
assign n13311 =  ( n12902 ) ? ( VREG_12_12 ) : ( n13310 ) ;
assign n13312 =  ( n12901 ) ? ( VREG_12_13 ) : ( n13311 ) ;
assign n13313 =  ( n12900 ) ? ( VREG_12_14 ) : ( n13312 ) ;
assign n13314 =  ( n12899 ) ? ( VREG_12_15 ) : ( n13313 ) ;
assign n13315 =  ( n12898 ) ? ( VREG_13_0 ) : ( n13314 ) ;
assign n13316 =  ( n12897 ) ? ( VREG_13_1 ) : ( n13315 ) ;
assign n13317 =  ( n12896 ) ? ( VREG_13_2 ) : ( n13316 ) ;
assign n13318 =  ( n12895 ) ? ( VREG_13_3 ) : ( n13317 ) ;
assign n13319 =  ( n12894 ) ? ( VREG_13_4 ) : ( n13318 ) ;
assign n13320 =  ( n12893 ) ? ( VREG_13_5 ) : ( n13319 ) ;
assign n13321 =  ( n12892 ) ? ( VREG_13_6 ) : ( n13320 ) ;
assign n13322 =  ( n12891 ) ? ( VREG_13_7 ) : ( n13321 ) ;
assign n13323 =  ( n12890 ) ? ( VREG_13_8 ) : ( n13322 ) ;
assign n13324 =  ( n12889 ) ? ( VREG_13_9 ) : ( n13323 ) ;
assign n13325 =  ( n12888 ) ? ( VREG_13_10 ) : ( n13324 ) ;
assign n13326 =  ( n12887 ) ? ( VREG_13_11 ) : ( n13325 ) ;
assign n13327 =  ( n12886 ) ? ( VREG_13_12 ) : ( n13326 ) ;
assign n13328 =  ( n12885 ) ? ( VREG_13_13 ) : ( n13327 ) ;
assign n13329 =  ( n12884 ) ? ( VREG_13_14 ) : ( n13328 ) ;
assign n13330 =  ( n12883 ) ? ( VREG_13_15 ) : ( n13329 ) ;
assign n13331 =  ( n12882 ) ? ( VREG_14_0 ) : ( n13330 ) ;
assign n13332 =  ( n12881 ) ? ( VREG_14_1 ) : ( n13331 ) ;
assign n13333 =  ( n12880 ) ? ( VREG_14_2 ) : ( n13332 ) ;
assign n13334 =  ( n12879 ) ? ( VREG_14_3 ) : ( n13333 ) ;
assign n13335 =  ( n12878 ) ? ( VREG_14_4 ) : ( n13334 ) ;
assign n13336 =  ( n12877 ) ? ( VREG_14_5 ) : ( n13335 ) ;
assign n13337 =  ( n12876 ) ? ( VREG_14_6 ) : ( n13336 ) ;
assign n13338 =  ( n12875 ) ? ( VREG_14_7 ) : ( n13337 ) ;
assign n13339 =  ( n12874 ) ? ( VREG_14_8 ) : ( n13338 ) ;
assign n13340 =  ( n12873 ) ? ( VREG_14_9 ) : ( n13339 ) ;
assign n13341 =  ( n12872 ) ? ( VREG_14_10 ) : ( n13340 ) ;
assign n13342 =  ( n12871 ) ? ( VREG_14_11 ) : ( n13341 ) ;
assign n13343 =  ( n12870 ) ? ( VREG_14_12 ) : ( n13342 ) ;
assign n13344 =  ( n12869 ) ? ( VREG_14_13 ) : ( n13343 ) ;
assign n13345 =  ( n12868 ) ? ( VREG_14_14 ) : ( n13344 ) ;
assign n13346 =  ( n12867 ) ? ( VREG_14_15 ) : ( n13345 ) ;
assign n13347 =  ( n12866 ) ? ( VREG_15_0 ) : ( n13346 ) ;
assign n13348 =  ( n12865 ) ? ( VREG_15_1 ) : ( n13347 ) ;
assign n13349 =  ( n12864 ) ? ( VREG_15_2 ) : ( n13348 ) ;
assign n13350 =  ( n12863 ) ? ( VREG_15_3 ) : ( n13349 ) ;
assign n13351 =  ( n12862 ) ? ( VREG_15_4 ) : ( n13350 ) ;
assign n13352 =  ( n12861 ) ? ( VREG_15_5 ) : ( n13351 ) ;
assign n13353 =  ( n12860 ) ? ( VREG_15_6 ) : ( n13352 ) ;
assign n13354 =  ( n12859 ) ? ( VREG_15_7 ) : ( n13353 ) ;
assign n13355 =  ( n12858 ) ? ( VREG_15_8 ) : ( n13354 ) ;
assign n13356 =  ( n12857 ) ? ( VREG_15_9 ) : ( n13355 ) ;
assign n13357 =  ( n12856 ) ? ( VREG_15_10 ) : ( n13356 ) ;
assign n13358 =  ( n12855 ) ? ( VREG_15_11 ) : ( n13357 ) ;
assign n13359 =  ( n12854 ) ? ( VREG_15_12 ) : ( n13358 ) ;
assign n13360 =  ( n12853 ) ? ( VREG_15_13 ) : ( n13359 ) ;
assign n13361 =  ( n12852 ) ? ( VREG_15_14 ) : ( n13360 ) ;
assign n13362 =  ( n12851 ) ? ( VREG_15_15 ) : ( n13361 ) ;
assign n13363 =  ( n12850 ) ? ( VREG_16_0 ) : ( n13362 ) ;
assign n13364 =  ( n12849 ) ? ( VREG_16_1 ) : ( n13363 ) ;
assign n13365 =  ( n12848 ) ? ( VREG_16_2 ) : ( n13364 ) ;
assign n13366 =  ( n12847 ) ? ( VREG_16_3 ) : ( n13365 ) ;
assign n13367 =  ( n12846 ) ? ( VREG_16_4 ) : ( n13366 ) ;
assign n13368 =  ( n12845 ) ? ( VREG_16_5 ) : ( n13367 ) ;
assign n13369 =  ( n12844 ) ? ( VREG_16_6 ) : ( n13368 ) ;
assign n13370 =  ( n12843 ) ? ( VREG_16_7 ) : ( n13369 ) ;
assign n13371 =  ( n12842 ) ? ( VREG_16_8 ) : ( n13370 ) ;
assign n13372 =  ( n12841 ) ? ( VREG_16_9 ) : ( n13371 ) ;
assign n13373 =  ( n12840 ) ? ( VREG_16_10 ) : ( n13372 ) ;
assign n13374 =  ( n12839 ) ? ( VREG_16_11 ) : ( n13373 ) ;
assign n13375 =  ( n12838 ) ? ( VREG_16_12 ) : ( n13374 ) ;
assign n13376 =  ( n12837 ) ? ( VREG_16_13 ) : ( n13375 ) ;
assign n13377 =  ( n12836 ) ? ( VREG_16_14 ) : ( n13376 ) ;
assign n13378 =  ( n12835 ) ? ( VREG_16_15 ) : ( n13377 ) ;
assign n13379 =  ( n12834 ) ? ( VREG_17_0 ) : ( n13378 ) ;
assign n13380 =  ( n12833 ) ? ( VREG_17_1 ) : ( n13379 ) ;
assign n13381 =  ( n12832 ) ? ( VREG_17_2 ) : ( n13380 ) ;
assign n13382 =  ( n12831 ) ? ( VREG_17_3 ) : ( n13381 ) ;
assign n13383 =  ( n12830 ) ? ( VREG_17_4 ) : ( n13382 ) ;
assign n13384 =  ( n12829 ) ? ( VREG_17_5 ) : ( n13383 ) ;
assign n13385 =  ( n12828 ) ? ( VREG_17_6 ) : ( n13384 ) ;
assign n13386 =  ( n12827 ) ? ( VREG_17_7 ) : ( n13385 ) ;
assign n13387 =  ( n12826 ) ? ( VREG_17_8 ) : ( n13386 ) ;
assign n13388 =  ( n12825 ) ? ( VREG_17_9 ) : ( n13387 ) ;
assign n13389 =  ( n12824 ) ? ( VREG_17_10 ) : ( n13388 ) ;
assign n13390 =  ( n12823 ) ? ( VREG_17_11 ) : ( n13389 ) ;
assign n13391 =  ( n12822 ) ? ( VREG_17_12 ) : ( n13390 ) ;
assign n13392 =  ( n12821 ) ? ( VREG_17_13 ) : ( n13391 ) ;
assign n13393 =  ( n12820 ) ? ( VREG_17_14 ) : ( n13392 ) ;
assign n13394 =  ( n12819 ) ? ( VREG_17_15 ) : ( n13393 ) ;
assign n13395 =  ( n12818 ) ? ( VREG_18_0 ) : ( n13394 ) ;
assign n13396 =  ( n12817 ) ? ( VREG_18_1 ) : ( n13395 ) ;
assign n13397 =  ( n12816 ) ? ( VREG_18_2 ) : ( n13396 ) ;
assign n13398 =  ( n12815 ) ? ( VREG_18_3 ) : ( n13397 ) ;
assign n13399 =  ( n12814 ) ? ( VREG_18_4 ) : ( n13398 ) ;
assign n13400 =  ( n12813 ) ? ( VREG_18_5 ) : ( n13399 ) ;
assign n13401 =  ( n12812 ) ? ( VREG_18_6 ) : ( n13400 ) ;
assign n13402 =  ( n12811 ) ? ( VREG_18_7 ) : ( n13401 ) ;
assign n13403 =  ( n12810 ) ? ( VREG_18_8 ) : ( n13402 ) ;
assign n13404 =  ( n12809 ) ? ( VREG_18_9 ) : ( n13403 ) ;
assign n13405 =  ( n12808 ) ? ( VREG_18_10 ) : ( n13404 ) ;
assign n13406 =  ( n12807 ) ? ( VREG_18_11 ) : ( n13405 ) ;
assign n13407 =  ( n12806 ) ? ( VREG_18_12 ) : ( n13406 ) ;
assign n13408 =  ( n12805 ) ? ( VREG_18_13 ) : ( n13407 ) ;
assign n13409 =  ( n12804 ) ? ( VREG_18_14 ) : ( n13408 ) ;
assign n13410 =  ( n12803 ) ? ( VREG_18_15 ) : ( n13409 ) ;
assign n13411 =  ( n12802 ) ? ( VREG_19_0 ) : ( n13410 ) ;
assign n13412 =  ( n12801 ) ? ( VREG_19_1 ) : ( n13411 ) ;
assign n13413 =  ( n12800 ) ? ( VREG_19_2 ) : ( n13412 ) ;
assign n13414 =  ( n12799 ) ? ( VREG_19_3 ) : ( n13413 ) ;
assign n13415 =  ( n12798 ) ? ( VREG_19_4 ) : ( n13414 ) ;
assign n13416 =  ( n12797 ) ? ( VREG_19_5 ) : ( n13415 ) ;
assign n13417 =  ( n12796 ) ? ( VREG_19_6 ) : ( n13416 ) ;
assign n13418 =  ( n12795 ) ? ( VREG_19_7 ) : ( n13417 ) ;
assign n13419 =  ( n12794 ) ? ( VREG_19_8 ) : ( n13418 ) ;
assign n13420 =  ( n12793 ) ? ( VREG_19_9 ) : ( n13419 ) ;
assign n13421 =  ( n12792 ) ? ( VREG_19_10 ) : ( n13420 ) ;
assign n13422 =  ( n12791 ) ? ( VREG_19_11 ) : ( n13421 ) ;
assign n13423 =  ( n12790 ) ? ( VREG_19_12 ) : ( n13422 ) ;
assign n13424 =  ( n12789 ) ? ( VREG_19_13 ) : ( n13423 ) ;
assign n13425 =  ( n12788 ) ? ( VREG_19_14 ) : ( n13424 ) ;
assign n13426 =  ( n12787 ) ? ( VREG_19_15 ) : ( n13425 ) ;
assign n13427 =  ( n12786 ) ? ( VREG_20_0 ) : ( n13426 ) ;
assign n13428 =  ( n12785 ) ? ( VREG_20_1 ) : ( n13427 ) ;
assign n13429 =  ( n12784 ) ? ( VREG_20_2 ) : ( n13428 ) ;
assign n13430 =  ( n12783 ) ? ( VREG_20_3 ) : ( n13429 ) ;
assign n13431 =  ( n12782 ) ? ( VREG_20_4 ) : ( n13430 ) ;
assign n13432 =  ( n12781 ) ? ( VREG_20_5 ) : ( n13431 ) ;
assign n13433 =  ( n12780 ) ? ( VREG_20_6 ) : ( n13432 ) ;
assign n13434 =  ( n12779 ) ? ( VREG_20_7 ) : ( n13433 ) ;
assign n13435 =  ( n12778 ) ? ( VREG_20_8 ) : ( n13434 ) ;
assign n13436 =  ( n12777 ) ? ( VREG_20_9 ) : ( n13435 ) ;
assign n13437 =  ( n12776 ) ? ( VREG_20_10 ) : ( n13436 ) ;
assign n13438 =  ( n12775 ) ? ( VREG_20_11 ) : ( n13437 ) ;
assign n13439 =  ( n12774 ) ? ( VREG_20_12 ) : ( n13438 ) ;
assign n13440 =  ( n12773 ) ? ( VREG_20_13 ) : ( n13439 ) ;
assign n13441 =  ( n12772 ) ? ( VREG_20_14 ) : ( n13440 ) ;
assign n13442 =  ( n12771 ) ? ( VREG_20_15 ) : ( n13441 ) ;
assign n13443 =  ( n12770 ) ? ( VREG_21_0 ) : ( n13442 ) ;
assign n13444 =  ( n12769 ) ? ( VREG_21_1 ) : ( n13443 ) ;
assign n13445 =  ( n12768 ) ? ( VREG_21_2 ) : ( n13444 ) ;
assign n13446 =  ( n12767 ) ? ( VREG_21_3 ) : ( n13445 ) ;
assign n13447 =  ( n12766 ) ? ( VREG_21_4 ) : ( n13446 ) ;
assign n13448 =  ( n12765 ) ? ( VREG_21_5 ) : ( n13447 ) ;
assign n13449 =  ( n12764 ) ? ( VREG_21_6 ) : ( n13448 ) ;
assign n13450 =  ( n12763 ) ? ( VREG_21_7 ) : ( n13449 ) ;
assign n13451 =  ( n12762 ) ? ( VREG_21_8 ) : ( n13450 ) ;
assign n13452 =  ( n12761 ) ? ( VREG_21_9 ) : ( n13451 ) ;
assign n13453 =  ( n12760 ) ? ( VREG_21_10 ) : ( n13452 ) ;
assign n13454 =  ( n12759 ) ? ( VREG_21_11 ) : ( n13453 ) ;
assign n13455 =  ( n12758 ) ? ( VREG_21_12 ) : ( n13454 ) ;
assign n13456 =  ( n12757 ) ? ( VREG_21_13 ) : ( n13455 ) ;
assign n13457 =  ( n12756 ) ? ( VREG_21_14 ) : ( n13456 ) ;
assign n13458 =  ( n12755 ) ? ( VREG_21_15 ) : ( n13457 ) ;
assign n13459 =  ( n12754 ) ? ( VREG_22_0 ) : ( n13458 ) ;
assign n13460 =  ( n12753 ) ? ( VREG_22_1 ) : ( n13459 ) ;
assign n13461 =  ( n12752 ) ? ( VREG_22_2 ) : ( n13460 ) ;
assign n13462 =  ( n12751 ) ? ( VREG_22_3 ) : ( n13461 ) ;
assign n13463 =  ( n12750 ) ? ( VREG_22_4 ) : ( n13462 ) ;
assign n13464 =  ( n12749 ) ? ( VREG_22_5 ) : ( n13463 ) ;
assign n13465 =  ( n12748 ) ? ( VREG_22_6 ) : ( n13464 ) ;
assign n13466 =  ( n12747 ) ? ( VREG_22_7 ) : ( n13465 ) ;
assign n13467 =  ( n12746 ) ? ( VREG_22_8 ) : ( n13466 ) ;
assign n13468 =  ( n12745 ) ? ( VREG_22_9 ) : ( n13467 ) ;
assign n13469 =  ( n12744 ) ? ( VREG_22_10 ) : ( n13468 ) ;
assign n13470 =  ( n12743 ) ? ( VREG_22_11 ) : ( n13469 ) ;
assign n13471 =  ( n12742 ) ? ( VREG_22_12 ) : ( n13470 ) ;
assign n13472 =  ( n12741 ) ? ( VREG_22_13 ) : ( n13471 ) ;
assign n13473 =  ( n12740 ) ? ( VREG_22_14 ) : ( n13472 ) ;
assign n13474 =  ( n12739 ) ? ( VREG_22_15 ) : ( n13473 ) ;
assign n13475 =  ( n12738 ) ? ( VREG_23_0 ) : ( n13474 ) ;
assign n13476 =  ( n12737 ) ? ( VREG_23_1 ) : ( n13475 ) ;
assign n13477 =  ( n12736 ) ? ( VREG_23_2 ) : ( n13476 ) ;
assign n13478 =  ( n12735 ) ? ( VREG_23_3 ) : ( n13477 ) ;
assign n13479 =  ( n12734 ) ? ( VREG_23_4 ) : ( n13478 ) ;
assign n13480 =  ( n12733 ) ? ( VREG_23_5 ) : ( n13479 ) ;
assign n13481 =  ( n12732 ) ? ( VREG_23_6 ) : ( n13480 ) ;
assign n13482 =  ( n12731 ) ? ( VREG_23_7 ) : ( n13481 ) ;
assign n13483 =  ( n12730 ) ? ( VREG_23_8 ) : ( n13482 ) ;
assign n13484 =  ( n12729 ) ? ( VREG_23_9 ) : ( n13483 ) ;
assign n13485 =  ( n12728 ) ? ( VREG_23_10 ) : ( n13484 ) ;
assign n13486 =  ( n12727 ) ? ( VREG_23_11 ) : ( n13485 ) ;
assign n13487 =  ( n12726 ) ? ( VREG_23_12 ) : ( n13486 ) ;
assign n13488 =  ( n12725 ) ? ( VREG_23_13 ) : ( n13487 ) ;
assign n13489 =  ( n12724 ) ? ( VREG_23_14 ) : ( n13488 ) ;
assign n13490 =  ( n12723 ) ? ( VREG_23_15 ) : ( n13489 ) ;
assign n13491 =  ( n12722 ) ? ( VREG_24_0 ) : ( n13490 ) ;
assign n13492 =  ( n12721 ) ? ( VREG_24_1 ) : ( n13491 ) ;
assign n13493 =  ( n12720 ) ? ( VREG_24_2 ) : ( n13492 ) ;
assign n13494 =  ( n12719 ) ? ( VREG_24_3 ) : ( n13493 ) ;
assign n13495 =  ( n12718 ) ? ( VREG_24_4 ) : ( n13494 ) ;
assign n13496 =  ( n12717 ) ? ( VREG_24_5 ) : ( n13495 ) ;
assign n13497 =  ( n12716 ) ? ( VREG_24_6 ) : ( n13496 ) ;
assign n13498 =  ( n12715 ) ? ( VREG_24_7 ) : ( n13497 ) ;
assign n13499 =  ( n12714 ) ? ( VREG_24_8 ) : ( n13498 ) ;
assign n13500 =  ( n12713 ) ? ( VREG_24_9 ) : ( n13499 ) ;
assign n13501 =  ( n12712 ) ? ( VREG_24_10 ) : ( n13500 ) ;
assign n13502 =  ( n12711 ) ? ( VREG_24_11 ) : ( n13501 ) ;
assign n13503 =  ( n12710 ) ? ( VREG_24_12 ) : ( n13502 ) ;
assign n13504 =  ( n12709 ) ? ( VREG_24_13 ) : ( n13503 ) ;
assign n13505 =  ( n12708 ) ? ( VREG_24_14 ) : ( n13504 ) ;
assign n13506 =  ( n12707 ) ? ( VREG_24_15 ) : ( n13505 ) ;
assign n13507 =  ( n12706 ) ? ( VREG_25_0 ) : ( n13506 ) ;
assign n13508 =  ( n12705 ) ? ( VREG_25_1 ) : ( n13507 ) ;
assign n13509 =  ( n12704 ) ? ( VREG_25_2 ) : ( n13508 ) ;
assign n13510 =  ( n12703 ) ? ( VREG_25_3 ) : ( n13509 ) ;
assign n13511 =  ( n12702 ) ? ( VREG_25_4 ) : ( n13510 ) ;
assign n13512 =  ( n12701 ) ? ( VREG_25_5 ) : ( n13511 ) ;
assign n13513 =  ( n12700 ) ? ( VREG_25_6 ) : ( n13512 ) ;
assign n13514 =  ( n12699 ) ? ( VREG_25_7 ) : ( n13513 ) ;
assign n13515 =  ( n12698 ) ? ( VREG_25_8 ) : ( n13514 ) ;
assign n13516 =  ( n12697 ) ? ( VREG_25_9 ) : ( n13515 ) ;
assign n13517 =  ( n12696 ) ? ( VREG_25_10 ) : ( n13516 ) ;
assign n13518 =  ( n12695 ) ? ( VREG_25_11 ) : ( n13517 ) ;
assign n13519 =  ( n12694 ) ? ( VREG_25_12 ) : ( n13518 ) ;
assign n13520 =  ( n12693 ) ? ( VREG_25_13 ) : ( n13519 ) ;
assign n13521 =  ( n12692 ) ? ( VREG_25_14 ) : ( n13520 ) ;
assign n13522 =  ( n12691 ) ? ( VREG_25_15 ) : ( n13521 ) ;
assign n13523 =  ( n12690 ) ? ( VREG_26_0 ) : ( n13522 ) ;
assign n13524 =  ( n12689 ) ? ( VREG_26_1 ) : ( n13523 ) ;
assign n13525 =  ( n12688 ) ? ( VREG_26_2 ) : ( n13524 ) ;
assign n13526 =  ( n12687 ) ? ( VREG_26_3 ) : ( n13525 ) ;
assign n13527 =  ( n12686 ) ? ( VREG_26_4 ) : ( n13526 ) ;
assign n13528 =  ( n12685 ) ? ( VREG_26_5 ) : ( n13527 ) ;
assign n13529 =  ( n12684 ) ? ( VREG_26_6 ) : ( n13528 ) ;
assign n13530 =  ( n12683 ) ? ( VREG_26_7 ) : ( n13529 ) ;
assign n13531 =  ( n12682 ) ? ( VREG_26_8 ) : ( n13530 ) ;
assign n13532 =  ( n12681 ) ? ( VREG_26_9 ) : ( n13531 ) ;
assign n13533 =  ( n12680 ) ? ( VREG_26_10 ) : ( n13532 ) ;
assign n13534 =  ( n12679 ) ? ( VREG_26_11 ) : ( n13533 ) ;
assign n13535 =  ( n12678 ) ? ( VREG_26_12 ) : ( n13534 ) ;
assign n13536 =  ( n12677 ) ? ( VREG_26_13 ) : ( n13535 ) ;
assign n13537 =  ( n12676 ) ? ( VREG_26_14 ) : ( n13536 ) ;
assign n13538 =  ( n12675 ) ? ( VREG_26_15 ) : ( n13537 ) ;
assign n13539 =  ( n12674 ) ? ( VREG_27_0 ) : ( n13538 ) ;
assign n13540 =  ( n12673 ) ? ( VREG_27_1 ) : ( n13539 ) ;
assign n13541 =  ( n12672 ) ? ( VREG_27_2 ) : ( n13540 ) ;
assign n13542 =  ( n12671 ) ? ( VREG_27_3 ) : ( n13541 ) ;
assign n13543 =  ( n12670 ) ? ( VREG_27_4 ) : ( n13542 ) ;
assign n13544 =  ( n12669 ) ? ( VREG_27_5 ) : ( n13543 ) ;
assign n13545 =  ( n12668 ) ? ( VREG_27_6 ) : ( n13544 ) ;
assign n13546 =  ( n12667 ) ? ( VREG_27_7 ) : ( n13545 ) ;
assign n13547 =  ( n12666 ) ? ( VREG_27_8 ) : ( n13546 ) ;
assign n13548 =  ( n12665 ) ? ( VREG_27_9 ) : ( n13547 ) ;
assign n13549 =  ( n12664 ) ? ( VREG_27_10 ) : ( n13548 ) ;
assign n13550 =  ( n12663 ) ? ( VREG_27_11 ) : ( n13549 ) ;
assign n13551 =  ( n12662 ) ? ( VREG_27_12 ) : ( n13550 ) ;
assign n13552 =  ( n12661 ) ? ( VREG_27_13 ) : ( n13551 ) ;
assign n13553 =  ( n12660 ) ? ( VREG_27_14 ) : ( n13552 ) ;
assign n13554 =  ( n12659 ) ? ( VREG_27_15 ) : ( n13553 ) ;
assign n13555 =  ( n12658 ) ? ( VREG_28_0 ) : ( n13554 ) ;
assign n13556 =  ( n12657 ) ? ( VREG_28_1 ) : ( n13555 ) ;
assign n13557 =  ( n12656 ) ? ( VREG_28_2 ) : ( n13556 ) ;
assign n13558 =  ( n12655 ) ? ( VREG_28_3 ) : ( n13557 ) ;
assign n13559 =  ( n12654 ) ? ( VREG_28_4 ) : ( n13558 ) ;
assign n13560 =  ( n12653 ) ? ( VREG_28_5 ) : ( n13559 ) ;
assign n13561 =  ( n12652 ) ? ( VREG_28_6 ) : ( n13560 ) ;
assign n13562 =  ( n12651 ) ? ( VREG_28_7 ) : ( n13561 ) ;
assign n13563 =  ( n12650 ) ? ( VREG_28_8 ) : ( n13562 ) ;
assign n13564 =  ( n12649 ) ? ( VREG_28_9 ) : ( n13563 ) ;
assign n13565 =  ( n12648 ) ? ( VREG_28_10 ) : ( n13564 ) ;
assign n13566 =  ( n12647 ) ? ( VREG_28_11 ) : ( n13565 ) ;
assign n13567 =  ( n12646 ) ? ( VREG_28_12 ) : ( n13566 ) ;
assign n13568 =  ( n12645 ) ? ( VREG_28_13 ) : ( n13567 ) ;
assign n13569 =  ( n12644 ) ? ( VREG_28_14 ) : ( n13568 ) ;
assign n13570 =  ( n12643 ) ? ( VREG_28_15 ) : ( n13569 ) ;
assign n13571 =  ( n12642 ) ? ( VREG_29_0 ) : ( n13570 ) ;
assign n13572 =  ( n12641 ) ? ( VREG_29_1 ) : ( n13571 ) ;
assign n13573 =  ( n12640 ) ? ( VREG_29_2 ) : ( n13572 ) ;
assign n13574 =  ( n12639 ) ? ( VREG_29_3 ) : ( n13573 ) ;
assign n13575 =  ( n12638 ) ? ( VREG_29_4 ) : ( n13574 ) ;
assign n13576 =  ( n12637 ) ? ( VREG_29_5 ) : ( n13575 ) ;
assign n13577 =  ( n12636 ) ? ( VREG_29_6 ) : ( n13576 ) ;
assign n13578 =  ( n12635 ) ? ( VREG_29_7 ) : ( n13577 ) ;
assign n13579 =  ( n12634 ) ? ( VREG_29_8 ) : ( n13578 ) ;
assign n13580 =  ( n12633 ) ? ( VREG_29_9 ) : ( n13579 ) ;
assign n13581 =  ( n12632 ) ? ( VREG_29_10 ) : ( n13580 ) ;
assign n13582 =  ( n12631 ) ? ( VREG_29_11 ) : ( n13581 ) ;
assign n13583 =  ( n12630 ) ? ( VREG_29_12 ) : ( n13582 ) ;
assign n13584 =  ( n12629 ) ? ( VREG_29_13 ) : ( n13583 ) ;
assign n13585 =  ( n12628 ) ? ( VREG_29_14 ) : ( n13584 ) ;
assign n13586 =  ( n12627 ) ? ( VREG_29_15 ) : ( n13585 ) ;
assign n13587 =  ( n12626 ) ? ( VREG_30_0 ) : ( n13586 ) ;
assign n13588 =  ( n12625 ) ? ( VREG_30_1 ) : ( n13587 ) ;
assign n13589 =  ( n12624 ) ? ( VREG_30_2 ) : ( n13588 ) ;
assign n13590 =  ( n12623 ) ? ( VREG_30_3 ) : ( n13589 ) ;
assign n13591 =  ( n12622 ) ? ( VREG_30_4 ) : ( n13590 ) ;
assign n13592 =  ( n12621 ) ? ( VREG_30_5 ) : ( n13591 ) ;
assign n13593 =  ( n12620 ) ? ( VREG_30_6 ) : ( n13592 ) ;
assign n13594 =  ( n12619 ) ? ( VREG_30_7 ) : ( n13593 ) ;
assign n13595 =  ( n12618 ) ? ( VREG_30_8 ) : ( n13594 ) ;
assign n13596 =  ( n12617 ) ? ( VREG_30_9 ) : ( n13595 ) ;
assign n13597 =  ( n12616 ) ? ( VREG_30_10 ) : ( n13596 ) ;
assign n13598 =  ( n12615 ) ? ( VREG_30_11 ) : ( n13597 ) ;
assign n13599 =  ( n12614 ) ? ( VREG_30_12 ) : ( n13598 ) ;
assign n13600 =  ( n12613 ) ? ( VREG_30_13 ) : ( n13599 ) ;
assign n13601 =  ( n12612 ) ? ( VREG_30_14 ) : ( n13600 ) ;
assign n13602 =  ( n12611 ) ? ( VREG_30_15 ) : ( n13601 ) ;
assign n13603 =  ( n12610 ) ? ( VREG_31_0 ) : ( n13602 ) ;
assign n13604 =  ( n12609 ) ? ( VREG_31_1 ) : ( n13603 ) ;
assign n13605 =  ( n12608 ) ? ( VREG_31_2 ) : ( n13604 ) ;
assign n13606 =  ( n12607 ) ? ( VREG_31_3 ) : ( n13605 ) ;
assign n13607 =  ( n12606 ) ? ( VREG_31_4 ) : ( n13606 ) ;
assign n13608 =  ( n12605 ) ? ( VREG_31_5 ) : ( n13607 ) ;
assign n13609 =  ( n12604 ) ? ( VREG_31_6 ) : ( n13608 ) ;
assign n13610 =  ( n12603 ) ? ( VREG_31_7 ) : ( n13609 ) ;
assign n13611 =  ( n12602 ) ? ( VREG_31_8 ) : ( n13610 ) ;
assign n13612 =  ( n12601 ) ? ( VREG_31_9 ) : ( n13611 ) ;
assign n13613 =  ( n12600 ) ? ( VREG_31_10 ) : ( n13612 ) ;
assign n13614 =  ( n12599 ) ? ( VREG_31_11 ) : ( n13613 ) ;
assign n13615 =  ( n12598 ) ? ( VREG_31_12 ) : ( n13614 ) ;
assign n13616 =  ( n12597 ) ? ( VREG_31_13 ) : ( n13615 ) ;
assign n13617 =  ( n12596 ) ? ( VREG_31_14 ) : ( n13616 ) ;
assign n13618 =  ( n12595 ) ? ( VREG_31_15 ) : ( n13617 ) ;
assign n13619 =  ( n12584 ) + ( n13618 )  ;
assign n13620 =  ( n12584 ) - ( n13618 )  ;
assign n13621 =  ( n12584 ) & ( n13618 )  ;
assign n13622 =  ( n12584 ) | ( n13618 )  ;
assign n13623 =  ( ( n12584 ) * ( n13618 ))  ;
assign n13624 =  ( n148 ) ? ( n13623 ) : ( VREG_0_13 ) ;
assign n13625 =  ( n146 ) ? ( n13622 ) : ( n13624 ) ;
assign n13626 =  ( n144 ) ? ( n13621 ) : ( n13625 ) ;
assign n13627 =  ( n142 ) ? ( n13620 ) : ( n13626 ) ;
assign n13628 =  ( n10 ) ? ( n13619 ) : ( n13627 ) ;
assign n13629 = n3030[13:13] ;
assign n13630 =  ( n13629 ) == ( 1'd0 )  ;
assign n13631 =  ( n13630 ) ? ( VREG_0_13 ) : ( n12594 ) ;
assign n13632 =  ( n13630 ) ? ( VREG_0_13 ) : ( n13628 ) ;
assign n13633 =  ( n3034 ) ? ( n13632 ) : ( VREG_0_13 ) ;
assign n13634 =  ( n2965 ) ? ( n13631 ) : ( n13633 ) ;
assign n13635 =  ( n1930 ) ? ( n13628 ) : ( n13634 ) ;
assign n13636 =  ( n879 ) ? ( n12594 ) : ( n13635 ) ;
assign n13637 =  ( n12584 ) + ( n164 )  ;
assign n13638 =  ( n12584 ) - ( n164 )  ;
assign n13639 =  ( n12584 ) & ( n164 )  ;
assign n13640 =  ( n12584 ) | ( n164 )  ;
assign n13641 =  ( ( n12584 ) * ( n164 ))  ;
assign n13642 =  ( n172 ) ? ( n13641 ) : ( VREG_0_13 ) ;
assign n13643 =  ( n170 ) ? ( n13640 ) : ( n13642 ) ;
assign n13644 =  ( n168 ) ? ( n13639 ) : ( n13643 ) ;
assign n13645 =  ( n166 ) ? ( n13638 ) : ( n13644 ) ;
assign n13646 =  ( n162 ) ? ( n13637 ) : ( n13645 ) ;
assign n13647 =  ( n12584 ) + ( n180 )  ;
assign n13648 =  ( n12584 ) - ( n180 )  ;
assign n13649 =  ( n12584 ) & ( n180 )  ;
assign n13650 =  ( n12584 ) | ( n180 )  ;
assign n13651 =  ( ( n12584 ) * ( n180 ))  ;
assign n13652 =  ( n172 ) ? ( n13651 ) : ( VREG_0_13 ) ;
assign n13653 =  ( n170 ) ? ( n13650 ) : ( n13652 ) ;
assign n13654 =  ( n168 ) ? ( n13649 ) : ( n13653 ) ;
assign n13655 =  ( n166 ) ? ( n13648 ) : ( n13654 ) ;
assign n13656 =  ( n162 ) ? ( n13647 ) : ( n13655 ) ;
assign n13657 =  ( n13630 ) ? ( VREG_0_13 ) : ( n13656 ) ;
assign n13658 =  ( n3051 ) ? ( n13657 ) : ( VREG_0_13 ) ;
assign n13659 =  ( n3040 ) ? ( n13646 ) : ( n13658 ) ;
assign n13660 =  ( n192 ) ? ( VREG_0_13 ) : ( VREG_0_13 ) ;
assign n13661 =  ( n157 ) ? ( n13659 ) : ( n13660 ) ;
assign n13662 =  ( n6 ) ? ( n13636 ) : ( n13661 ) ;
assign n13663 =  ( n4 ) ? ( n13662 ) : ( VREG_0_13 ) ;
assign n13664 =  ( 32'd14 ) == ( 32'd15 )  ;
assign n13665 =  ( n12 ) & ( n13664 )  ;
assign n13666 =  ( 32'd14 ) == ( 32'd14 )  ;
assign n13667 =  ( n12 ) & ( n13666 )  ;
assign n13668 =  ( 32'd14 ) == ( 32'd13 )  ;
assign n13669 =  ( n12 ) & ( n13668 )  ;
assign n13670 =  ( 32'd14 ) == ( 32'd12 )  ;
assign n13671 =  ( n12 ) & ( n13670 )  ;
assign n13672 =  ( 32'd14 ) == ( 32'd11 )  ;
assign n13673 =  ( n12 ) & ( n13672 )  ;
assign n13674 =  ( 32'd14 ) == ( 32'd10 )  ;
assign n13675 =  ( n12 ) & ( n13674 )  ;
assign n13676 =  ( 32'd14 ) == ( 32'd9 )  ;
assign n13677 =  ( n12 ) & ( n13676 )  ;
assign n13678 =  ( 32'd14 ) == ( 32'd8 )  ;
assign n13679 =  ( n12 ) & ( n13678 )  ;
assign n13680 =  ( 32'd14 ) == ( 32'd7 )  ;
assign n13681 =  ( n12 ) & ( n13680 )  ;
assign n13682 =  ( 32'd14 ) == ( 32'd6 )  ;
assign n13683 =  ( n12 ) & ( n13682 )  ;
assign n13684 =  ( 32'd14 ) == ( 32'd5 )  ;
assign n13685 =  ( n12 ) & ( n13684 )  ;
assign n13686 =  ( 32'd14 ) == ( 32'd4 )  ;
assign n13687 =  ( n12 ) & ( n13686 )  ;
assign n13688 =  ( 32'd14 ) == ( 32'd3 )  ;
assign n13689 =  ( n12 ) & ( n13688 )  ;
assign n13690 =  ( 32'd14 ) == ( 32'd2 )  ;
assign n13691 =  ( n12 ) & ( n13690 )  ;
assign n13692 =  ( 32'd14 ) == ( 32'd1 )  ;
assign n13693 =  ( n12 ) & ( n13692 )  ;
assign n13694 =  ( 32'd14 ) == ( 32'd0 )  ;
assign n13695 =  ( n12 ) & ( n13694 )  ;
assign n13696 =  ( n13 ) & ( n13664 )  ;
assign n13697 =  ( n13 ) & ( n13666 )  ;
assign n13698 =  ( n13 ) & ( n13668 )  ;
assign n13699 =  ( n13 ) & ( n13670 )  ;
assign n13700 =  ( n13 ) & ( n13672 )  ;
assign n13701 =  ( n13 ) & ( n13674 )  ;
assign n13702 =  ( n13 ) & ( n13676 )  ;
assign n13703 =  ( n13 ) & ( n13678 )  ;
assign n13704 =  ( n13 ) & ( n13680 )  ;
assign n13705 =  ( n13 ) & ( n13682 )  ;
assign n13706 =  ( n13 ) & ( n13684 )  ;
assign n13707 =  ( n13 ) & ( n13686 )  ;
assign n13708 =  ( n13 ) & ( n13688 )  ;
assign n13709 =  ( n13 ) & ( n13690 )  ;
assign n13710 =  ( n13 ) & ( n13692 )  ;
assign n13711 =  ( n13 ) & ( n13694 )  ;
assign n13712 =  ( n14 ) & ( n13664 )  ;
assign n13713 =  ( n14 ) & ( n13666 )  ;
assign n13714 =  ( n14 ) & ( n13668 )  ;
assign n13715 =  ( n14 ) & ( n13670 )  ;
assign n13716 =  ( n14 ) & ( n13672 )  ;
assign n13717 =  ( n14 ) & ( n13674 )  ;
assign n13718 =  ( n14 ) & ( n13676 )  ;
assign n13719 =  ( n14 ) & ( n13678 )  ;
assign n13720 =  ( n14 ) & ( n13680 )  ;
assign n13721 =  ( n14 ) & ( n13682 )  ;
assign n13722 =  ( n14 ) & ( n13684 )  ;
assign n13723 =  ( n14 ) & ( n13686 )  ;
assign n13724 =  ( n14 ) & ( n13688 )  ;
assign n13725 =  ( n14 ) & ( n13690 )  ;
assign n13726 =  ( n14 ) & ( n13692 )  ;
assign n13727 =  ( n14 ) & ( n13694 )  ;
assign n13728 =  ( n15 ) & ( n13664 )  ;
assign n13729 =  ( n15 ) & ( n13666 )  ;
assign n13730 =  ( n15 ) & ( n13668 )  ;
assign n13731 =  ( n15 ) & ( n13670 )  ;
assign n13732 =  ( n15 ) & ( n13672 )  ;
assign n13733 =  ( n15 ) & ( n13674 )  ;
assign n13734 =  ( n15 ) & ( n13676 )  ;
assign n13735 =  ( n15 ) & ( n13678 )  ;
assign n13736 =  ( n15 ) & ( n13680 )  ;
assign n13737 =  ( n15 ) & ( n13682 )  ;
assign n13738 =  ( n15 ) & ( n13684 )  ;
assign n13739 =  ( n15 ) & ( n13686 )  ;
assign n13740 =  ( n15 ) & ( n13688 )  ;
assign n13741 =  ( n15 ) & ( n13690 )  ;
assign n13742 =  ( n15 ) & ( n13692 )  ;
assign n13743 =  ( n15 ) & ( n13694 )  ;
assign n13744 =  ( n16 ) & ( n13664 )  ;
assign n13745 =  ( n16 ) & ( n13666 )  ;
assign n13746 =  ( n16 ) & ( n13668 )  ;
assign n13747 =  ( n16 ) & ( n13670 )  ;
assign n13748 =  ( n16 ) & ( n13672 )  ;
assign n13749 =  ( n16 ) & ( n13674 )  ;
assign n13750 =  ( n16 ) & ( n13676 )  ;
assign n13751 =  ( n16 ) & ( n13678 )  ;
assign n13752 =  ( n16 ) & ( n13680 )  ;
assign n13753 =  ( n16 ) & ( n13682 )  ;
assign n13754 =  ( n16 ) & ( n13684 )  ;
assign n13755 =  ( n16 ) & ( n13686 )  ;
assign n13756 =  ( n16 ) & ( n13688 )  ;
assign n13757 =  ( n16 ) & ( n13690 )  ;
assign n13758 =  ( n16 ) & ( n13692 )  ;
assign n13759 =  ( n16 ) & ( n13694 )  ;
assign n13760 =  ( n17 ) & ( n13664 )  ;
assign n13761 =  ( n17 ) & ( n13666 )  ;
assign n13762 =  ( n17 ) & ( n13668 )  ;
assign n13763 =  ( n17 ) & ( n13670 )  ;
assign n13764 =  ( n17 ) & ( n13672 )  ;
assign n13765 =  ( n17 ) & ( n13674 )  ;
assign n13766 =  ( n17 ) & ( n13676 )  ;
assign n13767 =  ( n17 ) & ( n13678 )  ;
assign n13768 =  ( n17 ) & ( n13680 )  ;
assign n13769 =  ( n17 ) & ( n13682 )  ;
assign n13770 =  ( n17 ) & ( n13684 )  ;
assign n13771 =  ( n17 ) & ( n13686 )  ;
assign n13772 =  ( n17 ) & ( n13688 )  ;
assign n13773 =  ( n17 ) & ( n13690 )  ;
assign n13774 =  ( n17 ) & ( n13692 )  ;
assign n13775 =  ( n17 ) & ( n13694 )  ;
assign n13776 =  ( n18 ) & ( n13664 )  ;
assign n13777 =  ( n18 ) & ( n13666 )  ;
assign n13778 =  ( n18 ) & ( n13668 )  ;
assign n13779 =  ( n18 ) & ( n13670 )  ;
assign n13780 =  ( n18 ) & ( n13672 )  ;
assign n13781 =  ( n18 ) & ( n13674 )  ;
assign n13782 =  ( n18 ) & ( n13676 )  ;
assign n13783 =  ( n18 ) & ( n13678 )  ;
assign n13784 =  ( n18 ) & ( n13680 )  ;
assign n13785 =  ( n18 ) & ( n13682 )  ;
assign n13786 =  ( n18 ) & ( n13684 )  ;
assign n13787 =  ( n18 ) & ( n13686 )  ;
assign n13788 =  ( n18 ) & ( n13688 )  ;
assign n13789 =  ( n18 ) & ( n13690 )  ;
assign n13790 =  ( n18 ) & ( n13692 )  ;
assign n13791 =  ( n18 ) & ( n13694 )  ;
assign n13792 =  ( n19 ) & ( n13664 )  ;
assign n13793 =  ( n19 ) & ( n13666 )  ;
assign n13794 =  ( n19 ) & ( n13668 )  ;
assign n13795 =  ( n19 ) & ( n13670 )  ;
assign n13796 =  ( n19 ) & ( n13672 )  ;
assign n13797 =  ( n19 ) & ( n13674 )  ;
assign n13798 =  ( n19 ) & ( n13676 )  ;
assign n13799 =  ( n19 ) & ( n13678 )  ;
assign n13800 =  ( n19 ) & ( n13680 )  ;
assign n13801 =  ( n19 ) & ( n13682 )  ;
assign n13802 =  ( n19 ) & ( n13684 )  ;
assign n13803 =  ( n19 ) & ( n13686 )  ;
assign n13804 =  ( n19 ) & ( n13688 )  ;
assign n13805 =  ( n19 ) & ( n13690 )  ;
assign n13806 =  ( n19 ) & ( n13692 )  ;
assign n13807 =  ( n19 ) & ( n13694 )  ;
assign n13808 =  ( n20 ) & ( n13664 )  ;
assign n13809 =  ( n20 ) & ( n13666 )  ;
assign n13810 =  ( n20 ) & ( n13668 )  ;
assign n13811 =  ( n20 ) & ( n13670 )  ;
assign n13812 =  ( n20 ) & ( n13672 )  ;
assign n13813 =  ( n20 ) & ( n13674 )  ;
assign n13814 =  ( n20 ) & ( n13676 )  ;
assign n13815 =  ( n20 ) & ( n13678 )  ;
assign n13816 =  ( n20 ) & ( n13680 )  ;
assign n13817 =  ( n20 ) & ( n13682 )  ;
assign n13818 =  ( n20 ) & ( n13684 )  ;
assign n13819 =  ( n20 ) & ( n13686 )  ;
assign n13820 =  ( n20 ) & ( n13688 )  ;
assign n13821 =  ( n20 ) & ( n13690 )  ;
assign n13822 =  ( n20 ) & ( n13692 )  ;
assign n13823 =  ( n20 ) & ( n13694 )  ;
assign n13824 =  ( n21 ) & ( n13664 )  ;
assign n13825 =  ( n21 ) & ( n13666 )  ;
assign n13826 =  ( n21 ) & ( n13668 )  ;
assign n13827 =  ( n21 ) & ( n13670 )  ;
assign n13828 =  ( n21 ) & ( n13672 )  ;
assign n13829 =  ( n21 ) & ( n13674 )  ;
assign n13830 =  ( n21 ) & ( n13676 )  ;
assign n13831 =  ( n21 ) & ( n13678 )  ;
assign n13832 =  ( n21 ) & ( n13680 )  ;
assign n13833 =  ( n21 ) & ( n13682 )  ;
assign n13834 =  ( n21 ) & ( n13684 )  ;
assign n13835 =  ( n21 ) & ( n13686 )  ;
assign n13836 =  ( n21 ) & ( n13688 )  ;
assign n13837 =  ( n21 ) & ( n13690 )  ;
assign n13838 =  ( n21 ) & ( n13692 )  ;
assign n13839 =  ( n21 ) & ( n13694 )  ;
assign n13840 =  ( n22 ) & ( n13664 )  ;
assign n13841 =  ( n22 ) & ( n13666 )  ;
assign n13842 =  ( n22 ) & ( n13668 )  ;
assign n13843 =  ( n22 ) & ( n13670 )  ;
assign n13844 =  ( n22 ) & ( n13672 )  ;
assign n13845 =  ( n22 ) & ( n13674 )  ;
assign n13846 =  ( n22 ) & ( n13676 )  ;
assign n13847 =  ( n22 ) & ( n13678 )  ;
assign n13848 =  ( n22 ) & ( n13680 )  ;
assign n13849 =  ( n22 ) & ( n13682 )  ;
assign n13850 =  ( n22 ) & ( n13684 )  ;
assign n13851 =  ( n22 ) & ( n13686 )  ;
assign n13852 =  ( n22 ) & ( n13688 )  ;
assign n13853 =  ( n22 ) & ( n13690 )  ;
assign n13854 =  ( n22 ) & ( n13692 )  ;
assign n13855 =  ( n22 ) & ( n13694 )  ;
assign n13856 =  ( n23 ) & ( n13664 )  ;
assign n13857 =  ( n23 ) & ( n13666 )  ;
assign n13858 =  ( n23 ) & ( n13668 )  ;
assign n13859 =  ( n23 ) & ( n13670 )  ;
assign n13860 =  ( n23 ) & ( n13672 )  ;
assign n13861 =  ( n23 ) & ( n13674 )  ;
assign n13862 =  ( n23 ) & ( n13676 )  ;
assign n13863 =  ( n23 ) & ( n13678 )  ;
assign n13864 =  ( n23 ) & ( n13680 )  ;
assign n13865 =  ( n23 ) & ( n13682 )  ;
assign n13866 =  ( n23 ) & ( n13684 )  ;
assign n13867 =  ( n23 ) & ( n13686 )  ;
assign n13868 =  ( n23 ) & ( n13688 )  ;
assign n13869 =  ( n23 ) & ( n13690 )  ;
assign n13870 =  ( n23 ) & ( n13692 )  ;
assign n13871 =  ( n23 ) & ( n13694 )  ;
assign n13872 =  ( n24 ) & ( n13664 )  ;
assign n13873 =  ( n24 ) & ( n13666 )  ;
assign n13874 =  ( n24 ) & ( n13668 )  ;
assign n13875 =  ( n24 ) & ( n13670 )  ;
assign n13876 =  ( n24 ) & ( n13672 )  ;
assign n13877 =  ( n24 ) & ( n13674 )  ;
assign n13878 =  ( n24 ) & ( n13676 )  ;
assign n13879 =  ( n24 ) & ( n13678 )  ;
assign n13880 =  ( n24 ) & ( n13680 )  ;
assign n13881 =  ( n24 ) & ( n13682 )  ;
assign n13882 =  ( n24 ) & ( n13684 )  ;
assign n13883 =  ( n24 ) & ( n13686 )  ;
assign n13884 =  ( n24 ) & ( n13688 )  ;
assign n13885 =  ( n24 ) & ( n13690 )  ;
assign n13886 =  ( n24 ) & ( n13692 )  ;
assign n13887 =  ( n24 ) & ( n13694 )  ;
assign n13888 =  ( n25 ) & ( n13664 )  ;
assign n13889 =  ( n25 ) & ( n13666 )  ;
assign n13890 =  ( n25 ) & ( n13668 )  ;
assign n13891 =  ( n25 ) & ( n13670 )  ;
assign n13892 =  ( n25 ) & ( n13672 )  ;
assign n13893 =  ( n25 ) & ( n13674 )  ;
assign n13894 =  ( n25 ) & ( n13676 )  ;
assign n13895 =  ( n25 ) & ( n13678 )  ;
assign n13896 =  ( n25 ) & ( n13680 )  ;
assign n13897 =  ( n25 ) & ( n13682 )  ;
assign n13898 =  ( n25 ) & ( n13684 )  ;
assign n13899 =  ( n25 ) & ( n13686 )  ;
assign n13900 =  ( n25 ) & ( n13688 )  ;
assign n13901 =  ( n25 ) & ( n13690 )  ;
assign n13902 =  ( n25 ) & ( n13692 )  ;
assign n13903 =  ( n25 ) & ( n13694 )  ;
assign n13904 =  ( n26 ) & ( n13664 )  ;
assign n13905 =  ( n26 ) & ( n13666 )  ;
assign n13906 =  ( n26 ) & ( n13668 )  ;
assign n13907 =  ( n26 ) & ( n13670 )  ;
assign n13908 =  ( n26 ) & ( n13672 )  ;
assign n13909 =  ( n26 ) & ( n13674 )  ;
assign n13910 =  ( n26 ) & ( n13676 )  ;
assign n13911 =  ( n26 ) & ( n13678 )  ;
assign n13912 =  ( n26 ) & ( n13680 )  ;
assign n13913 =  ( n26 ) & ( n13682 )  ;
assign n13914 =  ( n26 ) & ( n13684 )  ;
assign n13915 =  ( n26 ) & ( n13686 )  ;
assign n13916 =  ( n26 ) & ( n13688 )  ;
assign n13917 =  ( n26 ) & ( n13690 )  ;
assign n13918 =  ( n26 ) & ( n13692 )  ;
assign n13919 =  ( n26 ) & ( n13694 )  ;
assign n13920 =  ( n27 ) & ( n13664 )  ;
assign n13921 =  ( n27 ) & ( n13666 )  ;
assign n13922 =  ( n27 ) & ( n13668 )  ;
assign n13923 =  ( n27 ) & ( n13670 )  ;
assign n13924 =  ( n27 ) & ( n13672 )  ;
assign n13925 =  ( n27 ) & ( n13674 )  ;
assign n13926 =  ( n27 ) & ( n13676 )  ;
assign n13927 =  ( n27 ) & ( n13678 )  ;
assign n13928 =  ( n27 ) & ( n13680 )  ;
assign n13929 =  ( n27 ) & ( n13682 )  ;
assign n13930 =  ( n27 ) & ( n13684 )  ;
assign n13931 =  ( n27 ) & ( n13686 )  ;
assign n13932 =  ( n27 ) & ( n13688 )  ;
assign n13933 =  ( n27 ) & ( n13690 )  ;
assign n13934 =  ( n27 ) & ( n13692 )  ;
assign n13935 =  ( n27 ) & ( n13694 )  ;
assign n13936 =  ( n28 ) & ( n13664 )  ;
assign n13937 =  ( n28 ) & ( n13666 )  ;
assign n13938 =  ( n28 ) & ( n13668 )  ;
assign n13939 =  ( n28 ) & ( n13670 )  ;
assign n13940 =  ( n28 ) & ( n13672 )  ;
assign n13941 =  ( n28 ) & ( n13674 )  ;
assign n13942 =  ( n28 ) & ( n13676 )  ;
assign n13943 =  ( n28 ) & ( n13678 )  ;
assign n13944 =  ( n28 ) & ( n13680 )  ;
assign n13945 =  ( n28 ) & ( n13682 )  ;
assign n13946 =  ( n28 ) & ( n13684 )  ;
assign n13947 =  ( n28 ) & ( n13686 )  ;
assign n13948 =  ( n28 ) & ( n13688 )  ;
assign n13949 =  ( n28 ) & ( n13690 )  ;
assign n13950 =  ( n28 ) & ( n13692 )  ;
assign n13951 =  ( n28 ) & ( n13694 )  ;
assign n13952 =  ( n29 ) & ( n13664 )  ;
assign n13953 =  ( n29 ) & ( n13666 )  ;
assign n13954 =  ( n29 ) & ( n13668 )  ;
assign n13955 =  ( n29 ) & ( n13670 )  ;
assign n13956 =  ( n29 ) & ( n13672 )  ;
assign n13957 =  ( n29 ) & ( n13674 )  ;
assign n13958 =  ( n29 ) & ( n13676 )  ;
assign n13959 =  ( n29 ) & ( n13678 )  ;
assign n13960 =  ( n29 ) & ( n13680 )  ;
assign n13961 =  ( n29 ) & ( n13682 )  ;
assign n13962 =  ( n29 ) & ( n13684 )  ;
assign n13963 =  ( n29 ) & ( n13686 )  ;
assign n13964 =  ( n29 ) & ( n13688 )  ;
assign n13965 =  ( n29 ) & ( n13690 )  ;
assign n13966 =  ( n29 ) & ( n13692 )  ;
assign n13967 =  ( n29 ) & ( n13694 )  ;
assign n13968 =  ( n30 ) & ( n13664 )  ;
assign n13969 =  ( n30 ) & ( n13666 )  ;
assign n13970 =  ( n30 ) & ( n13668 )  ;
assign n13971 =  ( n30 ) & ( n13670 )  ;
assign n13972 =  ( n30 ) & ( n13672 )  ;
assign n13973 =  ( n30 ) & ( n13674 )  ;
assign n13974 =  ( n30 ) & ( n13676 )  ;
assign n13975 =  ( n30 ) & ( n13678 )  ;
assign n13976 =  ( n30 ) & ( n13680 )  ;
assign n13977 =  ( n30 ) & ( n13682 )  ;
assign n13978 =  ( n30 ) & ( n13684 )  ;
assign n13979 =  ( n30 ) & ( n13686 )  ;
assign n13980 =  ( n30 ) & ( n13688 )  ;
assign n13981 =  ( n30 ) & ( n13690 )  ;
assign n13982 =  ( n30 ) & ( n13692 )  ;
assign n13983 =  ( n30 ) & ( n13694 )  ;
assign n13984 =  ( n31 ) & ( n13664 )  ;
assign n13985 =  ( n31 ) & ( n13666 )  ;
assign n13986 =  ( n31 ) & ( n13668 )  ;
assign n13987 =  ( n31 ) & ( n13670 )  ;
assign n13988 =  ( n31 ) & ( n13672 )  ;
assign n13989 =  ( n31 ) & ( n13674 )  ;
assign n13990 =  ( n31 ) & ( n13676 )  ;
assign n13991 =  ( n31 ) & ( n13678 )  ;
assign n13992 =  ( n31 ) & ( n13680 )  ;
assign n13993 =  ( n31 ) & ( n13682 )  ;
assign n13994 =  ( n31 ) & ( n13684 )  ;
assign n13995 =  ( n31 ) & ( n13686 )  ;
assign n13996 =  ( n31 ) & ( n13688 )  ;
assign n13997 =  ( n31 ) & ( n13690 )  ;
assign n13998 =  ( n31 ) & ( n13692 )  ;
assign n13999 =  ( n31 ) & ( n13694 )  ;
assign n14000 =  ( n32 ) & ( n13664 )  ;
assign n14001 =  ( n32 ) & ( n13666 )  ;
assign n14002 =  ( n32 ) & ( n13668 )  ;
assign n14003 =  ( n32 ) & ( n13670 )  ;
assign n14004 =  ( n32 ) & ( n13672 )  ;
assign n14005 =  ( n32 ) & ( n13674 )  ;
assign n14006 =  ( n32 ) & ( n13676 )  ;
assign n14007 =  ( n32 ) & ( n13678 )  ;
assign n14008 =  ( n32 ) & ( n13680 )  ;
assign n14009 =  ( n32 ) & ( n13682 )  ;
assign n14010 =  ( n32 ) & ( n13684 )  ;
assign n14011 =  ( n32 ) & ( n13686 )  ;
assign n14012 =  ( n32 ) & ( n13688 )  ;
assign n14013 =  ( n32 ) & ( n13690 )  ;
assign n14014 =  ( n32 ) & ( n13692 )  ;
assign n14015 =  ( n32 ) & ( n13694 )  ;
assign n14016 =  ( n33 ) & ( n13664 )  ;
assign n14017 =  ( n33 ) & ( n13666 )  ;
assign n14018 =  ( n33 ) & ( n13668 )  ;
assign n14019 =  ( n33 ) & ( n13670 )  ;
assign n14020 =  ( n33 ) & ( n13672 )  ;
assign n14021 =  ( n33 ) & ( n13674 )  ;
assign n14022 =  ( n33 ) & ( n13676 )  ;
assign n14023 =  ( n33 ) & ( n13678 )  ;
assign n14024 =  ( n33 ) & ( n13680 )  ;
assign n14025 =  ( n33 ) & ( n13682 )  ;
assign n14026 =  ( n33 ) & ( n13684 )  ;
assign n14027 =  ( n33 ) & ( n13686 )  ;
assign n14028 =  ( n33 ) & ( n13688 )  ;
assign n14029 =  ( n33 ) & ( n13690 )  ;
assign n14030 =  ( n33 ) & ( n13692 )  ;
assign n14031 =  ( n33 ) & ( n13694 )  ;
assign n14032 =  ( n34 ) & ( n13664 )  ;
assign n14033 =  ( n34 ) & ( n13666 )  ;
assign n14034 =  ( n34 ) & ( n13668 )  ;
assign n14035 =  ( n34 ) & ( n13670 )  ;
assign n14036 =  ( n34 ) & ( n13672 )  ;
assign n14037 =  ( n34 ) & ( n13674 )  ;
assign n14038 =  ( n34 ) & ( n13676 )  ;
assign n14039 =  ( n34 ) & ( n13678 )  ;
assign n14040 =  ( n34 ) & ( n13680 )  ;
assign n14041 =  ( n34 ) & ( n13682 )  ;
assign n14042 =  ( n34 ) & ( n13684 )  ;
assign n14043 =  ( n34 ) & ( n13686 )  ;
assign n14044 =  ( n34 ) & ( n13688 )  ;
assign n14045 =  ( n34 ) & ( n13690 )  ;
assign n14046 =  ( n34 ) & ( n13692 )  ;
assign n14047 =  ( n34 ) & ( n13694 )  ;
assign n14048 =  ( n35 ) & ( n13664 )  ;
assign n14049 =  ( n35 ) & ( n13666 )  ;
assign n14050 =  ( n35 ) & ( n13668 )  ;
assign n14051 =  ( n35 ) & ( n13670 )  ;
assign n14052 =  ( n35 ) & ( n13672 )  ;
assign n14053 =  ( n35 ) & ( n13674 )  ;
assign n14054 =  ( n35 ) & ( n13676 )  ;
assign n14055 =  ( n35 ) & ( n13678 )  ;
assign n14056 =  ( n35 ) & ( n13680 )  ;
assign n14057 =  ( n35 ) & ( n13682 )  ;
assign n14058 =  ( n35 ) & ( n13684 )  ;
assign n14059 =  ( n35 ) & ( n13686 )  ;
assign n14060 =  ( n35 ) & ( n13688 )  ;
assign n14061 =  ( n35 ) & ( n13690 )  ;
assign n14062 =  ( n35 ) & ( n13692 )  ;
assign n14063 =  ( n35 ) & ( n13694 )  ;
assign n14064 =  ( n36 ) & ( n13664 )  ;
assign n14065 =  ( n36 ) & ( n13666 )  ;
assign n14066 =  ( n36 ) & ( n13668 )  ;
assign n14067 =  ( n36 ) & ( n13670 )  ;
assign n14068 =  ( n36 ) & ( n13672 )  ;
assign n14069 =  ( n36 ) & ( n13674 )  ;
assign n14070 =  ( n36 ) & ( n13676 )  ;
assign n14071 =  ( n36 ) & ( n13678 )  ;
assign n14072 =  ( n36 ) & ( n13680 )  ;
assign n14073 =  ( n36 ) & ( n13682 )  ;
assign n14074 =  ( n36 ) & ( n13684 )  ;
assign n14075 =  ( n36 ) & ( n13686 )  ;
assign n14076 =  ( n36 ) & ( n13688 )  ;
assign n14077 =  ( n36 ) & ( n13690 )  ;
assign n14078 =  ( n36 ) & ( n13692 )  ;
assign n14079 =  ( n36 ) & ( n13694 )  ;
assign n14080 =  ( n37 ) & ( n13664 )  ;
assign n14081 =  ( n37 ) & ( n13666 )  ;
assign n14082 =  ( n37 ) & ( n13668 )  ;
assign n14083 =  ( n37 ) & ( n13670 )  ;
assign n14084 =  ( n37 ) & ( n13672 )  ;
assign n14085 =  ( n37 ) & ( n13674 )  ;
assign n14086 =  ( n37 ) & ( n13676 )  ;
assign n14087 =  ( n37 ) & ( n13678 )  ;
assign n14088 =  ( n37 ) & ( n13680 )  ;
assign n14089 =  ( n37 ) & ( n13682 )  ;
assign n14090 =  ( n37 ) & ( n13684 )  ;
assign n14091 =  ( n37 ) & ( n13686 )  ;
assign n14092 =  ( n37 ) & ( n13688 )  ;
assign n14093 =  ( n37 ) & ( n13690 )  ;
assign n14094 =  ( n37 ) & ( n13692 )  ;
assign n14095 =  ( n37 ) & ( n13694 )  ;
assign n14096 =  ( n38 ) & ( n13664 )  ;
assign n14097 =  ( n38 ) & ( n13666 )  ;
assign n14098 =  ( n38 ) & ( n13668 )  ;
assign n14099 =  ( n38 ) & ( n13670 )  ;
assign n14100 =  ( n38 ) & ( n13672 )  ;
assign n14101 =  ( n38 ) & ( n13674 )  ;
assign n14102 =  ( n38 ) & ( n13676 )  ;
assign n14103 =  ( n38 ) & ( n13678 )  ;
assign n14104 =  ( n38 ) & ( n13680 )  ;
assign n14105 =  ( n38 ) & ( n13682 )  ;
assign n14106 =  ( n38 ) & ( n13684 )  ;
assign n14107 =  ( n38 ) & ( n13686 )  ;
assign n14108 =  ( n38 ) & ( n13688 )  ;
assign n14109 =  ( n38 ) & ( n13690 )  ;
assign n14110 =  ( n38 ) & ( n13692 )  ;
assign n14111 =  ( n38 ) & ( n13694 )  ;
assign n14112 =  ( n39 ) & ( n13664 )  ;
assign n14113 =  ( n39 ) & ( n13666 )  ;
assign n14114 =  ( n39 ) & ( n13668 )  ;
assign n14115 =  ( n39 ) & ( n13670 )  ;
assign n14116 =  ( n39 ) & ( n13672 )  ;
assign n14117 =  ( n39 ) & ( n13674 )  ;
assign n14118 =  ( n39 ) & ( n13676 )  ;
assign n14119 =  ( n39 ) & ( n13678 )  ;
assign n14120 =  ( n39 ) & ( n13680 )  ;
assign n14121 =  ( n39 ) & ( n13682 )  ;
assign n14122 =  ( n39 ) & ( n13684 )  ;
assign n14123 =  ( n39 ) & ( n13686 )  ;
assign n14124 =  ( n39 ) & ( n13688 )  ;
assign n14125 =  ( n39 ) & ( n13690 )  ;
assign n14126 =  ( n39 ) & ( n13692 )  ;
assign n14127 =  ( n39 ) & ( n13694 )  ;
assign n14128 =  ( n40 ) & ( n13664 )  ;
assign n14129 =  ( n40 ) & ( n13666 )  ;
assign n14130 =  ( n40 ) & ( n13668 )  ;
assign n14131 =  ( n40 ) & ( n13670 )  ;
assign n14132 =  ( n40 ) & ( n13672 )  ;
assign n14133 =  ( n40 ) & ( n13674 )  ;
assign n14134 =  ( n40 ) & ( n13676 )  ;
assign n14135 =  ( n40 ) & ( n13678 )  ;
assign n14136 =  ( n40 ) & ( n13680 )  ;
assign n14137 =  ( n40 ) & ( n13682 )  ;
assign n14138 =  ( n40 ) & ( n13684 )  ;
assign n14139 =  ( n40 ) & ( n13686 )  ;
assign n14140 =  ( n40 ) & ( n13688 )  ;
assign n14141 =  ( n40 ) & ( n13690 )  ;
assign n14142 =  ( n40 ) & ( n13692 )  ;
assign n14143 =  ( n40 ) & ( n13694 )  ;
assign n14144 =  ( n41 ) & ( n13664 )  ;
assign n14145 =  ( n41 ) & ( n13666 )  ;
assign n14146 =  ( n41 ) & ( n13668 )  ;
assign n14147 =  ( n41 ) & ( n13670 )  ;
assign n14148 =  ( n41 ) & ( n13672 )  ;
assign n14149 =  ( n41 ) & ( n13674 )  ;
assign n14150 =  ( n41 ) & ( n13676 )  ;
assign n14151 =  ( n41 ) & ( n13678 )  ;
assign n14152 =  ( n41 ) & ( n13680 )  ;
assign n14153 =  ( n41 ) & ( n13682 )  ;
assign n14154 =  ( n41 ) & ( n13684 )  ;
assign n14155 =  ( n41 ) & ( n13686 )  ;
assign n14156 =  ( n41 ) & ( n13688 )  ;
assign n14157 =  ( n41 ) & ( n13690 )  ;
assign n14158 =  ( n41 ) & ( n13692 )  ;
assign n14159 =  ( n41 ) & ( n13694 )  ;
assign n14160 =  ( n42 ) & ( n13664 )  ;
assign n14161 =  ( n42 ) & ( n13666 )  ;
assign n14162 =  ( n42 ) & ( n13668 )  ;
assign n14163 =  ( n42 ) & ( n13670 )  ;
assign n14164 =  ( n42 ) & ( n13672 )  ;
assign n14165 =  ( n42 ) & ( n13674 )  ;
assign n14166 =  ( n42 ) & ( n13676 )  ;
assign n14167 =  ( n42 ) & ( n13678 )  ;
assign n14168 =  ( n42 ) & ( n13680 )  ;
assign n14169 =  ( n42 ) & ( n13682 )  ;
assign n14170 =  ( n42 ) & ( n13684 )  ;
assign n14171 =  ( n42 ) & ( n13686 )  ;
assign n14172 =  ( n42 ) & ( n13688 )  ;
assign n14173 =  ( n42 ) & ( n13690 )  ;
assign n14174 =  ( n42 ) & ( n13692 )  ;
assign n14175 =  ( n42 ) & ( n13694 )  ;
assign n14176 =  ( n43 ) & ( n13664 )  ;
assign n14177 =  ( n43 ) & ( n13666 )  ;
assign n14178 =  ( n43 ) & ( n13668 )  ;
assign n14179 =  ( n43 ) & ( n13670 )  ;
assign n14180 =  ( n43 ) & ( n13672 )  ;
assign n14181 =  ( n43 ) & ( n13674 )  ;
assign n14182 =  ( n43 ) & ( n13676 )  ;
assign n14183 =  ( n43 ) & ( n13678 )  ;
assign n14184 =  ( n43 ) & ( n13680 )  ;
assign n14185 =  ( n43 ) & ( n13682 )  ;
assign n14186 =  ( n43 ) & ( n13684 )  ;
assign n14187 =  ( n43 ) & ( n13686 )  ;
assign n14188 =  ( n43 ) & ( n13688 )  ;
assign n14189 =  ( n43 ) & ( n13690 )  ;
assign n14190 =  ( n43 ) & ( n13692 )  ;
assign n14191 =  ( n43 ) & ( n13694 )  ;
assign n14192 =  ( n14191 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n14193 =  ( n14190 ) ? ( VREG_0_1 ) : ( n14192 ) ;
assign n14194 =  ( n14189 ) ? ( VREG_0_2 ) : ( n14193 ) ;
assign n14195 =  ( n14188 ) ? ( VREG_0_3 ) : ( n14194 ) ;
assign n14196 =  ( n14187 ) ? ( VREG_0_4 ) : ( n14195 ) ;
assign n14197 =  ( n14186 ) ? ( VREG_0_5 ) : ( n14196 ) ;
assign n14198 =  ( n14185 ) ? ( VREG_0_6 ) : ( n14197 ) ;
assign n14199 =  ( n14184 ) ? ( VREG_0_7 ) : ( n14198 ) ;
assign n14200 =  ( n14183 ) ? ( VREG_0_8 ) : ( n14199 ) ;
assign n14201 =  ( n14182 ) ? ( VREG_0_9 ) : ( n14200 ) ;
assign n14202 =  ( n14181 ) ? ( VREG_0_10 ) : ( n14201 ) ;
assign n14203 =  ( n14180 ) ? ( VREG_0_11 ) : ( n14202 ) ;
assign n14204 =  ( n14179 ) ? ( VREG_0_12 ) : ( n14203 ) ;
assign n14205 =  ( n14178 ) ? ( VREG_0_13 ) : ( n14204 ) ;
assign n14206 =  ( n14177 ) ? ( VREG_0_14 ) : ( n14205 ) ;
assign n14207 =  ( n14176 ) ? ( VREG_0_15 ) : ( n14206 ) ;
assign n14208 =  ( n14175 ) ? ( VREG_1_0 ) : ( n14207 ) ;
assign n14209 =  ( n14174 ) ? ( VREG_1_1 ) : ( n14208 ) ;
assign n14210 =  ( n14173 ) ? ( VREG_1_2 ) : ( n14209 ) ;
assign n14211 =  ( n14172 ) ? ( VREG_1_3 ) : ( n14210 ) ;
assign n14212 =  ( n14171 ) ? ( VREG_1_4 ) : ( n14211 ) ;
assign n14213 =  ( n14170 ) ? ( VREG_1_5 ) : ( n14212 ) ;
assign n14214 =  ( n14169 ) ? ( VREG_1_6 ) : ( n14213 ) ;
assign n14215 =  ( n14168 ) ? ( VREG_1_7 ) : ( n14214 ) ;
assign n14216 =  ( n14167 ) ? ( VREG_1_8 ) : ( n14215 ) ;
assign n14217 =  ( n14166 ) ? ( VREG_1_9 ) : ( n14216 ) ;
assign n14218 =  ( n14165 ) ? ( VREG_1_10 ) : ( n14217 ) ;
assign n14219 =  ( n14164 ) ? ( VREG_1_11 ) : ( n14218 ) ;
assign n14220 =  ( n14163 ) ? ( VREG_1_12 ) : ( n14219 ) ;
assign n14221 =  ( n14162 ) ? ( VREG_1_13 ) : ( n14220 ) ;
assign n14222 =  ( n14161 ) ? ( VREG_1_14 ) : ( n14221 ) ;
assign n14223 =  ( n14160 ) ? ( VREG_1_15 ) : ( n14222 ) ;
assign n14224 =  ( n14159 ) ? ( VREG_2_0 ) : ( n14223 ) ;
assign n14225 =  ( n14158 ) ? ( VREG_2_1 ) : ( n14224 ) ;
assign n14226 =  ( n14157 ) ? ( VREG_2_2 ) : ( n14225 ) ;
assign n14227 =  ( n14156 ) ? ( VREG_2_3 ) : ( n14226 ) ;
assign n14228 =  ( n14155 ) ? ( VREG_2_4 ) : ( n14227 ) ;
assign n14229 =  ( n14154 ) ? ( VREG_2_5 ) : ( n14228 ) ;
assign n14230 =  ( n14153 ) ? ( VREG_2_6 ) : ( n14229 ) ;
assign n14231 =  ( n14152 ) ? ( VREG_2_7 ) : ( n14230 ) ;
assign n14232 =  ( n14151 ) ? ( VREG_2_8 ) : ( n14231 ) ;
assign n14233 =  ( n14150 ) ? ( VREG_2_9 ) : ( n14232 ) ;
assign n14234 =  ( n14149 ) ? ( VREG_2_10 ) : ( n14233 ) ;
assign n14235 =  ( n14148 ) ? ( VREG_2_11 ) : ( n14234 ) ;
assign n14236 =  ( n14147 ) ? ( VREG_2_12 ) : ( n14235 ) ;
assign n14237 =  ( n14146 ) ? ( VREG_2_13 ) : ( n14236 ) ;
assign n14238 =  ( n14145 ) ? ( VREG_2_14 ) : ( n14237 ) ;
assign n14239 =  ( n14144 ) ? ( VREG_2_15 ) : ( n14238 ) ;
assign n14240 =  ( n14143 ) ? ( VREG_3_0 ) : ( n14239 ) ;
assign n14241 =  ( n14142 ) ? ( VREG_3_1 ) : ( n14240 ) ;
assign n14242 =  ( n14141 ) ? ( VREG_3_2 ) : ( n14241 ) ;
assign n14243 =  ( n14140 ) ? ( VREG_3_3 ) : ( n14242 ) ;
assign n14244 =  ( n14139 ) ? ( VREG_3_4 ) : ( n14243 ) ;
assign n14245 =  ( n14138 ) ? ( VREG_3_5 ) : ( n14244 ) ;
assign n14246 =  ( n14137 ) ? ( VREG_3_6 ) : ( n14245 ) ;
assign n14247 =  ( n14136 ) ? ( VREG_3_7 ) : ( n14246 ) ;
assign n14248 =  ( n14135 ) ? ( VREG_3_8 ) : ( n14247 ) ;
assign n14249 =  ( n14134 ) ? ( VREG_3_9 ) : ( n14248 ) ;
assign n14250 =  ( n14133 ) ? ( VREG_3_10 ) : ( n14249 ) ;
assign n14251 =  ( n14132 ) ? ( VREG_3_11 ) : ( n14250 ) ;
assign n14252 =  ( n14131 ) ? ( VREG_3_12 ) : ( n14251 ) ;
assign n14253 =  ( n14130 ) ? ( VREG_3_13 ) : ( n14252 ) ;
assign n14254 =  ( n14129 ) ? ( VREG_3_14 ) : ( n14253 ) ;
assign n14255 =  ( n14128 ) ? ( VREG_3_15 ) : ( n14254 ) ;
assign n14256 =  ( n14127 ) ? ( VREG_4_0 ) : ( n14255 ) ;
assign n14257 =  ( n14126 ) ? ( VREG_4_1 ) : ( n14256 ) ;
assign n14258 =  ( n14125 ) ? ( VREG_4_2 ) : ( n14257 ) ;
assign n14259 =  ( n14124 ) ? ( VREG_4_3 ) : ( n14258 ) ;
assign n14260 =  ( n14123 ) ? ( VREG_4_4 ) : ( n14259 ) ;
assign n14261 =  ( n14122 ) ? ( VREG_4_5 ) : ( n14260 ) ;
assign n14262 =  ( n14121 ) ? ( VREG_4_6 ) : ( n14261 ) ;
assign n14263 =  ( n14120 ) ? ( VREG_4_7 ) : ( n14262 ) ;
assign n14264 =  ( n14119 ) ? ( VREG_4_8 ) : ( n14263 ) ;
assign n14265 =  ( n14118 ) ? ( VREG_4_9 ) : ( n14264 ) ;
assign n14266 =  ( n14117 ) ? ( VREG_4_10 ) : ( n14265 ) ;
assign n14267 =  ( n14116 ) ? ( VREG_4_11 ) : ( n14266 ) ;
assign n14268 =  ( n14115 ) ? ( VREG_4_12 ) : ( n14267 ) ;
assign n14269 =  ( n14114 ) ? ( VREG_4_13 ) : ( n14268 ) ;
assign n14270 =  ( n14113 ) ? ( VREG_4_14 ) : ( n14269 ) ;
assign n14271 =  ( n14112 ) ? ( VREG_4_15 ) : ( n14270 ) ;
assign n14272 =  ( n14111 ) ? ( VREG_5_0 ) : ( n14271 ) ;
assign n14273 =  ( n14110 ) ? ( VREG_5_1 ) : ( n14272 ) ;
assign n14274 =  ( n14109 ) ? ( VREG_5_2 ) : ( n14273 ) ;
assign n14275 =  ( n14108 ) ? ( VREG_5_3 ) : ( n14274 ) ;
assign n14276 =  ( n14107 ) ? ( VREG_5_4 ) : ( n14275 ) ;
assign n14277 =  ( n14106 ) ? ( VREG_5_5 ) : ( n14276 ) ;
assign n14278 =  ( n14105 ) ? ( VREG_5_6 ) : ( n14277 ) ;
assign n14279 =  ( n14104 ) ? ( VREG_5_7 ) : ( n14278 ) ;
assign n14280 =  ( n14103 ) ? ( VREG_5_8 ) : ( n14279 ) ;
assign n14281 =  ( n14102 ) ? ( VREG_5_9 ) : ( n14280 ) ;
assign n14282 =  ( n14101 ) ? ( VREG_5_10 ) : ( n14281 ) ;
assign n14283 =  ( n14100 ) ? ( VREG_5_11 ) : ( n14282 ) ;
assign n14284 =  ( n14099 ) ? ( VREG_5_12 ) : ( n14283 ) ;
assign n14285 =  ( n14098 ) ? ( VREG_5_13 ) : ( n14284 ) ;
assign n14286 =  ( n14097 ) ? ( VREG_5_14 ) : ( n14285 ) ;
assign n14287 =  ( n14096 ) ? ( VREG_5_15 ) : ( n14286 ) ;
assign n14288 =  ( n14095 ) ? ( VREG_6_0 ) : ( n14287 ) ;
assign n14289 =  ( n14094 ) ? ( VREG_6_1 ) : ( n14288 ) ;
assign n14290 =  ( n14093 ) ? ( VREG_6_2 ) : ( n14289 ) ;
assign n14291 =  ( n14092 ) ? ( VREG_6_3 ) : ( n14290 ) ;
assign n14292 =  ( n14091 ) ? ( VREG_6_4 ) : ( n14291 ) ;
assign n14293 =  ( n14090 ) ? ( VREG_6_5 ) : ( n14292 ) ;
assign n14294 =  ( n14089 ) ? ( VREG_6_6 ) : ( n14293 ) ;
assign n14295 =  ( n14088 ) ? ( VREG_6_7 ) : ( n14294 ) ;
assign n14296 =  ( n14087 ) ? ( VREG_6_8 ) : ( n14295 ) ;
assign n14297 =  ( n14086 ) ? ( VREG_6_9 ) : ( n14296 ) ;
assign n14298 =  ( n14085 ) ? ( VREG_6_10 ) : ( n14297 ) ;
assign n14299 =  ( n14084 ) ? ( VREG_6_11 ) : ( n14298 ) ;
assign n14300 =  ( n14083 ) ? ( VREG_6_12 ) : ( n14299 ) ;
assign n14301 =  ( n14082 ) ? ( VREG_6_13 ) : ( n14300 ) ;
assign n14302 =  ( n14081 ) ? ( VREG_6_14 ) : ( n14301 ) ;
assign n14303 =  ( n14080 ) ? ( VREG_6_15 ) : ( n14302 ) ;
assign n14304 =  ( n14079 ) ? ( VREG_7_0 ) : ( n14303 ) ;
assign n14305 =  ( n14078 ) ? ( VREG_7_1 ) : ( n14304 ) ;
assign n14306 =  ( n14077 ) ? ( VREG_7_2 ) : ( n14305 ) ;
assign n14307 =  ( n14076 ) ? ( VREG_7_3 ) : ( n14306 ) ;
assign n14308 =  ( n14075 ) ? ( VREG_7_4 ) : ( n14307 ) ;
assign n14309 =  ( n14074 ) ? ( VREG_7_5 ) : ( n14308 ) ;
assign n14310 =  ( n14073 ) ? ( VREG_7_6 ) : ( n14309 ) ;
assign n14311 =  ( n14072 ) ? ( VREG_7_7 ) : ( n14310 ) ;
assign n14312 =  ( n14071 ) ? ( VREG_7_8 ) : ( n14311 ) ;
assign n14313 =  ( n14070 ) ? ( VREG_7_9 ) : ( n14312 ) ;
assign n14314 =  ( n14069 ) ? ( VREG_7_10 ) : ( n14313 ) ;
assign n14315 =  ( n14068 ) ? ( VREG_7_11 ) : ( n14314 ) ;
assign n14316 =  ( n14067 ) ? ( VREG_7_12 ) : ( n14315 ) ;
assign n14317 =  ( n14066 ) ? ( VREG_7_13 ) : ( n14316 ) ;
assign n14318 =  ( n14065 ) ? ( VREG_7_14 ) : ( n14317 ) ;
assign n14319 =  ( n14064 ) ? ( VREG_7_15 ) : ( n14318 ) ;
assign n14320 =  ( n14063 ) ? ( VREG_8_0 ) : ( n14319 ) ;
assign n14321 =  ( n14062 ) ? ( VREG_8_1 ) : ( n14320 ) ;
assign n14322 =  ( n14061 ) ? ( VREG_8_2 ) : ( n14321 ) ;
assign n14323 =  ( n14060 ) ? ( VREG_8_3 ) : ( n14322 ) ;
assign n14324 =  ( n14059 ) ? ( VREG_8_4 ) : ( n14323 ) ;
assign n14325 =  ( n14058 ) ? ( VREG_8_5 ) : ( n14324 ) ;
assign n14326 =  ( n14057 ) ? ( VREG_8_6 ) : ( n14325 ) ;
assign n14327 =  ( n14056 ) ? ( VREG_8_7 ) : ( n14326 ) ;
assign n14328 =  ( n14055 ) ? ( VREG_8_8 ) : ( n14327 ) ;
assign n14329 =  ( n14054 ) ? ( VREG_8_9 ) : ( n14328 ) ;
assign n14330 =  ( n14053 ) ? ( VREG_8_10 ) : ( n14329 ) ;
assign n14331 =  ( n14052 ) ? ( VREG_8_11 ) : ( n14330 ) ;
assign n14332 =  ( n14051 ) ? ( VREG_8_12 ) : ( n14331 ) ;
assign n14333 =  ( n14050 ) ? ( VREG_8_13 ) : ( n14332 ) ;
assign n14334 =  ( n14049 ) ? ( VREG_8_14 ) : ( n14333 ) ;
assign n14335 =  ( n14048 ) ? ( VREG_8_15 ) : ( n14334 ) ;
assign n14336 =  ( n14047 ) ? ( VREG_9_0 ) : ( n14335 ) ;
assign n14337 =  ( n14046 ) ? ( VREG_9_1 ) : ( n14336 ) ;
assign n14338 =  ( n14045 ) ? ( VREG_9_2 ) : ( n14337 ) ;
assign n14339 =  ( n14044 ) ? ( VREG_9_3 ) : ( n14338 ) ;
assign n14340 =  ( n14043 ) ? ( VREG_9_4 ) : ( n14339 ) ;
assign n14341 =  ( n14042 ) ? ( VREG_9_5 ) : ( n14340 ) ;
assign n14342 =  ( n14041 ) ? ( VREG_9_6 ) : ( n14341 ) ;
assign n14343 =  ( n14040 ) ? ( VREG_9_7 ) : ( n14342 ) ;
assign n14344 =  ( n14039 ) ? ( VREG_9_8 ) : ( n14343 ) ;
assign n14345 =  ( n14038 ) ? ( VREG_9_9 ) : ( n14344 ) ;
assign n14346 =  ( n14037 ) ? ( VREG_9_10 ) : ( n14345 ) ;
assign n14347 =  ( n14036 ) ? ( VREG_9_11 ) : ( n14346 ) ;
assign n14348 =  ( n14035 ) ? ( VREG_9_12 ) : ( n14347 ) ;
assign n14349 =  ( n14034 ) ? ( VREG_9_13 ) : ( n14348 ) ;
assign n14350 =  ( n14033 ) ? ( VREG_9_14 ) : ( n14349 ) ;
assign n14351 =  ( n14032 ) ? ( VREG_9_15 ) : ( n14350 ) ;
assign n14352 =  ( n14031 ) ? ( VREG_10_0 ) : ( n14351 ) ;
assign n14353 =  ( n14030 ) ? ( VREG_10_1 ) : ( n14352 ) ;
assign n14354 =  ( n14029 ) ? ( VREG_10_2 ) : ( n14353 ) ;
assign n14355 =  ( n14028 ) ? ( VREG_10_3 ) : ( n14354 ) ;
assign n14356 =  ( n14027 ) ? ( VREG_10_4 ) : ( n14355 ) ;
assign n14357 =  ( n14026 ) ? ( VREG_10_5 ) : ( n14356 ) ;
assign n14358 =  ( n14025 ) ? ( VREG_10_6 ) : ( n14357 ) ;
assign n14359 =  ( n14024 ) ? ( VREG_10_7 ) : ( n14358 ) ;
assign n14360 =  ( n14023 ) ? ( VREG_10_8 ) : ( n14359 ) ;
assign n14361 =  ( n14022 ) ? ( VREG_10_9 ) : ( n14360 ) ;
assign n14362 =  ( n14021 ) ? ( VREG_10_10 ) : ( n14361 ) ;
assign n14363 =  ( n14020 ) ? ( VREG_10_11 ) : ( n14362 ) ;
assign n14364 =  ( n14019 ) ? ( VREG_10_12 ) : ( n14363 ) ;
assign n14365 =  ( n14018 ) ? ( VREG_10_13 ) : ( n14364 ) ;
assign n14366 =  ( n14017 ) ? ( VREG_10_14 ) : ( n14365 ) ;
assign n14367 =  ( n14016 ) ? ( VREG_10_15 ) : ( n14366 ) ;
assign n14368 =  ( n14015 ) ? ( VREG_11_0 ) : ( n14367 ) ;
assign n14369 =  ( n14014 ) ? ( VREG_11_1 ) : ( n14368 ) ;
assign n14370 =  ( n14013 ) ? ( VREG_11_2 ) : ( n14369 ) ;
assign n14371 =  ( n14012 ) ? ( VREG_11_3 ) : ( n14370 ) ;
assign n14372 =  ( n14011 ) ? ( VREG_11_4 ) : ( n14371 ) ;
assign n14373 =  ( n14010 ) ? ( VREG_11_5 ) : ( n14372 ) ;
assign n14374 =  ( n14009 ) ? ( VREG_11_6 ) : ( n14373 ) ;
assign n14375 =  ( n14008 ) ? ( VREG_11_7 ) : ( n14374 ) ;
assign n14376 =  ( n14007 ) ? ( VREG_11_8 ) : ( n14375 ) ;
assign n14377 =  ( n14006 ) ? ( VREG_11_9 ) : ( n14376 ) ;
assign n14378 =  ( n14005 ) ? ( VREG_11_10 ) : ( n14377 ) ;
assign n14379 =  ( n14004 ) ? ( VREG_11_11 ) : ( n14378 ) ;
assign n14380 =  ( n14003 ) ? ( VREG_11_12 ) : ( n14379 ) ;
assign n14381 =  ( n14002 ) ? ( VREG_11_13 ) : ( n14380 ) ;
assign n14382 =  ( n14001 ) ? ( VREG_11_14 ) : ( n14381 ) ;
assign n14383 =  ( n14000 ) ? ( VREG_11_15 ) : ( n14382 ) ;
assign n14384 =  ( n13999 ) ? ( VREG_12_0 ) : ( n14383 ) ;
assign n14385 =  ( n13998 ) ? ( VREG_12_1 ) : ( n14384 ) ;
assign n14386 =  ( n13997 ) ? ( VREG_12_2 ) : ( n14385 ) ;
assign n14387 =  ( n13996 ) ? ( VREG_12_3 ) : ( n14386 ) ;
assign n14388 =  ( n13995 ) ? ( VREG_12_4 ) : ( n14387 ) ;
assign n14389 =  ( n13994 ) ? ( VREG_12_5 ) : ( n14388 ) ;
assign n14390 =  ( n13993 ) ? ( VREG_12_6 ) : ( n14389 ) ;
assign n14391 =  ( n13992 ) ? ( VREG_12_7 ) : ( n14390 ) ;
assign n14392 =  ( n13991 ) ? ( VREG_12_8 ) : ( n14391 ) ;
assign n14393 =  ( n13990 ) ? ( VREG_12_9 ) : ( n14392 ) ;
assign n14394 =  ( n13989 ) ? ( VREG_12_10 ) : ( n14393 ) ;
assign n14395 =  ( n13988 ) ? ( VREG_12_11 ) : ( n14394 ) ;
assign n14396 =  ( n13987 ) ? ( VREG_12_12 ) : ( n14395 ) ;
assign n14397 =  ( n13986 ) ? ( VREG_12_13 ) : ( n14396 ) ;
assign n14398 =  ( n13985 ) ? ( VREG_12_14 ) : ( n14397 ) ;
assign n14399 =  ( n13984 ) ? ( VREG_12_15 ) : ( n14398 ) ;
assign n14400 =  ( n13983 ) ? ( VREG_13_0 ) : ( n14399 ) ;
assign n14401 =  ( n13982 ) ? ( VREG_13_1 ) : ( n14400 ) ;
assign n14402 =  ( n13981 ) ? ( VREG_13_2 ) : ( n14401 ) ;
assign n14403 =  ( n13980 ) ? ( VREG_13_3 ) : ( n14402 ) ;
assign n14404 =  ( n13979 ) ? ( VREG_13_4 ) : ( n14403 ) ;
assign n14405 =  ( n13978 ) ? ( VREG_13_5 ) : ( n14404 ) ;
assign n14406 =  ( n13977 ) ? ( VREG_13_6 ) : ( n14405 ) ;
assign n14407 =  ( n13976 ) ? ( VREG_13_7 ) : ( n14406 ) ;
assign n14408 =  ( n13975 ) ? ( VREG_13_8 ) : ( n14407 ) ;
assign n14409 =  ( n13974 ) ? ( VREG_13_9 ) : ( n14408 ) ;
assign n14410 =  ( n13973 ) ? ( VREG_13_10 ) : ( n14409 ) ;
assign n14411 =  ( n13972 ) ? ( VREG_13_11 ) : ( n14410 ) ;
assign n14412 =  ( n13971 ) ? ( VREG_13_12 ) : ( n14411 ) ;
assign n14413 =  ( n13970 ) ? ( VREG_13_13 ) : ( n14412 ) ;
assign n14414 =  ( n13969 ) ? ( VREG_13_14 ) : ( n14413 ) ;
assign n14415 =  ( n13968 ) ? ( VREG_13_15 ) : ( n14414 ) ;
assign n14416 =  ( n13967 ) ? ( VREG_14_0 ) : ( n14415 ) ;
assign n14417 =  ( n13966 ) ? ( VREG_14_1 ) : ( n14416 ) ;
assign n14418 =  ( n13965 ) ? ( VREG_14_2 ) : ( n14417 ) ;
assign n14419 =  ( n13964 ) ? ( VREG_14_3 ) : ( n14418 ) ;
assign n14420 =  ( n13963 ) ? ( VREG_14_4 ) : ( n14419 ) ;
assign n14421 =  ( n13962 ) ? ( VREG_14_5 ) : ( n14420 ) ;
assign n14422 =  ( n13961 ) ? ( VREG_14_6 ) : ( n14421 ) ;
assign n14423 =  ( n13960 ) ? ( VREG_14_7 ) : ( n14422 ) ;
assign n14424 =  ( n13959 ) ? ( VREG_14_8 ) : ( n14423 ) ;
assign n14425 =  ( n13958 ) ? ( VREG_14_9 ) : ( n14424 ) ;
assign n14426 =  ( n13957 ) ? ( VREG_14_10 ) : ( n14425 ) ;
assign n14427 =  ( n13956 ) ? ( VREG_14_11 ) : ( n14426 ) ;
assign n14428 =  ( n13955 ) ? ( VREG_14_12 ) : ( n14427 ) ;
assign n14429 =  ( n13954 ) ? ( VREG_14_13 ) : ( n14428 ) ;
assign n14430 =  ( n13953 ) ? ( VREG_14_14 ) : ( n14429 ) ;
assign n14431 =  ( n13952 ) ? ( VREG_14_15 ) : ( n14430 ) ;
assign n14432 =  ( n13951 ) ? ( VREG_15_0 ) : ( n14431 ) ;
assign n14433 =  ( n13950 ) ? ( VREG_15_1 ) : ( n14432 ) ;
assign n14434 =  ( n13949 ) ? ( VREG_15_2 ) : ( n14433 ) ;
assign n14435 =  ( n13948 ) ? ( VREG_15_3 ) : ( n14434 ) ;
assign n14436 =  ( n13947 ) ? ( VREG_15_4 ) : ( n14435 ) ;
assign n14437 =  ( n13946 ) ? ( VREG_15_5 ) : ( n14436 ) ;
assign n14438 =  ( n13945 ) ? ( VREG_15_6 ) : ( n14437 ) ;
assign n14439 =  ( n13944 ) ? ( VREG_15_7 ) : ( n14438 ) ;
assign n14440 =  ( n13943 ) ? ( VREG_15_8 ) : ( n14439 ) ;
assign n14441 =  ( n13942 ) ? ( VREG_15_9 ) : ( n14440 ) ;
assign n14442 =  ( n13941 ) ? ( VREG_15_10 ) : ( n14441 ) ;
assign n14443 =  ( n13940 ) ? ( VREG_15_11 ) : ( n14442 ) ;
assign n14444 =  ( n13939 ) ? ( VREG_15_12 ) : ( n14443 ) ;
assign n14445 =  ( n13938 ) ? ( VREG_15_13 ) : ( n14444 ) ;
assign n14446 =  ( n13937 ) ? ( VREG_15_14 ) : ( n14445 ) ;
assign n14447 =  ( n13936 ) ? ( VREG_15_15 ) : ( n14446 ) ;
assign n14448 =  ( n13935 ) ? ( VREG_16_0 ) : ( n14447 ) ;
assign n14449 =  ( n13934 ) ? ( VREG_16_1 ) : ( n14448 ) ;
assign n14450 =  ( n13933 ) ? ( VREG_16_2 ) : ( n14449 ) ;
assign n14451 =  ( n13932 ) ? ( VREG_16_3 ) : ( n14450 ) ;
assign n14452 =  ( n13931 ) ? ( VREG_16_4 ) : ( n14451 ) ;
assign n14453 =  ( n13930 ) ? ( VREG_16_5 ) : ( n14452 ) ;
assign n14454 =  ( n13929 ) ? ( VREG_16_6 ) : ( n14453 ) ;
assign n14455 =  ( n13928 ) ? ( VREG_16_7 ) : ( n14454 ) ;
assign n14456 =  ( n13927 ) ? ( VREG_16_8 ) : ( n14455 ) ;
assign n14457 =  ( n13926 ) ? ( VREG_16_9 ) : ( n14456 ) ;
assign n14458 =  ( n13925 ) ? ( VREG_16_10 ) : ( n14457 ) ;
assign n14459 =  ( n13924 ) ? ( VREG_16_11 ) : ( n14458 ) ;
assign n14460 =  ( n13923 ) ? ( VREG_16_12 ) : ( n14459 ) ;
assign n14461 =  ( n13922 ) ? ( VREG_16_13 ) : ( n14460 ) ;
assign n14462 =  ( n13921 ) ? ( VREG_16_14 ) : ( n14461 ) ;
assign n14463 =  ( n13920 ) ? ( VREG_16_15 ) : ( n14462 ) ;
assign n14464 =  ( n13919 ) ? ( VREG_17_0 ) : ( n14463 ) ;
assign n14465 =  ( n13918 ) ? ( VREG_17_1 ) : ( n14464 ) ;
assign n14466 =  ( n13917 ) ? ( VREG_17_2 ) : ( n14465 ) ;
assign n14467 =  ( n13916 ) ? ( VREG_17_3 ) : ( n14466 ) ;
assign n14468 =  ( n13915 ) ? ( VREG_17_4 ) : ( n14467 ) ;
assign n14469 =  ( n13914 ) ? ( VREG_17_5 ) : ( n14468 ) ;
assign n14470 =  ( n13913 ) ? ( VREG_17_6 ) : ( n14469 ) ;
assign n14471 =  ( n13912 ) ? ( VREG_17_7 ) : ( n14470 ) ;
assign n14472 =  ( n13911 ) ? ( VREG_17_8 ) : ( n14471 ) ;
assign n14473 =  ( n13910 ) ? ( VREG_17_9 ) : ( n14472 ) ;
assign n14474 =  ( n13909 ) ? ( VREG_17_10 ) : ( n14473 ) ;
assign n14475 =  ( n13908 ) ? ( VREG_17_11 ) : ( n14474 ) ;
assign n14476 =  ( n13907 ) ? ( VREG_17_12 ) : ( n14475 ) ;
assign n14477 =  ( n13906 ) ? ( VREG_17_13 ) : ( n14476 ) ;
assign n14478 =  ( n13905 ) ? ( VREG_17_14 ) : ( n14477 ) ;
assign n14479 =  ( n13904 ) ? ( VREG_17_15 ) : ( n14478 ) ;
assign n14480 =  ( n13903 ) ? ( VREG_18_0 ) : ( n14479 ) ;
assign n14481 =  ( n13902 ) ? ( VREG_18_1 ) : ( n14480 ) ;
assign n14482 =  ( n13901 ) ? ( VREG_18_2 ) : ( n14481 ) ;
assign n14483 =  ( n13900 ) ? ( VREG_18_3 ) : ( n14482 ) ;
assign n14484 =  ( n13899 ) ? ( VREG_18_4 ) : ( n14483 ) ;
assign n14485 =  ( n13898 ) ? ( VREG_18_5 ) : ( n14484 ) ;
assign n14486 =  ( n13897 ) ? ( VREG_18_6 ) : ( n14485 ) ;
assign n14487 =  ( n13896 ) ? ( VREG_18_7 ) : ( n14486 ) ;
assign n14488 =  ( n13895 ) ? ( VREG_18_8 ) : ( n14487 ) ;
assign n14489 =  ( n13894 ) ? ( VREG_18_9 ) : ( n14488 ) ;
assign n14490 =  ( n13893 ) ? ( VREG_18_10 ) : ( n14489 ) ;
assign n14491 =  ( n13892 ) ? ( VREG_18_11 ) : ( n14490 ) ;
assign n14492 =  ( n13891 ) ? ( VREG_18_12 ) : ( n14491 ) ;
assign n14493 =  ( n13890 ) ? ( VREG_18_13 ) : ( n14492 ) ;
assign n14494 =  ( n13889 ) ? ( VREG_18_14 ) : ( n14493 ) ;
assign n14495 =  ( n13888 ) ? ( VREG_18_15 ) : ( n14494 ) ;
assign n14496 =  ( n13887 ) ? ( VREG_19_0 ) : ( n14495 ) ;
assign n14497 =  ( n13886 ) ? ( VREG_19_1 ) : ( n14496 ) ;
assign n14498 =  ( n13885 ) ? ( VREG_19_2 ) : ( n14497 ) ;
assign n14499 =  ( n13884 ) ? ( VREG_19_3 ) : ( n14498 ) ;
assign n14500 =  ( n13883 ) ? ( VREG_19_4 ) : ( n14499 ) ;
assign n14501 =  ( n13882 ) ? ( VREG_19_5 ) : ( n14500 ) ;
assign n14502 =  ( n13881 ) ? ( VREG_19_6 ) : ( n14501 ) ;
assign n14503 =  ( n13880 ) ? ( VREG_19_7 ) : ( n14502 ) ;
assign n14504 =  ( n13879 ) ? ( VREG_19_8 ) : ( n14503 ) ;
assign n14505 =  ( n13878 ) ? ( VREG_19_9 ) : ( n14504 ) ;
assign n14506 =  ( n13877 ) ? ( VREG_19_10 ) : ( n14505 ) ;
assign n14507 =  ( n13876 ) ? ( VREG_19_11 ) : ( n14506 ) ;
assign n14508 =  ( n13875 ) ? ( VREG_19_12 ) : ( n14507 ) ;
assign n14509 =  ( n13874 ) ? ( VREG_19_13 ) : ( n14508 ) ;
assign n14510 =  ( n13873 ) ? ( VREG_19_14 ) : ( n14509 ) ;
assign n14511 =  ( n13872 ) ? ( VREG_19_15 ) : ( n14510 ) ;
assign n14512 =  ( n13871 ) ? ( VREG_20_0 ) : ( n14511 ) ;
assign n14513 =  ( n13870 ) ? ( VREG_20_1 ) : ( n14512 ) ;
assign n14514 =  ( n13869 ) ? ( VREG_20_2 ) : ( n14513 ) ;
assign n14515 =  ( n13868 ) ? ( VREG_20_3 ) : ( n14514 ) ;
assign n14516 =  ( n13867 ) ? ( VREG_20_4 ) : ( n14515 ) ;
assign n14517 =  ( n13866 ) ? ( VREG_20_5 ) : ( n14516 ) ;
assign n14518 =  ( n13865 ) ? ( VREG_20_6 ) : ( n14517 ) ;
assign n14519 =  ( n13864 ) ? ( VREG_20_7 ) : ( n14518 ) ;
assign n14520 =  ( n13863 ) ? ( VREG_20_8 ) : ( n14519 ) ;
assign n14521 =  ( n13862 ) ? ( VREG_20_9 ) : ( n14520 ) ;
assign n14522 =  ( n13861 ) ? ( VREG_20_10 ) : ( n14521 ) ;
assign n14523 =  ( n13860 ) ? ( VREG_20_11 ) : ( n14522 ) ;
assign n14524 =  ( n13859 ) ? ( VREG_20_12 ) : ( n14523 ) ;
assign n14525 =  ( n13858 ) ? ( VREG_20_13 ) : ( n14524 ) ;
assign n14526 =  ( n13857 ) ? ( VREG_20_14 ) : ( n14525 ) ;
assign n14527 =  ( n13856 ) ? ( VREG_20_15 ) : ( n14526 ) ;
assign n14528 =  ( n13855 ) ? ( VREG_21_0 ) : ( n14527 ) ;
assign n14529 =  ( n13854 ) ? ( VREG_21_1 ) : ( n14528 ) ;
assign n14530 =  ( n13853 ) ? ( VREG_21_2 ) : ( n14529 ) ;
assign n14531 =  ( n13852 ) ? ( VREG_21_3 ) : ( n14530 ) ;
assign n14532 =  ( n13851 ) ? ( VREG_21_4 ) : ( n14531 ) ;
assign n14533 =  ( n13850 ) ? ( VREG_21_5 ) : ( n14532 ) ;
assign n14534 =  ( n13849 ) ? ( VREG_21_6 ) : ( n14533 ) ;
assign n14535 =  ( n13848 ) ? ( VREG_21_7 ) : ( n14534 ) ;
assign n14536 =  ( n13847 ) ? ( VREG_21_8 ) : ( n14535 ) ;
assign n14537 =  ( n13846 ) ? ( VREG_21_9 ) : ( n14536 ) ;
assign n14538 =  ( n13845 ) ? ( VREG_21_10 ) : ( n14537 ) ;
assign n14539 =  ( n13844 ) ? ( VREG_21_11 ) : ( n14538 ) ;
assign n14540 =  ( n13843 ) ? ( VREG_21_12 ) : ( n14539 ) ;
assign n14541 =  ( n13842 ) ? ( VREG_21_13 ) : ( n14540 ) ;
assign n14542 =  ( n13841 ) ? ( VREG_21_14 ) : ( n14541 ) ;
assign n14543 =  ( n13840 ) ? ( VREG_21_15 ) : ( n14542 ) ;
assign n14544 =  ( n13839 ) ? ( VREG_22_0 ) : ( n14543 ) ;
assign n14545 =  ( n13838 ) ? ( VREG_22_1 ) : ( n14544 ) ;
assign n14546 =  ( n13837 ) ? ( VREG_22_2 ) : ( n14545 ) ;
assign n14547 =  ( n13836 ) ? ( VREG_22_3 ) : ( n14546 ) ;
assign n14548 =  ( n13835 ) ? ( VREG_22_4 ) : ( n14547 ) ;
assign n14549 =  ( n13834 ) ? ( VREG_22_5 ) : ( n14548 ) ;
assign n14550 =  ( n13833 ) ? ( VREG_22_6 ) : ( n14549 ) ;
assign n14551 =  ( n13832 ) ? ( VREG_22_7 ) : ( n14550 ) ;
assign n14552 =  ( n13831 ) ? ( VREG_22_8 ) : ( n14551 ) ;
assign n14553 =  ( n13830 ) ? ( VREG_22_9 ) : ( n14552 ) ;
assign n14554 =  ( n13829 ) ? ( VREG_22_10 ) : ( n14553 ) ;
assign n14555 =  ( n13828 ) ? ( VREG_22_11 ) : ( n14554 ) ;
assign n14556 =  ( n13827 ) ? ( VREG_22_12 ) : ( n14555 ) ;
assign n14557 =  ( n13826 ) ? ( VREG_22_13 ) : ( n14556 ) ;
assign n14558 =  ( n13825 ) ? ( VREG_22_14 ) : ( n14557 ) ;
assign n14559 =  ( n13824 ) ? ( VREG_22_15 ) : ( n14558 ) ;
assign n14560 =  ( n13823 ) ? ( VREG_23_0 ) : ( n14559 ) ;
assign n14561 =  ( n13822 ) ? ( VREG_23_1 ) : ( n14560 ) ;
assign n14562 =  ( n13821 ) ? ( VREG_23_2 ) : ( n14561 ) ;
assign n14563 =  ( n13820 ) ? ( VREG_23_3 ) : ( n14562 ) ;
assign n14564 =  ( n13819 ) ? ( VREG_23_4 ) : ( n14563 ) ;
assign n14565 =  ( n13818 ) ? ( VREG_23_5 ) : ( n14564 ) ;
assign n14566 =  ( n13817 ) ? ( VREG_23_6 ) : ( n14565 ) ;
assign n14567 =  ( n13816 ) ? ( VREG_23_7 ) : ( n14566 ) ;
assign n14568 =  ( n13815 ) ? ( VREG_23_8 ) : ( n14567 ) ;
assign n14569 =  ( n13814 ) ? ( VREG_23_9 ) : ( n14568 ) ;
assign n14570 =  ( n13813 ) ? ( VREG_23_10 ) : ( n14569 ) ;
assign n14571 =  ( n13812 ) ? ( VREG_23_11 ) : ( n14570 ) ;
assign n14572 =  ( n13811 ) ? ( VREG_23_12 ) : ( n14571 ) ;
assign n14573 =  ( n13810 ) ? ( VREG_23_13 ) : ( n14572 ) ;
assign n14574 =  ( n13809 ) ? ( VREG_23_14 ) : ( n14573 ) ;
assign n14575 =  ( n13808 ) ? ( VREG_23_15 ) : ( n14574 ) ;
assign n14576 =  ( n13807 ) ? ( VREG_24_0 ) : ( n14575 ) ;
assign n14577 =  ( n13806 ) ? ( VREG_24_1 ) : ( n14576 ) ;
assign n14578 =  ( n13805 ) ? ( VREG_24_2 ) : ( n14577 ) ;
assign n14579 =  ( n13804 ) ? ( VREG_24_3 ) : ( n14578 ) ;
assign n14580 =  ( n13803 ) ? ( VREG_24_4 ) : ( n14579 ) ;
assign n14581 =  ( n13802 ) ? ( VREG_24_5 ) : ( n14580 ) ;
assign n14582 =  ( n13801 ) ? ( VREG_24_6 ) : ( n14581 ) ;
assign n14583 =  ( n13800 ) ? ( VREG_24_7 ) : ( n14582 ) ;
assign n14584 =  ( n13799 ) ? ( VREG_24_8 ) : ( n14583 ) ;
assign n14585 =  ( n13798 ) ? ( VREG_24_9 ) : ( n14584 ) ;
assign n14586 =  ( n13797 ) ? ( VREG_24_10 ) : ( n14585 ) ;
assign n14587 =  ( n13796 ) ? ( VREG_24_11 ) : ( n14586 ) ;
assign n14588 =  ( n13795 ) ? ( VREG_24_12 ) : ( n14587 ) ;
assign n14589 =  ( n13794 ) ? ( VREG_24_13 ) : ( n14588 ) ;
assign n14590 =  ( n13793 ) ? ( VREG_24_14 ) : ( n14589 ) ;
assign n14591 =  ( n13792 ) ? ( VREG_24_15 ) : ( n14590 ) ;
assign n14592 =  ( n13791 ) ? ( VREG_25_0 ) : ( n14591 ) ;
assign n14593 =  ( n13790 ) ? ( VREG_25_1 ) : ( n14592 ) ;
assign n14594 =  ( n13789 ) ? ( VREG_25_2 ) : ( n14593 ) ;
assign n14595 =  ( n13788 ) ? ( VREG_25_3 ) : ( n14594 ) ;
assign n14596 =  ( n13787 ) ? ( VREG_25_4 ) : ( n14595 ) ;
assign n14597 =  ( n13786 ) ? ( VREG_25_5 ) : ( n14596 ) ;
assign n14598 =  ( n13785 ) ? ( VREG_25_6 ) : ( n14597 ) ;
assign n14599 =  ( n13784 ) ? ( VREG_25_7 ) : ( n14598 ) ;
assign n14600 =  ( n13783 ) ? ( VREG_25_8 ) : ( n14599 ) ;
assign n14601 =  ( n13782 ) ? ( VREG_25_9 ) : ( n14600 ) ;
assign n14602 =  ( n13781 ) ? ( VREG_25_10 ) : ( n14601 ) ;
assign n14603 =  ( n13780 ) ? ( VREG_25_11 ) : ( n14602 ) ;
assign n14604 =  ( n13779 ) ? ( VREG_25_12 ) : ( n14603 ) ;
assign n14605 =  ( n13778 ) ? ( VREG_25_13 ) : ( n14604 ) ;
assign n14606 =  ( n13777 ) ? ( VREG_25_14 ) : ( n14605 ) ;
assign n14607 =  ( n13776 ) ? ( VREG_25_15 ) : ( n14606 ) ;
assign n14608 =  ( n13775 ) ? ( VREG_26_0 ) : ( n14607 ) ;
assign n14609 =  ( n13774 ) ? ( VREG_26_1 ) : ( n14608 ) ;
assign n14610 =  ( n13773 ) ? ( VREG_26_2 ) : ( n14609 ) ;
assign n14611 =  ( n13772 ) ? ( VREG_26_3 ) : ( n14610 ) ;
assign n14612 =  ( n13771 ) ? ( VREG_26_4 ) : ( n14611 ) ;
assign n14613 =  ( n13770 ) ? ( VREG_26_5 ) : ( n14612 ) ;
assign n14614 =  ( n13769 ) ? ( VREG_26_6 ) : ( n14613 ) ;
assign n14615 =  ( n13768 ) ? ( VREG_26_7 ) : ( n14614 ) ;
assign n14616 =  ( n13767 ) ? ( VREG_26_8 ) : ( n14615 ) ;
assign n14617 =  ( n13766 ) ? ( VREG_26_9 ) : ( n14616 ) ;
assign n14618 =  ( n13765 ) ? ( VREG_26_10 ) : ( n14617 ) ;
assign n14619 =  ( n13764 ) ? ( VREG_26_11 ) : ( n14618 ) ;
assign n14620 =  ( n13763 ) ? ( VREG_26_12 ) : ( n14619 ) ;
assign n14621 =  ( n13762 ) ? ( VREG_26_13 ) : ( n14620 ) ;
assign n14622 =  ( n13761 ) ? ( VREG_26_14 ) : ( n14621 ) ;
assign n14623 =  ( n13760 ) ? ( VREG_26_15 ) : ( n14622 ) ;
assign n14624 =  ( n13759 ) ? ( VREG_27_0 ) : ( n14623 ) ;
assign n14625 =  ( n13758 ) ? ( VREG_27_1 ) : ( n14624 ) ;
assign n14626 =  ( n13757 ) ? ( VREG_27_2 ) : ( n14625 ) ;
assign n14627 =  ( n13756 ) ? ( VREG_27_3 ) : ( n14626 ) ;
assign n14628 =  ( n13755 ) ? ( VREG_27_4 ) : ( n14627 ) ;
assign n14629 =  ( n13754 ) ? ( VREG_27_5 ) : ( n14628 ) ;
assign n14630 =  ( n13753 ) ? ( VREG_27_6 ) : ( n14629 ) ;
assign n14631 =  ( n13752 ) ? ( VREG_27_7 ) : ( n14630 ) ;
assign n14632 =  ( n13751 ) ? ( VREG_27_8 ) : ( n14631 ) ;
assign n14633 =  ( n13750 ) ? ( VREG_27_9 ) : ( n14632 ) ;
assign n14634 =  ( n13749 ) ? ( VREG_27_10 ) : ( n14633 ) ;
assign n14635 =  ( n13748 ) ? ( VREG_27_11 ) : ( n14634 ) ;
assign n14636 =  ( n13747 ) ? ( VREG_27_12 ) : ( n14635 ) ;
assign n14637 =  ( n13746 ) ? ( VREG_27_13 ) : ( n14636 ) ;
assign n14638 =  ( n13745 ) ? ( VREG_27_14 ) : ( n14637 ) ;
assign n14639 =  ( n13744 ) ? ( VREG_27_15 ) : ( n14638 ) ;
assign n14640 =  ( n13743 ) ? ( VREG_28_0 ) : ( n14639 ) ;
assign n14641 =  ( n13742 ) ? ( VREG_28_1 ) : ( n14640 ) ;
assign n14642 =  ( n13741 ) ? ( VREG_28_2 ) : ( n14641 ) ;
assign n14643 =  ( n13740 ) ? ( VREG_28_3 ) : ( n14642 ) ;
assign n14644 =  ( n13739 ) ? ( VREG_28_4 ) : ( n14643 ) ;
assign n14645 =  ( n13738 ) ? ( VREG_28_5 ) : ( n14644 ) ;
assign n14646 =  ( n13737 ) ? ( VREG_28_6 ) : ( n14645 ) ;
assign n14647 =  ( n13736 ) ? ( VREG_28_7 ) : ( n14646 ) ;
assign n14648 =  ( n13735 ) ? ( VREG_28_8 ) : ( n14647 ) ;
assign n14649 =  ( n13734 ) ? ( VREG_28_9 ) : ( n14648 ) ;
assign n14650 =  ( n13733 ) ? ( VREG_28_10 ) : ( n14649 ) ;
assign n14651 =  ( n13732 ) ? ( VREG_28_11 ) : ( n14650 ) ;
assign n14652 =  ( n13731 ) ? ( VREG_28_12 ) : ( n14651 ) ;
assign n14653 =  ( n13730 ) ? ( VREG_28_13 ) : ( n14652 ) ;
assign n14654 =  ( n13729 ) ? ( VREG_28_14 ) : ( n14653 ) ;
assign n14655 =  ( n13728 ) ? ( VREG_28_15 ) : ( n14654 ) ;
assign n14656 =  ( n13727 ) ? ( VREG_29_0 ) : ( n14655 ) ;
assign n14657 =  ( n13726 ) ? ( VREG_29_1 ) : ( n14656 ) ;
assign n14658 =  ( n13725 ) ? ( VREG_29_2 ) : ( n14657 ) ;
assign n14659 =  ( n13724 ) ? ( VREG_29_3 ) : ( n14658 ) ;
assign n14660 =  ( n13723 ) ? ( VREG_29_4 ) : ( n14659 ) ;
assign n14661 =  ( n13722 ) ? ( VREG_29_5 ) : ( n14660 ) ;
assign n14662 =  ( n13721 ) ? ( VREG_29_6 ) : ( n14661 ) ;
assign n14663 =  ( n13720 ) ? ( VREG_29_7 ) : ( n14662 ) ;
assign n14664 =  ( n13719 ) ? ( VREG_29_8 ) : ( n14663 ) ;
assign n14665 =  ( n13718 ) ? ( VREG_29_9 ) : ( n14664 ) ;
assign n14666 =  ( n13717 ) ? ( VREG_29_10 ) : ( n14665 ) ;
assign n14667 =  ( n13716 ) ? ( VREG_29_11 ) : ( n14666 ) ;
assign n14668 =  ( n13715 ) ? ( VREG_29_12 ) : ( n14667 ) ;
assign n14669 =  ( n13714 ) ? ( VREG_29_13 ) : ( n14668 ) ;
assign n14670 =  ( n13713 ) ? ( VREG_29_14 ) : ( n14669 ) ;
assign n14671 =  ( n13712 ) ? ( VREG_29_15 ) : ( n14670 ) ;
assign n14672 =  ( n13711 ) ? ( VREG_30_0 ) : ( n14671 ) ;
assign n14673 =  ( n13710 ) ? ( VREG_30_1 ) : ( n14672 ) ;
assign n14674 =  ( n13709 ) ? ( VREG_30_2 ) : ( n14673 ) ;
assign n14675 =  ( n13708 ) ? ( VREG_30_3 ) : ( n14674 ) ;
assign n14676 =  ( n13707 ) ? ( VREG_30_4 ) : ( n14675 ) ;
assign n14677 =  ( n13706 ) ? ( VREG_30_5 ) : ( n14676 ) ;
assign n14678 =  ( n13705 ) ? ( VREG_30_6 ) : ( n14677 ) ;
assign n14679 =  ( n13704 ) ? ( VREG_30_7 ) : ( n14678 ) ;
assign n14680 =  ( n13703 ) ? ( VREG_30_8 ) : ( n14679 ) ;
assign n14681 =  ( n13702 ) ? ( VREG_30_9 ) : ( n14680 ) ;
assign n14682 =  ( n13701 ) ? ( VREG_30_10 ) : ( n14681 ) ;
assign n14683 =  ( n13700 ) ? ( VREG_30_11 ) : ( n14682 ) ;
assign n14684 =  ( n13699 ) ? ( VREG_30_12 ) : ( n14683 ) ;
assign n14685 =  ( n13698 ) ? ( VREG_30_13 ) : ( n14684 ) ;
assign n14686 =  ( n13697 ) ? ( VREG_30_14 ) : ( n14685 ) ;
assign n14687 =  ( n13696 ) ? ( VREG_30_15 ) : ( n14686 ) ;
assign n14688 =  ( n13695 ) ? ( VREG_31_0 ) : ( n14687 ) ;
assign n14689 =  ( n13693 ) ? ( VREG_31_1 ) : ( n14688 ) ;
assign n14690 =  ( n13691 ) ? ( VREG_31_2 ) : ( n14689 ) ;
assign n14691 =  ( n13689 ) ? ( VREG_31_3 ) : ( n14690 ) ;
assign n14692 =  ( n13687 ) ? ( VREG_31_4 ) : ( n14691 ) ;
assign n14693 =  ( n13685 ) ? ( VREG_31_5 ) : ( n14692 ) ;
assign n14694 =  ( n13683 ) ? ( VREG_31_6 ) : ( n14693 ) ;
assign n14695 =  ( n13681 ) ? ( VREG_31_7 ) : ( n14694 ) ;
assign n14696 =  ( n13679 ) ? ( VREG_31_8 ) : ( n14695 ) ;
assign n14697 =  ( n13677 ) ? ( VREG_31_9 ) : ( n14696 ) ;
assign n14698 =  ( n13675 ) ? ( VREG_31_10 ) : ( n14697 ) ;
assign n14699 =  ( n13673 ) ? ( VREG_31_11 ) : ( n14698 ) ;
assign n14700 =  ( n13671 ) ? ( VREG_31_12 ) : ( n14699 ) ;
assign n14701 =  ( n13669 ) ? ( VREG_31_13 ) : ( n14700 ) ;
assign n14702 =  ( n13667 ) ? ( VREG_31_14 ) : ( n14701 ) ;
assign n14703 =  ( n13665 ) ? ( VREG_31_15 ) : ( n14702 ) ;
assign n14704 =  ( n14703 ) + ( n140 )  ;
assign n14705 =  ( n14703 ) - ( n140 )  ;
assign n14706 =  ( n14703 ) & ( n140 )  ;
assign n14707 =  ( n14703 ) | ( n140 )  ;
assign n14708 =  ( ( n14703 ) * ( n140 ))  ;
assign n14709 =  ( n148 ) ? ( n14708 ) : ( VREG_0_14 ) ;
assign n14710 =  ( n146 ) ? ( n14707 ) : ( n14709 ) ;
assign n14711 =  ( n144 ) ? ( n14706 ) : ( n14710 ) ;
assign n14712 =  ( n142 ) ? ( n14705 ) : ( n14711 ) ;
assign n14713 =  ( n10 ) ? ( n14704 ) : ( n14712 ) ;
assign n14714 =  ( n77 ) & ( n13664 )  ;
assign n14715 =  ( n77 ) & ( n13666 )  ;
assign n14716 =  ( n77 ) & ( n13668 )  ;
assign n14717 =  ( n77 ) & ( n13670 )  ;
assign n14718 =  ( n77 ) & ( n13672 )  ;
assign n14719 =  ( n77 ) & ( n13674 )  ;
assign n14720 =  ( n77 ) & ( n13676 )  ;
assign n14721 =  ( n77 ) & ( n13678 )  ;
assign n14722 =  ( n77 ) & ( n13680 )  ;
assign n14723 =  ( n77 ) & ( n13682 )  ;
assign n14724 =  ( n77 ) & ( n13684 )  ;
assign n14725 =  ( n77 ) & ( n13686 )  ;
assign n14726 =  ( n77 ) & ( n13688 )  ;
assign n14727 =  ( n77 ) & ( n13690 )  ;
assign n14728 =  ( n77 ) & ( n13692 )  ;
assign n14729 =  ( n77 ) & ( n13694 )  ;
assign n14730 =  ( n78 ) & ( n13664 )  ;
assign n14731 =  ( n78 ) & ( n13666 )  ;
assign n14732 =  ( n78 ) & ( n13668 )  ;
assign n14733 =  ( n78 ) & ( n13670 )  ;
assign n14734 =  ( n78 ) & ( n13672 )  ;
assign n14735 =  ( n78 ) & ( n13674 )  ;
assign n14736 =  ( n78 ) & ( n13676 )  ;
assign n14737 =  ( n78 ) & ( n13678 )  ;
assign n14738 =  ( n78 ) & ( n13680 )  ;
assign n14739 =  ( n78 ) & ( n13682 )  ;
assign n14740 =  ( n78 ) & ( n13684 )  ;
assign n14741 =  ( n78 ) & ( n13686 )  ;
assign n14742 =  ( n78 ) & ( n13688 )  ;
assign n14743 =  ( n78 ) & ( n13690 )  ;
assign n14744 =  ( n78 ) & ( n13692 )  ;
assign n14745 =  ( n78 ) & ( n13694 )  ;
assign n14746 =  ( n79 ) & ( n13664 )  ;
assign n14747 =  ( n79 ) & ( n13666 )  ;
assign n14748 =  ( n79 ) & ( n13668 )  ;
assign n14749 =  ( n79 ) & ( n13670 )  ;
assign n14750 =  ( n79 ) & ( n13672 )  ;
assign n14751 =  ( n79 ) & ( n13674 )  ;
assign n14752 =  ( n79 ) & ( n13676 )  ;
assign n14753 =  ( n79 ) & ( n13678 )  ;
assign n14754 =  ( n79 ) & ( n13680 )  ;
assign n14755 =  ( n79 ) & ( n13682 )  ;
assign n14756 =  ( n79 ) & ( n13684 )  ;
assign n14757 =  ( n79 ) & ( n13686 )  ;
assign n14758 =  ( n79 ) & ( n13688 )  ;
assign n14759 =  ( n79 ) & ( n13690 )  ;
assign n14760 =  ( n79 ) & ( n13692 )  ;
assign n14761 =  ( n79 ) & ( n13694 )  ;
assign n14762 =  ( n80 ) & ( n13664 )  ;
assign n14763 =  ( n80 ) & ( n13666 )  ;
assign n14764 =  ( n80 ) & ( n13668 )  ;
assign n14765 =  ( n80 ) & ( n13670 )  ;
assign n14766 =  ( n80 ) & ( n13672 )  ;
assign n14767 =  ( n80 ) & ( n13674 )  ;
assign n14768 =  ( n80 ) & ( n13676 )  ;
assign n14769 =  ( n80 ) & ( n13678 )  ;
assign n14770 =  ( n80 ) & ( n13680 )  ;
assign n14771 =  ( n80 ) & ( n13682 )  ;
assign n14772 =  ( n80 ) & ( n13684 )  ;
assign n14773 =  ( n80 ) & ( n13686 )  ;
assign n14774 =  ( n80 ) & ( n13688 )  ;
assign n14775 =  ( n80 ) & ( n13690 )  ;
assign n14776 =  ( n80 ) & ( n13692 )  ;
assign n14777 =  ( n80 ) & ( n13694 )  ;
assign n14778 =  ( n81 ) & ( n13664 )  ;
assign n14779 =  ( n81 ) & ( n13666 )  ;
assign n14780 =  ( n81 ) & ( n13668 )  ;
assign n14781 =  ( n81 ) & ( n13670 )  ;
assign n14782 =  ( n81 ) & ( n13672 )  ;
assign n14783 =  ( n81 ) & ( n13674 )  ;
assign n14784 =  ( n81 ) & ( n13676 )  ;
assign n14785 =  ( n81 ) & ( n13678 )  ;
assign n14786 =  ( n81 ) & ( n13680 )  ;
assign n14787 =  ( n81 ) & ( n13682 )  ;
assign n14788 =  ( n81 ) & ( n13684 )  ;
assign n14789 =  ( n81 ) & ( n13686 )  ;
assign n14790 =  ( n81 ) & ( n13688 )  ;
assign n14791 =  ( n81 ) & ( n13690 )  ;
assign n14792 =  ( n81 ) & ( n13692 )  ;
assign n14793 =  ( n81 ) & ( n13694 )  ;
assign n14794 =  ( n82 ) & ( n13664 )  ;
assign n14795 =  ( n82 ) & ( n13666 )  ;
assign n14796 =  ( n82 ) & ( n13668 )  ;
assign n14797 =  ( n82 ) & ( n13670 )  ;
assign n14798 =  ( n82 ) & ( n13672 )  ;
assign n14799 =  ( n82 ) & ( n13674 )  ;
assign n14800 =  ( n82 ) & ( n13676 )  ;
assign n14801 =  ( n82 ) & ( n13678 )  ;
assign n14802 =  ( n82 ) & ( n13680 )  ;
assign n14803 =  ( n82 ) & ( n13682 )  ;
assign n14804 =  ( n82 ) & ( n13684 )  ;
assign n14805 =  ( n82 ) & ( n13686 )  ;
assign n14806 =  ( n82 ) & ( n13688 )  ;
assign n14807 =  ( n82 ) & ( n13690 )  ;
assign n14808 =  ( n82 ) & ( n13692 )  ;
assign n14809 =  ( n82 ) & ( n13694 )  ;
assign n14810 =  ( n83 ) & ( n13664 )  ;
assign n14811 =  ( n83 ) & ( n13666 )  ;
assign n14812 =  ( n83 ) & ( n13668 )  ;
assign n14813 =  ( n83 ) & ( n13670 )  ;
assign n14814 =  ( n83 ) & ( n13672 )  ;
assign n14815 =  ( n83 ) & ( n13674 )  ;
assign n14816 =  ( n83 ) & ( n13676 )  ;
assign n14817 =  ( n83 ) & ( n13678 )  ;
assign n14818 =  ( n83 ) & ( n13680 )  ;
assign n14819 =  ( n83 ) & ( n13682 )  ;
assign n14820 =  ( n83 ) & ( n13684 )  ;
assign n14821 =  ( n83 ) & ( n13686 )  ;
assign n14822 =  ( n83 ) & ( n13688 )  ;
assign n14823 =  ( n83 ) & ( n13690 )  ;
assign n14824 =  ( n83 ) & ( n13692 )  ;
assign n14825 =  ( n83 ) & ( n13694 )  ;
assign n14826 =  ( n84 ) & ( n13664 )  ;
assign n14827 =  ( n84 ) & ( n13666 )  ;
assign n14828 =  ( n84 ) & ( n13668 )  ;
assign n14829 =  ( n84 ) & ( n13670 )  ;
assign n14830 =  ( n84 ) & ( n13672 )  ;
assign n14831 =  ( n84 ) & ( n13674 )  ;
assign n14832 =  ( n84 ) & ( n13676 )  ;
assign n14833 =  ( n84 ) & ( n13678 )  ;
assign n14834 =  ( n84 ) & ( n13680 )  ;
assign n14835 =  ( n84 ) & ( n13682 )  ;
assign n14836 =  ( n84 ) & ( n13684 )  ;
assign n14837 =  ( n84 ) & ( n13686 )  ;
assign n14838 =  ( n84 ) & ( n13688 )  ;
assign n14839 =  ( n84 ) & ( n13690 )  ;
assign n14840 =  ( n84 ) & ( n13692 )  ;
assign n14841 =  ( n84 ) & ( n13694 )  ;
assign n14842 =  ( n85 ) & ( n13664 )  ;
assign n14843 =  ( n85 ) & ( n13666 )  ;
assign n14844 =  ( n85 ) & ( n13668 )  ;
assign n14845 =  ( n85 ) & ( n13670 )  ;
assign n14846 =  ( n85 ) & ( n13672 )  ;
assign n14847 =  ( n85 ) & ( n13674 )  ;
assign n14848 =  ( n85 ) & ( n13676 )  ;
assign n14849 =  ( n85 ) & ( n13678 )  ;
assign n14850 =  ( n85 ) & ( n13680 )  ;
assign n14851 =  ( n85 ) & ( n13682 )  ;
assign n14852 =  ( n85 ) & ( n13684 )  ;
assign n14853 =  ( n85 ) & ( n13686 )  ;
assign n14854 =  ( n85 ) & ( n13688 )  ;
assign n14855 =  ( n85 ) & ( n13690 )  ;
assign n14856 =  ( n85 ) & ( n13692 )  ;
assign n14857 =  ( n85 ) & ( n13694 )  ;
assign n14858 =  ( n86 ) & ( n13664 )  ;
assign n14859 =  ( n86 ) & ( n13666 )  ;
assign n14860 =  ( n86 ) & ( n13668 )  ;
assign n14861 =  ( n86 ) & ( n13670 )  ;
assign n14862 =  ( n86 ) & ( n13672 )  ;
assign n14863 =  ( n86 ) & ( n13674 )  ;
assign n14864 =  ( n86 ) & ( n13676 )  ;
assign n14865 =  ( n86 ) & ( n13678 )  ;
assign n14866 =  ( n86 ) & ( n13680 )  ;
assign n14867 =  ( n86 ) & ( n13682 )  ;
assign n14868 =  ( n86 ) & ( n13684 )  ;
assign n14869 =  ( n86 ) & ( n13686 )  ;
assign n14870 =  ( n86 ) & ( n13688 )  ;
assign n14871 =  ( n86 ) & ( n13690 )  ;
assign n14872 =  ( n86 ) & ( n13692 )  ;
assign n14873 =  ( n86 ) & ( n13694 )  ;
assign n14874 =  ( n87 ) & ( n13664 )  ;
assign n14875 =  ( n87 ) & ( n13666 )  ;
assign n14876 =  ( n87 ) & ( n13668 )  ;
assign n14877 =  ( n87 ) & ( n13670 )  ;
assign n14878 =  ( n87 ) & ( n13672 )  ;
assign n14879 =  ( n87 ) & ( n13674 )  ;
assign n14880 =  ( n87 ) & ( n13676 )  ;
assign n14881 =  ( n87 ) & ( n13678 )  ;
assign n14882 =  ( n87 ) & ( n13680 )  ;
assign n14883 =  ( n87 ) & ( n13682 )  ;
assign n14884 =  ( n87 ) & ( n13684 )  ;
assign n14885 =  ( n87 ) & ( n13686 )  ;
assign n14886 =  ( n87 ) & ( n13688 )  ;
assign n14887 =  ( n87 ) & ( n13690 )  ;
assign n14888 =  ( n87 ) & ( n13692 )  ;
assign n14889 =  ( n87 ) & ( n13694 )  ;
assign n14890 =  ( n88 ) & ( n13664 )  ;
assign n14891 =  ( n88 ) & ( n13666 )  ;
assign n14892 =  ( n88 ) & ( n13668 )  ;
assign n14893 =  ( n88 ) & ( n13670 )  ;
assign n14894 =  ( n88 ) & ( n13672 )  ;
assign n14895 =  ( n88 ) & ( n13674 )  ;
assign n14896 =  ( n88 ) & ( n13676 )  ;
assign n14897 =  ( n88 ) & ( n13678 )  ;
assign n14898 =  ( n88 ) & ( n13680 )  ;
assign n14899 =  ( n88 ) & ( n13682 )  ;
assign n14900 =  ( n88 ) & ( n13684 )  ;
assign n14901 =  ( n88 ) & ( n13686 )  ;
assign n14902 =  ( n88 ) & ( n13688 )  ;
assign n14903 =  ( n88 ) & ( n13690 )  ;
assign n14904 =  ( n88 ) & ( n13692 )  ;
assign n14905 =  ( n88 ) & ( n13694 )  ;
assign n14906 =  ( n89 ) & ( n13664 )  ;
assign n14907 =  ( n89 ) & ( n13666 )  ;
assign n14908 =  ( n89 ) & ( n13668 )  ;
assign n14909 =  ( n89 ) & ( n13670 )  ;
assign n14910 =  ( n89 ) & ( n13672 )  ;
assign n14911 =  ( n89 ) & ( n13674 )  ;
assign n14912 =  ( n89 ) & ( n13676 )  ;
assign n14913 =  ( n89 ) & ( n13678 )  ;
assign n14914 =  ( n89 ) & ( n13680 )  ;
assign n14915 =  ( n89 ) & ( n13682 )  ;
assign n14916 =  ( n89 ) & ( n13684 )  ;
assign n14917 =  ( n89 ) & ( n13686 )  ;
assign n14918 =  ( n89 ) & ( n13688 )  ;
assign n14919 =  ( n89 ) & ( n13690 )  ;
assign n14920 =  ( n89 ) & ( n13692 )  ;
assign n14921 =  ( n89 ) & ( n13694 )  ;
assign n14922 =  ( n90 ) & ( n13664 )  ;
assign n14923 =  ( n90 ) & ( n13666 )  ;
assign n14924 =  ( n90 ) & ( n13668 )  ;
assign n14925 =  ( n90 ) & ( n13670 )  ;
assign n14926 =  ( n90 ) & ( n13672 )  ;
assign n14927 =  ( n90 ) & ( n13674 )  ;
assign n14928 =  ( n90 ) & ( n13676 )  ;
assign n14929 =  ( n90 ) & ( n13678 )  ;
assign n14930 =  ( n90 ) & ( n13680 )  ;
assign n14931 =  ( n90 ) & ( n13682 )  ;
assign n14932 =  ( n90 ) & ( n13684 )  ;
assign n14933 =  ( n90 ) & ( n13686 )  ;
assign n14934 =  ( n90 ) & ( n13688 )  ;
assign n14935 =  ( n90 ) & ( n13690 )  ;
assign n14936 =  ( n90 ) & ( n13692 )  ;
assign n14937 =  ( n90 ) & ( n13694 )  ;
assign n14938 =  ( n91 ) & ( n13664 )  ;
assign n14939 =  ( n91 ) & ( n13666 )  ;
assign n14940 =  ( n91 ) & ( n13668 )  ;
assign n14941 =  ( n91 ) & ( n13670 )  ;
assign n14942 =  ( n91 ) & ( n13672 )  ;
assign n14943 =  ( n91 ) & ( n13674 )  ;
assign n14944 =  ( n91 ) & ( n13676 )  ;
assign n14945 =  ( n91 ) & ( n13678 )  ;
assign n14946 =  ( n91 ) & ( n13680 )  ;
assign n14947 =  ( n91 ) & ( n13682 )  ;
assign n14948 =  ( n91 ) & ( n13684 )  ;
assign n14949 =  ( n91 ) & ( n13686 )  ;
assign n14950 =  ( n91 ) & ( n13688 )  ;
assign n14951 =  ( n91 ) & ( n13690 )  ;
assign n14952 =  ( n91 ) & ( n13692 )  ;
assign n14953 =  ( n91 ) & ( n13694 )  ;
assign n14954 =  ( n92 ) & ( n13664 )  ;
assign n14955 =  ( n92 ) & ( n13666 )  ;
assign n14956 =  ( n92 ) & ( n13668 )  ;
assign n14957 =  ( n92 ) & ( n13670 )  ;
assign n14958 =  ( n92 ) & ( n13672 )  ;
assign n14959 =  ( n92 ) & ( n13674 )  ;
assign n14960 =  ( n92 ) & ( n13676 )  ;
assign n14961 =  ( n92 ) & ( n13678 )  ;
assign n14962 =  ( n92 ) & ( n13680 )  ;
assign n14963 =  ( n92 ) & ( n13682 )  ;
assign n14964 =  ( n92 ) & ( n13684 )  ;
assign n14965 =  ( n92 ) & ( n13686 )  ;
assign n14966 =  ( n92 ) & ( n13688 )  ;
assign n14967 =  ( n92 ) & ( n13690 )  ;
assign n14968 =  ( n92 ) & ( n13692 )  ;
assign n14969 =  ( n92 ) & ( n13694 )  ;
assign n14970 =  ( n93 ) & ( n13664 )  ;
assign n14971 =  ( n93 ) & ( n13666 )  ;
assign n14972 =  ( n93 ) & ( n13668 )  ;
assign n14973 =  ( n93 ) & ( n13670 )  ;
assign n14974 =  ( n93 ) & ( n13672 )  ;
assign n14975 =  ( n93 ) & ( n13674 )  ;
assign n14976 =  ( n93 ) & ( n13676 )  ;
assign n14977 =  ( n93 ) & ( n13678 )  ;
assign n14978 =  ( n93 ) & ( n13680 )  ;
assign n14979 =  ( n93 ) & ( n13682 )  ;
assign n14980 =  ( n93 ) & ( n13684 )  ;
assign n14981 =  ( n93 ) & ( n13686 )  ;
assign n14982 =  ( n93 ) & ( n13688 )  ;
assign n14983 =  ( n93 ) & ( n13690 )  ;
assign n14984 =  ( n93 ) & ( n13692 )  ;
assign n14985 =  ( n93 ) & ( n13694 )  ;
assign n14986 =  ( n94 ) & ( n13664 )  ;
assign n14987 =  ( n94 ) & ( n13666 )  ;
assign n14988 =  ( n94 ) & ( n13668 )  ;
assign n14989 =  ( n94 ) & ( n13670 )  ;
assign n14990 =  ( n94 ) & ( n13672 )  ;
assign n14991 =  ( n94 ) & ( n13674 )  ;
assign n14992 =  ( n94 ) & ( n13676 )  ;
assign n14993 =  ( n94 ) & ( n13678 )  ;
assign n14994 =  ( n94 ) & ( n13680 )  ;
assign n14995 =  ( n94 ) & ( n13682 )  ;
assign n14996 =  ( n94 ) & ( n13684 )  ;
assign n14997 =  ( n94 ) & ( n13686 )  ;
assign n14998 =  ( n94 ) & ( n13688 )  ;
assign n14999 =  ( n94 ) & ( n13690 )  ;
assign n15000 =  ( n94 ) & ( n13692 )  ;
assign n15001 =  ( n94 ) & ( n13694 )  ;
assign n15002 =  ( n95 ) & ( n13664 )  ;
assign n15003 =  ( n95 ) & ( n13666 )  ;
assign n15004 =  ( n95 ) & ( n13668 )  ;
assign n15005 =  ( n95 ) & ( n13670 )  ;
assign n15006 =  ( n95 ) & ( n13672 )  ;
assign n15007 =  ( n95 ) & ( n13674 )  ;
assign n15008 =  ( n95 ) & ( n13676 )  ;
assign n15009 =  ( n95 ) & ( n13678 )  ;
assign n15010 =  ( n95 ) & ( n13680 )  ;
assign n15011 =  ( n95 ) & ( n13682 )  ;
assign n15012 =  ( n95 ) & ( n13684 )  ;
assign n15013 =  ( n95 ) & ( n13686 )  ;
assign n15014 =  ( n95 ) & ( n13688 )  ;
assign n15015 =  ( n95 ) & ( n13690 )  ;
assign n15016 =  ( n95 ) & ( n13692 )  ;
assign n15017 =  ( n95 ) & ( n13694 )  ;
assign n15018 =  ( n96 ) & ( n13664 )  ;
assign n15019 =  ( n96 ) & ( n13666 )  ;
assign n15020 =  ( n96 ) & ( n13668 )  ;
assign n15021 =  ( n96 ) & ( n13670 )  ;
assign n15022 =  ( n96 ) & ( n13672 )  ;
assign n15023 =  ( n96 ) & ( n13674 )  ;
assign n15024 =  ( n96 ) & ( n13676 )  ;
assign n15025 =  ( n96 ) & ( n13678 )  ;
assign n15026 =  ( n96 ) & ( n13680 )  ;
assign n15027 =  ( n96 ) & ( n13682 )  ;
assign n15028 =  ( n96 ) & ( n13684 )  ;
assign n15029 =  ( n96 ) & ( n13686 )  ;
assign n15030 =  ( n96 ) & ( n13688 )  ;
assign n15031 =  ( n96 ) & ( n13690 )  ;
assign n15032 =  ( n96 ) & ( n13692 )  ;
assign n15033 =  ( n96 ) & ( n13694 )  ;
assign n15034 =  ( n97 ) & ( n13664 )  ;
assign n15035 =  ( n97 ) & ( n13666 )  ;
assign n15036 =  ( n97 ) & ( n13668 )  ;
assign n15037 =  ( n97 ) & ( n13670 )  ;
assign n15038 =  ( n97 ) & ( n13672 )  ;
assign n15039 =  ( n97 ) & ( n13674 )  ;
assign n15040 =  ( n97 ) & ( n13676 )  ;
assign n15041 =  ( n97 ) & ( n13678 )  ;
assign n15042 =  ( n97 ) & ( n13680 )  ;
assign n15043 =  ( n97 ) & ( n13682 )  ;
assign n15044 =  ( n97 ) & ( n13684 )  ;
assign n15045 =  ( n97 ) & ( n13686 )  ;
assign n15046 =  ( n97 ) & ( n13688 )  ;
assign n15047 =  ( n97 ) & ( n13690 )  ;
assign n15048 =  ( n97 ) & ( n13692 )  ;
assign n15049 =  ( n97 ) & ( n13694 )  ;
assign n15050 =  ( n98 ) & ( n13664 )  ;
assign n15051 =  ( n98 ) & ( n13666 )  ;
assign n15052 =  ( n98 ) & ( n13668 )  ;
assign n15053 =  ( n98 ) & ( n13670 )  ;
assign n15054 =  ( n98 ) & ( n13672 )  ;
assign n15055 =  ( n98 ) & ( n13674 )  ;
assign n15056 =  ( n98 ) & ( n13676 )  ;
assign n15057 =  ( n98 ) & ( n13678 )  ;
assign n15058 =  ( n98 ) & ( n13680 )  ;
assign n15059 =  ( n98 ) & ( n13682 )  ;
assign n15060 =  ( n98 ) & ( n13684 )  ;
assign n15061 =  ( n98 ) & ( n13686 )  ;
assign n15062 =  ( n98 ) & ( n13688 )  ;
assign n15063 =  ( n98 ) & ( n13690 )  ;
assign n15064 =  ( n98 ) & ( n13692 )  ;
assign n15065 =  ( n98 ) & ( n13694 )  ;
assign n15066 =  ( n99 ) & ( n13664 )  ;
assign n15067 =  ( n99 ) & ( n13666 )  ;
assign n15068 =  ( n99 ) & ( n13668 )  ;
assign n15069 =  ( n99 ) & ( n13670 )  ;
assign n15070 =  ( n99 ) & ( n13672 )  ;
assign n15071 =  ( n99 ) & ( n13674 )  ;
assign n15072 =  ( n99 ) & ( n13676 )  ;
assign n15073 =  ( n99 ) & ( n13678 )  ;
assign n15074 =  ( n99 ) & ( n13680 )  ;
assign n15075 =  ( n99 ) & ( n13682 )  ;
assign n15076 =  ( n99 ) & ( n13684 )  ;
assign n15077 =  ( n99 ) & ( n13686 )  ;
assign n15078 =  ( n99 ) & ( n13688 )  ;
assign n15079 =  ( n99 ) & ( n13690 )  ;
assign n15080 =  ( n99 ) & ( n13692 )  ;
assign n15081 =  ( n99 ) & ( n13694 )  ;
assign n15082 =  ( n100 ) & ( n13664 )  ;
assign n15083 =  ( n100 ) & ( n13666 )  ;
assign n15084 =  ( n100 ) & ( n13668 )  ;
assign n15085 =  ( n100 ) & ( n13670 )  ;
assign n15086 =  ( n100 ) & ( n13672 )  ;
assign n15087 =  ( n100 ) & ( n13674 )  ;
assign n15088 =  ( n100 ) & ( n13676 )  ;
assign n15089 =  ( n100 ) & ( n13678 )  ;
assign n15090 =  ( n100 ) & ( n13680 )  ;
assign n15091 =  ( n100 ) & ( n13682 )  ;
assign n15092 =  ( n100 ) & ( n13684 )  ;
assign n15093 =  ( n100 ) & ( n13686 )  ;
assign n15094 =  ( n100 ) & ( n13688 )  ;
assign n15095 =  ( n100 ) & ( n13690 )  ;
assign n15096 =  ( n100 ) & ( n13692 )  ;
assign n15097 =  ( n100 ) & ( n13694 )  ;
assign n15098 =  ( n101 ) & ( n13664 )  ;
assign n15099 =  ( n101 ) & ( n13666 )  ;
assign n15100 =  ( n101 ) & ( n13668 )  ;
assign n15101 =  ( n101 ) & ( n13670 )  ;
assign n15102 =  ( n101 ) & ( n13672 )  ;
assign n15103 =  ( n101 ) & ( n13674 )  ;
assign n15104 =  ( n101 ) & ( n13676 )  ;
assign n15105 =  ( n101 ) & ( n13678 )  ;
assign n15106 =  ( n101 ) & ( n13680 )  ;
assign n15107 =  ( n101 ) & ( n13682 )  ;
assign n15108 =  ( n101 ) & ( n13684 )  ;
assign n15109 =  ( n101 ) & ( n13686 )  ;
assign n15110 =  ( n101 ) & ( n13688 )  ;
assign n15111 =  ( n101 ) & ( n13690 )  ;
assign n15112 =  ( n101 ) & ( n13692 )  ;
assign n15113 =  ( n101 ) & ( n13694 )  ;
assign n15114 =  ( n102 ) & ( n13664 )  ;
assign n15115 =  ( n102 ) & ( n13666 )  ;
assign n15116 =  ( n102 ) & ( n13668 )  ;
assign n15117 =  ( n102 ) & ( n13670 )  ;
assign n15118 =  ( n102 ) & ( n13672 )  ;
assign n15119 =  ( n102 ) & ( n13674 )  ;
assign n15120 =  ( n102 ) & ( n13676 )  ;
assign n15121 =  ( n102 ) & ( n13678 )  ;
assign n15122 =  ( n102 ) & ( n13680 )  ;
assign n15123 =  ( n102 ) & ( n13682 )  ;
assign n15124 =  ( n102 ) & ( n13684 )  ;
assign n15125 =  ( n102 ) & ( n13686 )  ;
assign n15126 =  ( n102 ) & ( n13688 )  ;
assign n15127 =  ( n102 ) & ( n13690 )  ;
assign n15128 =  ( n102 ) & ( n13692 )  ;
assign n15129 =  ( n102 ) & ( n13694 )  ;
assign n15130 =  ( n103 ) & ( n13664 )  ;
assign n15131 =  ( n103 ) & ( n13666 )  ;
assign n15132 =  ( n103 ) & ( n13668 )  ;
assign n15133 =  ( n103 ) & ( n13670 )  ;
assign n15134 =  ( n103 ) & ( n13672 )  ;
assign n15135 =  ( n103 ) & ( n13674 )  ;
assign n15136 =  ( n103 ) & ( n13676 )  ;
assign n15137 =  ( n103 ) & ( n13678 )  ;
assign n15138 =  ( n103 ) & ( n13680 )  ;
assign n15139 =  ( n103 ) & ( n13682 )  ;
assign n15140 =  ( n103 ) & ( n13684 )  ;
assign n15141 =  ( n103 ) & ( n13686 )  ;
assign n15142 =  ( n103 ) & ( n13688 )  ;
assign n15143 =  ( n103 ) & ( n13690 )  ;
assign n15144 =  ( n103 ) & ( n13692 )  ;
assign n15145 =  ( n103 ) & ( n13694 )  ;
assign n15146 =  ( n104 ) & ( n13664 )  ;
assign n15147 =  ( n104 ) & ( n13666 )  ;
assign n15148 =  ( n104 ) & ( n13668 )  ;
assign n15149 =  ( n104 ) & ( n13670 )  ;
assign n15150 =  ( n104 ) & ( n13672 )  ;
assign n15151 =  ( n104 ) & ( n13674 )  ;
assign n15152 =  ( n104 ) & ( n13676 )  ;
assign n15153 =  ( n104 ) & ( n13678 )  ;
assign n15154 =  ( n104 ) & ( n13680 )  ;
assign n15155 =  ( n104 ) & ( n13682 )  ;
assign n15156 =  ( n104 ) & ( n13684 )  ;
assign n15157 =  ( n104 ) & ( n13686 )  ;
assign n15158 =  ( n104 ) & ( n13688 )  ;
assign n15159 =  ( n104 ) & ( n13690 )  ;
assign n15160 =  ( n104 ) & ( n13692 )  ;
assign n15161 =  ( n104 ) & ( n13694 )  ;
assign n15162 =  ( n105 ) & ( n13664 )  ;
assign n15163 =  ( n105 ) & ( n13666 )  ;
assign n15164 =  ( n105 ) & ( n13668 )  ;
assign n15165 =  ( n105 ) & ( n13670 )  ;
assign n15166 =  ( n105 ) & ( n13672 )  ;
assign n15167 =  ( n105 ) & ( n13674 )  ;
assign n15168 =  ( n105 ) & ( n13676 )  ;
assign n15169 =  ( n105 ) & ( n13678 )  ;
assign n15170 =  ( n105 ) & ( n13680 )  ;
assign n15171 =  ( n105 ) & ( n13682 )  ;
assign n15172 =  ( n105 ) & ( n13684 )  ;
assign n15173 =  ( n105 ) & ( n13686 )  ;
assign n15174 =  ( n105 ) & ( n13688 )  ;
assign n15175 =  ( n105 ) & ( n13690 )  ;
assign n15176 =  ( n105 ) & ( n13692 )  ;
assign n15177 =  ( n105 ) & ( n13694 )  ;
assign n15178 =  ( n106 ) & ( n13664 )  ;
assign n15179 =  ( n106 ) & ( n13666 )  ;
assign n15180 =  ( n106 ) & ( n13668 )  ;
assign n15181 =  ( n106 ) & ( n13670 )  ;
assign n15182 =  ( n106 ) & ( n13672 )  ;
assign n15183 =  ( n106 ) & ( n13674 )  ;
assign n15184 =  ( n106 ) & ( n13676 )  ;
assign n15185 =  ( n106 ) & ( n13678 )  ;
assign n15186 =  ( n106 ) & ( n13680 )  ;
assign n15187 =  ( n106 ) & ( n13682 )  ;
assign n15188 =  ( n106 ) & ( n13684 )  ;
assign n15189 =  ( n106 ) & ( n13686 )  ;
assign n15190 =  ( n106 ) & ( n13688 )  ;
assign n15191 =  ( n106 ) & ( n13690 )  ;
assign n15192 =  ( n106 ) & ( n13692 )  ;
assign n15193 =  ( n106 ) & ( n13694 )  ;
assign n15194 =  ( n107 ) & ( n13664 )  ;
assign n15195 =  ( n107 ) & ( n13666 )  ;
assign n15196 =  ( n107 ) & ( n13668 )  ;
assign n15197 =  ( n107 ) & ( n13670 )  ;
assign n15198 =  ( n107 ) & ( n13672 )  ;
assign n15199 =  ( n107 ) & ( n13674 )  ;
assign n15200 =  ( n107 ) & ( n13676 )  ;
assign n15201 =  ( n107 ) & ( n13678 )  ;
assign n15202 =  ( n107 ) & ( n13680 )  ;
assign n15203 =  ( n107 ) & ( n13682 )  ;
assign n15204 =  ( n107 ) & ( n13684 )  ;
assign n15205 =  ( n107 ) & ( n13686 )  ;
assign n15206 =  ( n107 ) & ( n13688 )  ;
assign n15207 =  ( n107 ) & ( n13690 )  ;
assign n15208 =  ( n107 ) & ( n13692 )  ;
assign n15209 =  ( n107 ) & ( n13694 )  ;
assign n15210 =  ( n108 ) & ( n13664 )  ;
assign n15211 =  ( n108 ) & ( n13666 )  ;
assign n15212 =  ( n108 ) & ( n13668 )  ;
assign n15213 =  ( n108 ) & ( n13670 )  ;
assign n15214 =  ( n108 ) & ( n13672 )  ;
assign n15215 =  ( n108 ) & ( n13674 )  ;
assign n15216 =  ( n108 ) & ( n13676 )  ;
assign n15217 =  ( n108 ) & ( n13678 )  ;
assign n15218 =  ( n108 ) & ( n13680 )  ;
assign n15219 =  ( n108 ) & ( n13682 )  ;
assign n15220 =  ( n108 ) & ( n13684 )  ;
assign n15221 =  ( n108 ) & ( n13686 )  ;
assign n15222 =  ( n108 ) & ( n13688 )  ;
assign n15223 =  ( n108 ) & ( n13690 )  ;
assign n15224 =  ( n108 ) & ( n13692 )  ;
assign n15225 =  ( n108 ) & ( n13694 )  ;
assign n15226 =  ( n15225 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n15227 =  ( n15224 ) ? ( VREG_0_1 ) : ( n15226 ) ;
assign n15228 =  ( n15223 ) ? ( VREG_0_2 ) : ( n15227 ) ;
assign n15229 =  ( n15222 ) ? ( VREG_0_3 ) : ( n15228 ) ;
assign n15230 =  ( n15221 ) ? ( VREG_0_4 ) : ( n15229 ) ;
assign n15231 =  ( n15220 ) ? ( VREG_0_5 ) : ( n15230 ) ;
assign n15232 =  ( n15219 ) ? ( VREG_0_6 ) : ( n15231 ) ;
assign n15233 =  ( n15218 ) ? ( VREG_0_7 ) : ( n15232 ) ;
assign n15234 =  ( n15217 ) ? ( VREG_0_8 ) : ( n15233 ) ;
assign n15235 =  ( n15216 ) ? ( VREG_0_9 ) : ( n15234 ) ;
assign n15236 =  ( n15215 ) ? ( VREG_0_10 ) : ( n15235 ) ;
assign n15237 =  ( n15214 ) ? ( VREG_0_11 ) : ( n15236 ) ;
assign n15238 =  ( n15213 ) ? ( VREG_0_12 ) : ( n15237 ) ;
assign n15239 =  ( n15212 ) ? ( VREG_0_13 ) : ( n15238 ) ;
assign n15240 =  ( n15211 ) ? ( VREG_0_14 ) : ( n15239 ) ;
assign n15241 =  ( n15210 ) ? ( VREG_0_15 ) : ( n15240 ) ;
assign n15242 =  ( n15209 ) ? ( VREG_1_0 ) : ( n15241 ) ;
assign n15243 =  ( n15208 ) ? ( VREG_1_1 ) : ( n15242 ) ;
assign n15244 =  ( n15207 ) ? ( VREG_1_2 ) : ( n15243 ) ;
assign n15245 =  ( n15206 ) ? ( VREG_1_3 ) : ( n15244 ) ;
assign n15246 =  ( n15205 ) ? ( VREG_1_4 ) : ( n15245 ) ;
assign n15247 =  ( n15204 ) ? ( VREG_1_5 ) : ( n15246 ) ;
assign n15248 =  ( n15203 ) ? ( VREG_1_6 ) : ( n15247 ) ;
assign n15249 =  ( n15202 ) ? ( VREG_1_7 ) : ( n15248 ) ;
assign n15250 =  ( n15201 ) ? ( VREG_1_8 ) : ( n15249 ) ;
assign n15251 =  ( n15200 ) ? ( VREG_1_9 ) : ( n15250 ) ;
assign n15252 =  ( n15199 ) ? ( VREG_1_10 ) : ( n15251 ) ;
assign n15253 =  ( n15198 ) ? ( VREG_1_11 ) : ( n15252 ) ;
assign n15254 =  ( n15197 ) ? ( VREG_1_12 ) : ( n15253 ) ;
assign n15255 =  ( n15196 ) ? ( VREG_1_13 ) : ( n15254 ) ;
assign n15256 =  ( n15195 ) ? ( VREG_1_14 ) : ( n15255 ) ;
assign n15257 =  ( n15194 ) ? ( VREG_1_15 ) : ( n15256 ) ;
assign n15258 =  ( n15193 ) ? ( VREG_2_0 ) : ( n15257 ) ;
assign n15259 =  ( n15192 ) ? ( VREG_2_1 ) : ( n15258 ) ;
assign n15260 =  ( n15191 ) ? ( VREG_2_2 ) : ( n15259 ) ;
assign n15261 =  ( n15190 ) ? ( VREG_2_3 ) : ( n15260 ) ;
assign n15262 =  ( n15189 ) ? ( VREG_2_4 ) : ( n15261 ) ;
assign n15263 =  ( n15188 ) ? ( VREG_2_5 ) : ( n15262 ) ;
assign n15264 =  ( n15187 ) ? ( VREG_2_6 ) : ( n15263 ) ;
assign n15265 =  ( n15186 ) ? ( VREG_2_7 ) : ( n15264 ) ;
assign n15266 =  ( n15185 ) ? ( VREG_2_8 ) : ( n15265 ) ;
assign n15267 =  ( n15184 ) ? ( VREG_2_9 ) : ( n15266 ) ;
assign n15268 =  ( n15183 ) ? ( VREG_2_10 ) : ( n15267 ) ;
assign n15269 =  ( n15182 ) ? ( VREG_2_11 ) : ( n15268 ) ;
assign n15270 =  ( n15181 ) ? ( VREG_2_12 ) : ( n15269 ) ;
assign n15271 =  ( n15180 ) ? ( VREG_2_13 ) : ( n15270 ) ;
assign n15272 =  ( n15179 ) ? ( VREG_2_14 ) : ( n15271 ) ;
assign n15273 =  ( n15178 ) ? ( VREG_2_15 ) : ( n15272 ) ;
assign n15274 =  ( n15177 ) ? ( VREG_3_0 ) : ( n15273 ) ;
assign n15275 =  ( n15176 ) ? ( VREG_3_1 ) : ( n15274 ) ;
assign n15276 =  ( n15175 ) ? ( VREG_3_2 ) : ( n15275 ) ;
assign n15277 =  ( n15174 ) ? ( VREG_3_3 ) : ( n15276 ) ;
assign n15278 =  ( n15173 ) ? ( VREG_3_4 ) : ( n15277 ) ;
assign n15279 =  ( n15172 ) ? ( VREG_3_5 ) : ( n15278 ) ;
assign n15280 =  ( n15171 ) ? ( VREG_3_6 ) : ( n15279 ) ;
assign n15281 =  ( n15170 ) ? ( VREG_3_7 ) : ( n15280 ) ;
assign n15282 =  ( n15169 ) ? ( VREG_3_8 ) : ( n15281 ) ;
assign n15283 =  ( n15168 ) ? ( VREG_3_9 ) : ( n15282 ) ;
assign n15284 =  ( n15167 ) ? ( VREG_3_10 ) : ( n15283 ) ;
assign n15285 =  ( n15166 ) ? ( VREG_3_11 ) : ( n15284 ) ;
assign n15286 =  ( n15165 ) ? ( VREG_3_12 ) : ( n15285 ) ;
assign n15287 =  ( n15164 ) ? ( VREG_3_13 ) : ( n15286 ) ;
assign n15288 =  ( n15163 ) ? ( VREG_3_14 ) : ( n15287 ) ;
assign n15289 =  ( n15162 ) ? ( VREG_3_15 ) : ( n15288 ) ;
assign n15290 =  ( n15161 ) ? ( VREG_4_0 ) : ( n15289 ) ;
assign n15291 =  ( n15160 ) ? ( VREG_4_1 ) : ( n15290 ) ;
assign n15292 =  ( n15159 ) ? ( VREG_4_2 ) : ( n15291 ) ;
assign n15293 =  ( n15158 ) ? ( VREG_4_3 ) : ( n15292 ) ;
assign n15294 =  ( n15157 ) ? ( VREG_4_4 ) : ( n15293 ) ;
assign n15295 =  ( n15156 ) ? ( VREG_4_5 ) : ( n15294 ) ;
assign n15296 =  ( n15155 ) ? ( VREG_4_6 ) : ( n15295 ) ;
assign n15297 =  ( n15154 ) ? ( VREG_4_7 ) : ( n15296 ) ;
assign n15298 =  ( n15153 ) ? ( VREG_4_8 ) : ( n15297 ) ;
assign n15299 =  ( n15152 ) ? ( VREG_4_9 ) : ( n15298 ) ;
assign n15300 =  ( n15151 ) ? ( VREG_4_10 ) : ( n15299 ) ;
assign n15301 =  ( n15150 ) ? ( VREG_4_11 ) : ( n15300 ) ;
assign n15302 =  ( n15149 ) ? ( VREG_4_12 ) : ( n15301 ) ;
assign n15303 =  ( n15148 ) ? ( VREG_4_13 ) : ( n15302 ) ;
assign n15304 =  ( n15147 ) ? ( VREG_4_14 ) : ( n15303 ) ;
assign n15305 =  ( n15146 ) ? ( VREG_4_15 ) : ( n15304 ) ;
assign n15306 =  ( n15145 ) ? ( VREG_5_0 ) : ( n15305 ) ;
assign n15307 =  ( n15144 ) ? ( VREG_5_1 ) : ( n15306 ) ;
assign n15308 =  ( n15143 ) ? ( VREG_5_2 ) : ( n15307 ) ;
assign n15309 =  ( n15142 ) ? ( VREG_5_3 ) : ( n15308 ) ;
assign n15310 =  ( n15141 ) ? ( VREG_5_4 ) : ( n15309 ) ;
assign n15311 =  ( n15140 ) ? ( VREG_5_5 ) : ( n15310 ) ;
assign n15312 =  ( n15139 ) ? ( VREG_5_6 ) : ( n15311 ) ;
assign n15313 =  ( n15138 ) ? ( VREG_5_7 ) : ( n15312 ) ;
assign n15314 =  ( n15137 ) ? ( VREG_5_8 ) : ( n15313 ) ;
assign n15315 =  ( n15136 ) ? ( VREG_5_9 ) : ( n15314 ) ;
assign n15316 =  ( n15135 ) ? ( VREG_5_10 ) : ( n15315 ) ;
assign n15317 =  ( n15134 ) ? ( VREG_5_11 ) : ( n15316 ) ;
assign n15318 =  ( n15133 ) ? ( VREG_5_12 ) : ( n15317 ) ;
assign n15319 =  ( n15132 ) ? ( VREG_5_13 ) : ( n15318 ) ;
assign n15320 =  ( n15131 ) ? ( VREG_5_14 ) : ( n15319 ) ;
assign n15321 =  ( n15130 ) ? ( VREG_5_15 ) : ( n15320 ) ;
assign n15322 =  ( n15129 ) ? ( VREG_6_0 ) : ( n15321 ) ;
assign n15323 =  ( n15128 ) ? ( VREG_6_1 ) : ( n15322 ) ;
assign n15324 =  ( n15127 ) ? ( VREG_6_2 ) : ( n15323 ) ;
assign n15325 =  ( n15126 ) ? ( VREG_6_3 ) : ( n15324 ) ;
assign n15326 =  ( n15125 ) ? ( VREG_6_4 ) : ( n15325 ) ;
assign n15327 =  ( n15124 ) ? ( VREG_6_5 ) : ( n15326 ) ;
assign n15328 =  ( n15123 ) ? ( VREG_6_6 ) : ( n15327 ) ;
assign n15329 =  ( n15122 ) ? ( VREG_6_7 ) : ( n15328 ) ;
assign n15330 =  ( n15121 ) ? ( VREG_6_8 ) : ( n15329 ) ;
assign n15331 =  ( n15120 ) ? ( VREG_6_9 ) : ( n15330 ) ;
assign n15332 =  ( n15119 ) ? ( VREG_6_10 ) : ( n15331 ) ;
assign n15333 =  ( n15118 ) ? ( VREG_6_11 ) : ( n15332 ) ;
assign n15334 =  ( n15117 ) ? ( VREG_6_12 ) : ( n15333 ) ;
assign n15335 =  ( n15116 ) ? ( VREG_6_13 ) : ( n15334 ) ;
assign n15336 =  ( n15115 ) ? ( VREG_6_14 ) : ( n15335 ) ;
assign n15337 =  ( n15114 ) ? ( VREG_6_15 ) : ( n15336 ) ;
assign n15338 =  ( n15113 ) ? ( VREG_7_0 ) : ( n15337 ) ;
assign n15339 =  ( n15112 ) ? ( VREG_7_1 ) : ( n15338 ) ;
assign n15340 =  ( n15111 ) ? ( VREG_7_2 ) : ( n15339 ) ;
assign n15341 =  ( n15110 ) ? ( VREG_7_3 ) : ( n15340 ) ;
assign n15342 =  ( n15109 ) ? ( VREG_7_4 ) : ( n15341 ) ;
assign n15343 =  ( n15108 ) ? ( VREG_7_5 ) : ( n15342 ) ;
assign n15344 =  ( n15107 ) ? ( VREG_7_6 ) : ( n15343 ) ;
assign n15345 =  ( n15106 ) ? ( VREG_7_7 ) : ( n15344 ) ;
assign n15346 =  ( n15105 ) ? ( VREG_7_8 ) : ( n15345 ) ;
assign n15347 =  ( n15104 ) ? ( VREG_7_9 ) : ( n15346 ) ;
assign n15348 =  ( n15103 ) ? ( VREG_7_10 ) : ( n15347 ) ;
assign n15349 =  ( n15102 ) ? ( VREG_7_11 ) : ( n15348 ) ;
assign n15350 =  ( n15101 ) ? ( VREG_7_12 ) : ( n15349 ) ;
assign n15351 =  ( n15100 ) ? ( VREG_7_13 ) : ( n15350 ) ;
assign n15352 =  ( n15099 ) ? ( VREG_7_14 ) : ( n15351 ) ;
assign n15353 =  ( n15098 ) ? ( VREG_7_15 ) : ( n15352 ) ;
assign n15354 =  ( n15097 ) ? ( VREG_8_0 ) : ( n15353 ) ;
assign n15355 =  ( n15096 ) ? ( VREG_8_1 ) : ( n15354 ) ;
assign n15356 =  ( n15095 ) ? ( VREG_8_2 ) : ( n15355 ) ;
assign n15357 =  ( n15094 ) ? ( VREG_8_3 ) : ( n15356 ) ;
assign n15358 =  ( n15093 ) ? ( VREG_8_4 ) : ( n15357 ) ;
assign n15359 =  ( n15092 ) ? ( VREG_8_5 ) : ( n15358 ) ;
assign n15360 =  ( n15091 ) ? ( VREG_8_6 ) : ( n15359 ) ;
assign n15361 =  ( n15090 ) ? ( VREG_8_7 ) : ( n15360 ) ;
assign n15362 =  ( n15089 ) ? ( VREG_8_8 ) : ( n15361 ) ;
assign n15363 =  ( n15088 ) ? ( VREG_8_9 ) : ( n15362 ) ;
assign n15364 =  ( n15087 ) ? ( VREG_8_10 ) : ( n15363 ) ;
assign n15365 =  ( n15086 ) ? ( VREG_8_11 ) : ( n15364 ) ;
assign n15366 =  ( n15085 ) ? ( VREG_8_12 ) : ( n15365 ) ;
assign n15367 =  ( n15084 ) ? ( VREG_8_13 ) : ( n15366 ) ;
assign n15368 =  ( n15083 ) ? ( VREG_8_14 ) : ( n15367 ) ;
assign n15369 =  ( n15082 ) ? ( VREG_8_15 ) : ( n15368 ) ;
assign n15370 =  ( n15081 ) ? ( VREG_9_0 ) : ( n15369 ) ;
assign n15371 =  ( n15080 ) ? ( VREG_9_1 ) : ( n15370 ) ;
assign n15372 =  ( n15079 ) ? ( VREG_9_2 ) : ( n15371 ) ;
assign n15373 =  ( n15078 ) ? ( VREG_9_3 ) : ( n15372 ) ;
assign n15374 =  ( n15077 ) ? ( VREG_9_4 ) : ( n15373 ) ;
assign n15375 =  ( n15076 ) ? ( VREG_9_5 ) : ( n15374 ) ;
assign n15376 =  ( n15075 ) ? ( VREG_9_6 ) : ( n15375 ) ;
assign n15377 =  ( n15074 ) ? ( VREG_9_7 ) : ( n15376 ) ;
assign n15378 =  ( n15073 ) ? ( VREG_9_8 ) : ( n15377 ) ;
assign n15379 =  ( n15072 ) ? ( VREG_9_9 ) : ( n15378 ) ;
assign n15380 =  ( n15071 ) ? ( VREG_9_10 ) : ( n15379 ) ;
assign n15381 =  ( n15070 ) ? ( VREG_9_11 ) : ( n15380 ) ;
assign n15382 =  ( n15069 ) ? ( VREG_9_12 ) : ( n15381 ) ;
assign n15383 =  ( n15068 ) ? ( VREG_9_13 ) : ( n15382 ) ;
assign n15384 =  ( n15067 ) ? ( VREG_9_14 ) : ( n15383 ) ;
assign n15385 =  ( n15066 ) ? ( VREG_9_15 ) : ( n15384 ) ;
assign n15386 =  ( n15065 ) ? ( VREG_10_0 ) : ( n15385 ) ;
assign n15387 =  ( n15064 ) ? ( VREG_10_1 ) : ( n15386 ) ;
assign n15388 =  ( n15063 ) ? ( VREG_10_2 ) : ( n15387 ) ;
assign n15389 =  ( n15062 ) ? ( VREG_10_3 ) : ( n15388 ) ;
assign n15390 =  ( n15061 ) ? ( VREG_10_4 ) : ( n15389 ) ;
assign n15391 =  ( n15060 ) ? ( VREG_10_5 ) : ( n15390 ) ;
assign n15392 =  ( n15059 ) ? ( VREG_10_6 ) : ( n15391 ) ;
assign n15393 =  ( n15058 ) ? ( VREG_10_7 ) : ( n15392 ) ;
assign n15394 =  ( n15057 ) ? ( VREG_10_8 ) : ( n15393 ) ;
assign n15395 =  ( n15056 ) ? ( VREG_10_9 ) : ( n15394 ) ;
assign n15396 =  ( n15055 ) ? ( VREG_10_10 ) : ( n15395 ) ;
assign n15397 =  ( n15054 ) ? ( VREG_10_11 ) : ( n15396 ) ;
assign n15398 =  ( n15053 ) ? ( VREG_10_12 ) : ( n15397 ) ;
assign n15399 =  ( n15052 ) ? ( VREG_10_13 ) : ( n15398 ) ;
assign n15400 =  ( n15051 ) ? ( VREG_10_14 ) : ( n15399 ) ;
assign n15401 =  ( n15050 ) ? ( VREG_10_15 ) : ( n15400 ) ;
assign n15402 =  ( n15049 ) ? ( VREG_11_0 ) : ( n15401 ) ;
assign n15403 =  ( n15048 ) ? ( VREG_11_1 ) : ( n15402 ) ;
assign n15404 =  ( n15047 ) ? ( VREG_11_2 ) : ( n15403 ) ;
assign n15405 =  ( n15046 ) ? ( VREG_11_3 ) : ( n15404 ) ;
assign n15406 =  ( n15045 ) ? ( VREG_11_4 ) : ( n15405 ) ;
assign n15407 =  ( n15044 ) ? ( VREG_11_5 ) : ( n15406 ) ;
assign n15408 =  ( n15043 ) ? ( VREG_11_6 ) : ( n15407 ) ;
assign n15409 =  ( n15042 ) ? ( VREG_11_7 ) : ( n15408 ) ;
assign n15410 =  ( n15041 ) ? ( VREG_11_8 ) : ( n15409 ) ;
assign n15411 =  ( n15040 ) ? ( VREG_11_9 ) : ( n15410 ) ;
assign n15412 =  ( n15039 ) ? ( VREG_11_10 ) : ( n15411 ) ;
assign n15413 =  ( n15038 ) ? ( VREG_11_11 ) : ( n15412 ) ;
assign n15414 =  ( n15037 ) ? ( VREG_11_12 ) : ( n15413 ) ;
assign n15415 =  ( n15036 ) ? ( VREG_11_13 ) : ( n15414 ) ;
assign n15416 =  ( n15035 ) ? ( VREG_11_14 ) : ( n15415 ) ;
assign n15417 =  ( n15034 ) ? ( VREG_11_15 ) : ( n15416 ) ;
assign n15418 =  ( n15033 ) ? ( VREG_12_0 ) : ( n15417 ) ;
assign n15419 =  ( n15032 ) ? ( VREG_12_1 ) : ( n15418 ) ;
assign n15420 =  ( n15031 ) ? ( VREG_12_2 ) : ( n15419 ) ;
assign n15421 =  ( n15030 ) ? ( VREG_12_3 ) : ( n15420 ) ;
assign n15422 =  ( n15029 ) ? ( VREG_12_4 ) : ( n15421 ) ;
assign n15423 =  ( n15028 ) ? ( VREG_12_5 ) : ( n15422 ) ;
assign n15424 =  ( n15027 ) ? ( VREG_12_6 ) : ( n15423 ) ;
assign n15425 =  ( n15026 ) ? ( VREG_12_7 ) : ( n15424 ) ;
assign n15426 =  ( n15025 ) ? ( VREG_12_8 ) : ( n15425 ) ;
assign n15427 =  ( n15024 ) ? ( VREG_12_9 ) : ( n15426 ) ;
assign n15428 =  ( n15023 ) ? ( VREG_12_10 ) : ( n15427 ) ;
assign n15429 =  ( n15022 ) ? ( VREG_12_11 ) : ( n15428 ) ;
assign n15430 =  ( n15021 ) ? ( VREG_12_12 ) : ( n15429 ) ;
assign n15431 =  ( n15020 ) ? ( VREG_12_13 ) : ( n15430 ) ;
assign n15432 =  ( n15019 ) ? ( VREG_12_14 ) : ( n15431 ) ;
assign n15433 =  ( n15018 ) ? ( VREG_12_15 ) : ( n15432 ) ;
assign n15434 =  ( n15017 ) ? ( VREG_13_0 ) : ( n15433 ) ;
assign n15435 =  ( n15016 ) ? ( VREG_13_1 ) : ( n15434 ) ;
assign n15436 =  ( n15015 ) ? ( VREG_13_2 ) : ( n15435 ) ;
assign n15437 =  ( n15014 ) ? ( VREG_13_3 ) : ( n15436 ) ;
assign n15438 =  ( n15013 ) ? ( VREG_13_4 ) : ( n15437 ) ;
assign n15439 =  ( n15012 ) ? ( VREG_13_5 ) : ( n15438 ) ;
assign n15440 =  ( n15011 ) ? ( VREG_13_6 ) : ( n15439 ) ;
assign n15441 =  ( n15010 ) ? ( VREG_13_7 ) : ( n15440 ) ;
assign n15442 =  ( n15009 ) ? ( VREG_13_8 ) : ( n15441 ) ;
assign n15443 =  ( n15008 ) ? ( VREG_13_9 ) : ( n15442 ) ;
assign n15444 =  ( n15007 ) ? ( VREG_13_10 ) : ( n15443 ) ;
assign n15445 =  ( n15006 ) ? ( VREG_13_11 ) : ( n15444 ) ;
assign n15446 =  ( n15005 ) ? ( VREG_13_12 ) : ( n15445 ) ;
assign n15447 =  ( n15004 ) ? ( VREG_13_13 ) : ( n15446 ) ;
assign n15448 =  ( n15003 ) ? ( VREG_13_14 ) : ( n15447 ) ;
assign n15449 =  ( n15002 ) ? ( VREG_13_15 ) : ( n15448 ) ;
assign n15450 =  ( n15001 ) ? ( VREG_14_0 ) : ( n15449 ) ;
assign n15451 =  ( n15000 ) ? ( VREG_14_1 ) : ( n15450 ) ;
assign n15452 =  ( n14999 ) ? ( VREG_14_2 ) : ( n15451 ) ;
assign n15453 =  ( n14998 ) ? ( VREG_14_3 ) : ( n15452 ) ;
assign n15454 =  ( n14997 ) ? ( VREG_14_4 ) : ( n15453 ) ;
assign n15455 =  ( n14996 ) ? ( VREG_14_5 ) : ( n15454 ) ;
assign n15456 =  ( n14995 ) ? ( VREG_14_6 ) : ( n15455 ) ;
assign n15457 =  ( n14994 ) ? ( VREG_14_7 ) : ( n15456 ) ;
assign n15458 =  ( n14993 ) ? ( VREG_14_8 ) : ( n15457 ) ;
assign n15459 =  ( n14992 ) ? ( VREG_14_9 ) : ( n15458 ) ;
assign n15460 =  ( n14991 ) ? ( VREG_14_10 ) : ( n15459 ) ;
assign n15461 =  ( n14990 ) ? ( VREG_14_11 ) : ( n15460 ) ;
assign n15462 =  ( n14989 ) ? ( VREG_14_12 ) : ( n15461 ) ;
assign n15463 =  ( n14988 ) ? ( VREG_14_13 ) : ( n15462 ) ;
assign n15464 =  ( n14987 ) ? ( VREG_14_14 ) : ( n15463 ) ;
assign n15465 =  ( n14986 ) ? ( VREG_14_15 ) : ( n15464 ) ;
assign n15466 =  ( n14985 ) ? ( VREG_15_0 ) : ( n15465 ) ;
assign n15467 =  ( n14984 ) ? ( VREG_15_1 ) : ( n15466 ) ;
assign n15468 =  ( n14983 ) ? ( VREG_15_2 ) : ( n15467 ) ;
assign n15469 =  ( n14982 ) ? ( VREG_15_3 ) : ( n15468 ) ;
assign n15470 =  ( n14981 ) ? ( VREG_15_4 ) : ( n15469 ) ;
assign n15471 =  ( n14980 ) ? ( VREG_15_5 ) : ( n15470 ) ;
assign n15472 =  ( n14979 ) ? ( VREG_15_6 ) : ( n15471 ) ;
assign n15473 =  ( n14978 ) ? ( VREG_15_7 ) : ( n15472 ) ;
assign n15474 =  ( n14977 ) ? ( VREG_15_8 ) : ( n15473 ) ;
assign n15475 =  ( n14976 ) ? ( VREG_15_9 ) : ( n15474 ) ;
assign n15476 =  ( n14975 ) ? ( VREG_15_10 ) : ( n15475 ) ;
assign n15477 =  ( n14974 ) ? ( VREG_15_11 ) : ( n15476 ) ;
assign n15478 =  ( n14973 ) ? ( VREG_15_12 ) : ( n15477 ) ;
assign n15479 =  ( n14972 ) ? ( VREG_15_13 ) : ( n15478 ) ;
assign n15480 =  ( n14971 ) ? ( VREG_15_14 ) : ( n15479 ) ;
assign n15481 =  ( n14970 ) ? ( VREG_15_15 ) : ( n15480 ) ;
assign n15482 =  ( n14969 ) ? ( VREG_16_0 ) : ( n15481 ) ;
assign n15483 =  ( n14968 ) ? ( VREG_16_1 ) : ( n15482 ) ;
assign n15484 =  ( n14967 ) ? ( VREG_16_2 ) : ( n15483 ) ;
assign n15485 =  ( n14966 ) ? ( VREG_16_3 ) : ( n15484 ) ;
assign n15486 =  ( n14965 ) ? ( VREG_16_4 ) : ( n15485 ) ;
assign n15487 =  ( n14964 ) ? ( VREG_16_5 ) : ( n15486 ) ;
assign n15488 =  ( n14963 ) ? ( VREG_16_6 ) : ( n15487 ) ;
assign n15489 =  ( n14962 ) ? ( VREG_16_7 ) : ( n15488 ) ;
assign n15490 =  ( n14961 ) ? ( VREG_16_8 ) : ( n15489 ) ;
assign n15491 =  ( n14960 ) ? ( VREG_16_9 ) : ( n15490 ) ;
assign n15492 =  ( n14959 ) ? ( VREG_16_10 ) : ( n15491 ) ;
assign n15493 =  ( n14958 ) ? ( VREG_16_11 ) : ( n15492 ) ;
assign n15494 =  ( n14957 ) ? ( VREG_16_12 ) : ( n15493 ) ;
assign n15495 =  ( n14956 ) ? ( VREG_16_13 ) : ( n15494 ) ;
assign n15496 =  ( n14955 ) ? ( VREG_16_14 ) : ( n15495 ) ;
assign n15497 =  ( n14954 ) ? ( VREG_16_15 ) : ( n15496 ) ;
assign n15498 =  ( n14953 ) ? ( VREG_17_0 ) : ( n15497 ) ;
assign n15499 =  ( n14952 ) ? ( VREG_17_1 ) : ( n15498 ) ;
assign n15500 =  ( n14951 ) ? ( VREG_17_2 ) : ( n15499 ) ;
assign n15501 =  ( n14950 ) ? ( VREG_17_3 ) : ( n15500 ) ;
assign n15502 =  ( n14949 ) ? ( VREG_17_4 ) : ( n15501 ) ;
assign n15503 =  ( n14948 ) ? ( VREG_17_5 ) : ( n15502 ) ;
assign n15504 =  ( n14947 ) ? ( VREG_17_6 ) : ( n15503 ) ;
assign n15505 =  ( n14946 ) ? ( VREG_17_7 ) : ( n15504 ) ;
assign n15506 =  ( n14945 ) ? ( VREG_17_8 ) : ( n15505 ) ;
assign n15507 =  ( n14944 ) ? ( VREG_17_9 ) : ( n15506 ) ;
assign n15508 =  ( n14943 ) ? ( VREG_17_10 ) : ( n15507 ) ;
assign n15509 =  ( n14942 ) ? ( VREG_17_11 ) : ( n15508 ) ;
assign n15510 =  ( n14941 ) ? ( VREG_17_12 ) : ( n15509 ) ;
assign n15511 =  ( n14940 ) ? ( VREG_17_13 ) : ( n15510 ) ;
assign n15512 =  ( n14939 ) ? ( VREG_17_14 ) : ( n15511 ) ;
assign n15513 =  ( n14938 ) ? ( VREG_17_15 ) : ( n15512 ) ;
assign n15514 =  ( n14937 ) ? ( VREG_18_0 ) : ( n15513 ) ;
assign n15515 =  ( n14936 ) ? ( VREG_18_1 ) : ( n15514 ) ;
assign n15516 =  ( n14935 ) ? ( VREG_18_2 ) : ( n15515 ) ;
assign n15517 =  ( n14934 ) ? ( VREG_18_3 ) : ( n15516 ) ;
assign n15518 =  ( n14933 ) ? ( VREG_18_4 ) : ( n15517 ) ;
assign n15519 =  ( n14932 ) ? ( VREG_18_5 ) : ( n15518 ) ;
assign n15520 =  ( n14931 ) ? ( VREG_18_6 ) : ( n15519 ) ;
assign n15521 =  ( n14930 ) ? ( VREG_18_7 ) : ( n15520 ) ;
assign n15522 =  ( n14929 ) ? ( VREG_18_8 ) : ( n15521 ) ;
assign n15523 =  ( n14928 ) ? ( VREG_18_9 ) : ( n15522 ) ;
assign n15524 =  ( n14927 ) ? ( VREG_18_10 ) : ( n15523 ) ;
assign n15525 =  ( n14926 ) ? ( VREG_18_11 ) : ( n15524 ) ;
assign n15526 =  ( n14925 ) ? ( VREG_18_12 ) : ( n15525 ) ;
assign n15527 =  ( n14924 ) ? ( VREG_18_13 ) : ( n15526 ) ;
assign n15528 =  ( n14923 ) ? ( VREG_18_14 ) : ( n15527 ) ;
assign n15529 =  ( n14922 ) ? ( VREG_18_15 ) : ( n15528 ) ;
assign n15530 =  ( n14921 ) ? ( VREG_19_0 ) : ( n15529 ) ;
assign n15531 =  ( n14920 ) ? ( VREG_19_1 ) : ( n15530 ) ;
assign n15532 =  ( n14919 ) ? ( VREG_19_2 ) : ( n15531 ) ;
assign n15533 =  ( n14918 ) ? ( VREG_19_3 ) : ( n15532 ) ;
assign n15534 =  ( n14917 ) ? ( VREG_19_4 ) : ( n15533 ) ;
assign n15535 =  ( n14916 ) ? ( VREG_19_5 ) : ( n15534 ) ;
assign n15536 =  ( n14915 ) ? ( VREG_19_6 ) : ( n15535 ) ;
assign n15537 =  ( n14914 ) ? ( VREG_19_7 ) : ( n15536 ) ;
assign n15538 =  ( n14913 ) ? ( VREG_19_8 ) : ( n15537 ) ;
assign n15539 =  ( n14912 ) ? ( VREG_19_9 ) : ( n15538 ) ;
assign n15540 =  ( n14911 ) ? ( VREG_19_10 ) : ( n15539 ) ;
assign n15541 =  ( n14910 ) ? ( VREG_19_11 ) : ( n15540 ) ;
assign n15542 =  ( n14909 ) ? ( VREG_19_12 ) : ( n15541 ) ;
assign n15543 =  ( n14908 ) ? ( VREG_19_13 ) : ( n15542 ) ;
assign n15544 =  ( n14907 ) ? ( VREG_19_14 ) : ( n15543 ) ;
assign n15545 =  ( n14906 ) ? ( VREG_19_15 ) : ( n15544 ) ;
assign n15546 =  ( n14905 ) ? ( VREG_20_0 ) : ( n15545 ) ;
assign n15547 =  ( n14904 ) ? ( VREG_20_1 ) : ( n15546 ) ;
assign n15548 =  ( n14903 ) ? ( VREG_20_2 ) : ( n15547 ) ;
assign n15549 =  ( n14902 ) ? ( VREG_20_3 ) : ( n15548 ) ;
assign n15550 =  ( n14901 ) ? ( VREG_20_4 ) : ( n15549 ) ;
assign n15551 =  ( n14900 ) ? ( VREG_20_5 ) : ( n15550 ) ;
assign n15552 =  ( n14899 ) ? ( VREG_20_6 ) : ( n15551 ) ;
assign n15553 =  ( n14898 ) ? ( VREG_20_7 ) : ( n15552 ) ;
assign n15554 =  ( n14897 ) ? ( VREG_20_8 ) : ( n15553 ) ;
assign n15555 =  ( n14896 ) ? ( VREG_20_9 ) : ( n15554 ) ;
assign n15556 =  ( n14895 ) ? ( VREG_20_10 ) : ( n15555 ) ;
assign n15557 =  ( n14894 ) ? ( VREG_20_11 ) : ( n15556 ) ;
assign n15558 =  ( n14893 ) ? ( VREG_20_12 ) : ( n15557 ) ;
assign n15559 =  ( n14892 ) ? ( VREG_20_13 ) : ( n15558 ) ;
assign n15560 =  ( n14891 ) ? ( VREG_20_14 ) : ( n15559 ) ;
assign n15561 =  ( n14890 ) ? ( VREG_20_15 ) : ( n15560 ) ;
assign n15562 =  ( n14889 ) ? ( VREG_21_0 ) : ( n15561 ) ;
assign n15563 =  ( n14888 ) ? ( VREG_21_1 ) : ( n15562 ) ;
assign n15564 =  ( n14887 ) ? ( VREG_21_2 ) : ( n15563 ) ;
assign n15565 =  ( n14886 ) ? ( VREG_21_3 ) : ( n15564 ) ;
assign n15566 =  ( n14885 ) ? ( VREG_21_4 ) : ( n15565 ) ;
assign n15567 =  ( n14884 ) ? ( VREG_21_5 ) : ( n15566 ) ;
assign n15568 =  ( n14883 ) ? ( VREG_21_6 ) : ( n15567 ) ;
assign n15569 =  ( n14882 ) ? ( VREG_21_7 ) : ( n15568 ) ;
assign n15570 =  ( n14881 ) ? ( VREG_21_8 ) : ( n15569 ) ;
assign n15571 =  ( n14880 ) ? ( VREG_21_9 ) : ( n15570 ) ;
assign n15572 =  ( n14879 ) ? ( VREG_21_10 ) : ( n15571 ) ;
assign n15573 =  ( n14878 ) ? ( VREG_21_11 ) : ( n15572 ) ;
assign n15574 =  ( n14877 ) ? ( VREG_21_12 ) : ( n15573 ) ;
assign n15575 =  ( n14876 ) ? ( VREG_21_13 ) : ( n15574 ) ;
assign n15576 =  ( n14875 ) ? ( VREG_21_14 ) : ( n15575 ) ;
assign n15577 =  ( n14874 ) ? ( VREG_21_15 ) : ( n15576 ) ;
assign n15578 =  ( n14873 ) ? ( VREG_22_0 ) : ( n15577 ) ;
assign n15579 =  ( n14872 ) ? ( VREG_22_1 ) : ( n15578 ) ;
assign n15580 =  ( n14871 ) ? ( VREG_22_2 ) : ( n15579 ) ;
assign n15581 =  ( n14870 ) ? ( VREG_22_3 ) : ( n15580 ) ;
assign n15582 =  ( n14869 ) ? ( VREG_22_4 ) : ( n15581 ) ;
assign n15583 =  ( n14868 ) ? ( VREG_22_5 ) : ( n15582 ) ;
assign n15584 =  ( n14867 ) ? ( VREG_22_6 ) : ( n15583 ) ;
assign n15585 =  ( n14866 ) ? ( VREG_22_7 ) : ( n15584 ) ;
assign n15586 =  ( n14865 ) ? ( VREG_22_8 ) : ( n15585 ) ;
assign n15587 =  ( n14864 ) ? ( VREG_22_9 ) : ( n15586 ) ;
assign n15588 =  ( n14863 ) ? ( VREG_22_10 ) : ( n15587 ) ;
assign n15589 =  ( n14862 ) ? ( VREG_22_11 ) : ( n15588 ) ;
assign n15590 =  ( n14861 ) ? ( VREG_22_12 ) : ( n15589 ) ;
assign n15591 =  ( n14860 ) ? ( VREG_22_13 ) : ( n15590 ) ;
assign n15592 =  ( n14859 ) ? ( VREG_22_14 ) : ( n15591 ) ;
assign n15593 =  ( n14858 ) ? ( VREG_22_15 ) : ( n15592 ) ;
assign n15594 =  ( n14857 ) ? ( VREG_23_0 ) : ( n15593 ) ;
assign n15595 =  ( n14856 ) ? ( VREG_23_1 ) : ( n15594 ) ;
assign n15596 =  ( n14855 ) ? ( VREG_23_2 ) : ( n15595 ) ;
assign n15597 =  ( n14854 ) ? ( VREG_23_3 ) : ( n15596 ) ;
assign n15598 =  ( n14853 ) ? ( VREG_23_4 ) : ( n15597 ) ;
assign n15599 =  ( n14852 ) ? ( VREG_23_5 ) : ( n15598 ) ;
assign n15600 =  ( n14851 ) ? ( VREG_23_6 ) : ( n15599 ) ;
assign n15601 =  ( n14850 ) ? ( VREG_23_7 ) : ( n15600 ) ;
assign n15602 =  ( n14849 ) ? ( VREG_23_8 ) : ( n15601 ) ;
assign n15603 =  ( n14848 ) ? ( VREG_23_9 ) : ( n15602 ) ;
assign n15604 =  ( n14847 ) ? ( VREG_23_10 ) : ( n15603 ) ;
assign n15605 =  ( n14846 ) ? ( VREG_23_11 ) : ( n15604 ) ;
assign n15606 =  ( n14845 ) ? ( VREG_23_12 ) : ( n15605 ) ;
assign n15607 =  ( n14844 ) ? ( VREG_23_13 ) : ( n15606 ) ;
assign n15608 =  ( n14843 ) ? ( VREG_23_14 ) : ( n15607 ) ;
assign n15609 =  ( n14842 ) ? ( VREG_23_15 ) : ( n15608 ) ;
assign n15610 =  ( n14841 ) ? ( VREG_24_0 ) : ( n15609 ) ;
assign n15611 =  ( n14840 ) ? ( VREG_24_1 ) : ( n15610 ) ;
assign n15612 =  ( n14839 ) ? ( VREG_24_2 ) : ( n15611 ) ;
assign n15613 =  ( n14838 ) ? ( VREG_24_3 ) : ( n15612 ) ;
assign n15614 =  ( n14837 ) ? ( VREG_24_4 ) : ( n15613 ) ;
assign n15615 =  ( n14836 ) ? ( VREG_24_5 ) : ( n15614 ) ;
assign n15616 =  ( n14835 ) ? ( VREG_24_6 ) : ( n15615 ) ;
assign n15617 =  ( n14834 ) ? ( VREG_24_7 ) : ( n15616 ) ;
assign n15618 =  ( n14833 ) ? ( VREG_24_8 ) : ( n15617 ) ;
assign n15619 =  ( n14832 ) ? ( VREG_24_9 ) : ( n15618 ) ;
assign n15620 =  ( n14831 ) ? ( VREG_24_10 ) : ( n15619 ) ;
assign n15621 =  ( n14830 ) ? ( VREG_24_11 ) : ( n15620 ) ;
assign n15622 =  ( n14829 ) ? ( VREG_24_12 ) : ( n15621 ) ;
assign n15623 =  ( n14828 ) ? ( VREG_24_13 ) : ( n15622 ) ;
assign n15624 =  ( n14827 ) ? ( VREG_24_14 ) : ( n15623 ) ;
assign n15625 =  ( n14826 ) ? ( VREG_24_15 ) : ( n15624 ) ;
assign n15626 =  ( n14825 ) ? ( VREG_25_0 ) : ( n15625 ) ;
assign n15627 =  ( n14824 ) ? ( VREG_25_1 ) : ( n15626 ) ;
assign n15628 =  ( n14823 ) ? ( VREG_25_2 ) : ( n15627 ) ;
assign n15629 =  ( n14822 ) ? ( VREG_25_3 ) : ( n15628 ) ;
assign n15630 =  ( n14821 ) ? ( VREG_25_4 ) : ( n15629 ) ;
assign n15631 =  ( n14820 ) ? ( VREG_25_5 ) : ( n15630 ) ;
assign n15632 =  ( n14819 ) ? ( VREG_25_6 ) : ( n15631 ) ;
assign n15633 =  ( n14818 ) ? ( VREG_25_7 ) : ( n15632 ) ;
assign n15634 =  ( n14817 ) ? ( VREG_25_8 ) : ( n15633 ) ;
assign n15635 =  ( n14816 ) ? ( VREG_25_9 ) : ( n15634 ) ;
assign n15636 =  ( n14815 ) ? ( VREG_25_10 ) : ( n15635 ) ;
assign n15637 =  ( n14814 ) ? ( VREG_25_11 ) : ( n15636 ) ;
assign n15638 =  ( n14813 ) ? ( VREG_25_12 ) : ( n15637 ) ;
assign n15639 =  ( n14812 ) ? ( VREG_25_13 ) : ( n15638 ) ;
assign n15640 =  ( n14811 ) ? ( VREG_25_14 ) : ( n15639 ) ;
assign n15641 =  ( n14810 ) ? ( VREG_25_15 ) : ( n15640 ) ;
assign n15642 =  ( n14809 ) ? ( VREG_26_0 ) : ( n15641 ) ;
assign n15643 =  ( n14808 ) ? ( VREG_26_1 ) : ( n15642 ) ;
assign n15644 =  ( n14807 ) ? ( VREG_26_2 ) : ( n15643 ) ;
assign n15645 =  ( n14806 ) ? ( VREG_26_3 ) : ( n15644 ) ;
assign n15646 =  ( n14805 ) ? ( VREG_26_4 ) : ( n15645 ) ;
assign n15647 =  ( n14804 ) ? ( VREG_26_5 ) : ( n15646 ) ;
assign n15648 =  ( n14803 ) ? ( VREG_26_6 ) : ( n15647 ) ;
assign n15649 =  ( n14802 ) ? ( VREG_26_7 ) : ( n15648 ) ;
assign n15650 =  ( n14801 ) ? ( VREG_26_8 ) : ( n15649 ) ;
assign n15651 =  ( n14800 ) ? ( VREG_26_9 ) : ( n15650 ) ;
assign n15652 =  ( n14799 ) ? ( VREG_26_10 ) : ( n15651 ) ;
assign n15653 =  ( n14798 ) ? ( VREG_26_11 ) : ( n15652 ) ;
assign n15654 =  ( n14797 ) ? ( VREG_26_12 ) : ( n15653 ) ;
assign n15655 =  ( n14796 ) ? ( VREG_26_13 ) : ( n15654 ) ;
assign n15656 =  ( n14795 ) ? ( VREG_26_14 ) : ( n15655 ) ;
assign n15657 =  ( n14794 ) ? ( VREG_26_15 ) : ( n15656 ) ;
assign n15658 =  ( n14793 ) ? ( VREG_27_0 ) : ( n15657 ) ;
assign n15659 =  ( n14792 ) ? ( VREG_27_1 ) : ( n15658 ) ;
assign n15660 =  ( n14791 ) ? ( VREG_27_2 ) : ( n15659 ) ;
assign n15661 =  ( n14790 ) ? ( VREG_27_3 ) : ( n15660 ) ;
assign n15662 =  ( n14789 ) ? ( VREG_27_4 ) : ( n15661 ) ;
assign n15663 =  ( n14788 ) ? ( VREG_27_5 ) : ( n15662 ) ;
assign n15664 =  ( n14787 ) ? ( VREG_27_6 ) : ( n15663 ) ;
assign n15665 =  ( n14786 ) ? ( VREG_27_7 ) : ( n15664 ) ;
assign n15666 =  ( n14785 ) ? ( VREG_27_8 ) : ( n15665 ) ;
assign n15667 =  ( n14784 ) ? ( VREG_27_9 ) : ( n15666 ) ;
assign n15668 =  ( n14783 ) ? ( VREG_27_10 ) : ( n15667 ) ;
assign n15669 =  ( n14782 ) ? ( VREG_27_11 ) : ( n15668 ) ;
assign n15670 =  ( n14781 ) ? ( VREG_27_12 ) : ( n15669 ) ;
assign n15671 =  ( n14780 ) ? ( VREG_27_13 ) : ( n15670 ) ;
assign n15672 =  ( n14779 ) ? ( VREG_27_14 ) : ( n15671 ) ;
assign n15673 =  ( n14778 ) ? ( VREG_27_15 ) : ( n15672 ) ;
assign n15674 =  ( n14777 ) ? ( VREG_28_0 ) : ( n15673 ) ;
assign n15675 =  ( n14776 ) ? ( VREG_28_1 ) : ( n15674 ) ;
assign n15676 =  ( n14775 ) ? ( VREG_28_2 ) : ( n15675 ) ;
assign n15677 =  ( n14774 ) ? ( VREG_28_3 ) : ( n15676 ) ;
assign n15678 =  ( n14773 ) ? ( VREG_28_4 ) : ( n15677 ) ;
assign n15679 =  ( n14772 ) ? ( VREG_28_5 ) : ( n15678 ) ;
assign n15680 =  ( n14771 ) ? ( VREG_28_6 ) : ( n15679 ) ;
assign n15681 =  ( n14770 ) ? ( VREG_28_7 ) : ( n15680 ) ;
assign n15682 =  ( n14769 ) ? ( VREG_28_8 ) : ( n15681 ) ;
assign n15683 =  ( n14768 ) ? ( VREG_28_9 ) : ( n15682 ) ;
assign n15684 =  ( n14767 ) ? ( VREG_28_10 ) : ( n15683 ) ;
assign n15685 =  ( n14766 ) ? ( VREG_28_11 ) : ( n15684 ) ;
assign n15686 =  ( n14765 ) ? ( VREG_28_12 ) : ( n15685 ) ;
assign n15687 =  ( n14764 ) ? ( VREG_28_13 ) : ( n15686 ) ;
assign n15688 =  ( n14763 ) ? ( VREG_28_14 ) : ( n15687 ) ;
assign n15689 =  ( n14762 ) ? ( VREG_28_15 ) : ( n15688 ) ;
assign n15690 =  ( n14761 ) ? ( VREG_29_0 ) : ( n15689 ) ;
assign n15691 =  ( n14760 ) ? ( VREG_29_1 ) : ( n15690 ) ;
assign n15692 =  ( n14759 ) ? ( VREG_29_2 ) : ( n15691 ) ;
assign n15693 =  ( n14758 ) ? ( VREG_29_3 ) : ( n15692 ) ;
assign n15694 =  ( n14757 ) ? ( VREG_29_4 ) : ( n15693 ) ;
assign n15695 =  ( n14756 ) ? ( VREG_29_5 ) : ( n15694 ) ;
assign n15696 =  ( n14755 ) ? ( VREG_29_6 ) : ( n15695 ) ;
assign n15697 =  ( n14754 ) ? ( VREG_29_7 ) : ( n15696 ) ;
assign n15698 =  ( n14753 ) ? ( VREG_29_8 ) : ( n15697 ) ;
assign n15699 =  ( n14752 ) ? ( VREG_29_9 ) : ( n15698 ) ;
assign n15700 =  ( n14751 ) ? ( VREG_29_10 ) : ( n15699 ) ;
assign n15701 =  ( n14750 ) ? ( VREG_29_11 ) : ( n15700 ) ;
assign n15702 =  ( n14749 ) ? ( VREG_29_12 ) : ( n15701 ) ;
assign n15703 =  ( n14748 ) ? ( VREG_29_13 ) : ( n15702 ) ;
assign n15704 =  ( n14747 ) ? ( VREG_29_14 ) : ( n15703 ) ;
assign n15705 =  ( n14746 ) ? ( VREG_29_15 ) : ( n15704 ) ;
assign n15706 =  ( n14745 ) ? ( VREG_30_0 ) : ( n15705 ) ;
assign n15707 =  ( n14744 ) ? ( VREG_30_1 ) : ( n15706 ) ;
assign n15708 =  ( n14743 ) ? ( VREG_30_2 ) : ( n15707 ) ;
assign n15709 =  ( n14742 ) ? ( VREG_30_3 ) : ( n15708 ) ;
assign n15710 =  ( n14741 ) ? ( VREG_30_4 ) : ( n15709 ) ;
assign n15711 =  ( n14740 ) ? ( VREG_30_5 ) : ( n15710 ) ;
assign n15712 =  ( n14739 ) ? ( VREG_30_6 ) : ( n15711 ) ;
assign n15713 =  ( n14738 ) ? ( VREG_30_7 ) : ( n15712 ) ;
assign n15714 =  ( n14737 ) ? ( VREG_30_8 ) : ( n15713 ) ;
assign n15715 =  ( n14736 ) ? ( VREG_30_9 ) : ( n15714 ) ;
assign n15716 =  ( n14735 ) ? ( VREG_30_10 ) : ( n15715 ) ;
assign n15717 =  ( n14734 ) ? ( VREG_30_11 ) : ( n15716 ) ;
assign n15718 =  ( n14733 ) ? ( VREG_30_12 ) : ( n15717 ) ;
assign n15719 =  ( n14732 ) ? ( VREG_30_13 ) : ( n15718 ) ;
assign n15720 =  ( n14731 ) ? ( VREG_30_14 ) : ( n15719 ) ;
assign n15721 =  ( n14730 ) ? ( VREG_30_15 ) : ( n15720 ) ;
assign n15722 =  ( n14729 ) ? ( VREG_31_0 ) : ( n15721 ) ;
assign n15723 =  ( n14728 ) ? ( VREG_31_1 ) : ( n15722 ) ;
assign n15724 =  ( n14727 ) ? ( VREG_31_2 ) : ( n15723 ) ;
assign n15725 =  ( n14726 ) ? ( VREG_31_3 ) : ( n15724 ) ;
assign n15726 =  ( n14725 ) ? ( VREG_31_4 ) : ( n15725 ) ;
assign n15727 =  ( n14724 ) ? ( VREG_31_5 ) : ( n15726 ) ;
assign n15728 =  ( n14723 ) ? ( VREG_31_6 ) : ( n15727 ) ;
assign n15729 =  ( n14722 ) ? ( VREG_31_7 ) : ( n15728 ) ;
assign n15730 =  ( n14721 ) ? ( VREG_31_8 ) : ( n15729 ) ;
assign n15731 =  ( n14720 ) ? ( VREG_31_9 ) : ( n15730 ) ;
assign n15732 =  ( n14719 ) ? ( VREG_31_10 ) : ( n15731 ) ;
assign n15733 =  ( n14718 ) ? ( VREG_31_11 ) : ( n15732 ) ;
assign n15734 =  ( n14717 ) ? ( VREG_31_12 ) : ( n15733 ) ;
assign n15735 =  ( n14716 ) ? ( VREG_31_13 ) : ( n15734 ) ;
assign n15736 =  ( n14715 ) ? ( VREG_31_14 ) : ( n15735 ) ;
assign n15737 =  ( n14714 ) ? ( VREG_31_15 ) : ( n15736 ) ;
assign n15738 =  ( n14703 ) + ( n15737 )  ;
assign n15739 =  ( n14703 ) - ( n15737 )  ;
assign n15740 =  ( n14703 ) & ( n15737 )  ;
assign n15741 =  ( n14703 ) | ( n15737 )  ;
assign n15742 =  ( ( n14703 ) * ( n15737 ))  ;
assign n15743 =  ( n148 ) ? ( n15742 ) : ( VREG_0_14 ) ;
assign n15744 =  ( n146 ) ? ( n15741 ) : ( n15743 ) ;
assign n15745 =  ( n144 ) ? ( n15740 ) : ( n15744 ) ;
assign n15746 =  ( n142 ) ? ( n15739 ) : ( n15745 ) ;
assign n15747 =  ( n10 ) ? ( n15738 ) : ( n15746 ) ;
assign n15748 = n3030[14:14] ;
assign n15749 =  ( n15748 ) == ( 1'd0 )  ;
assign n15750 =  ( n15749 ) ? ( VREG_0_14 ) : ( n14713 ) ;
assign n15751 =  ( n15749 ) ? ( VREG_0_14 ) : ( n15747 ) ;
assign n15752 =  ( n3034 ) ? ( n15751 ) : ( VREG_0_14 ) ;
assign n15753 =  ( n2965 ) ? ( n15750 ) : ( n15752 ) ;
assign n15754 =  ( n1930 ) ? ( n15747 ) : ( n15753 ) ;
assign n15755 =  ( n879 ) ? ( n14713 ) : ( n15754 ) ;
assign n15756 =  ( n14703 ) + ( n164 )  ;
assign n15757 =  ( n14703 ) - ( n164 )  ;
assign n15758 =  ( n14703 ) & ( n164 )  ;
assign n15759 =  ( n14703 ) | ( n164 )  ;
assign n15760 =  ( ( n14703 ) * ( n164 ))  ;
assign n15761 =  ( n172 ) ? ( n15760 ) : ( VREG_0_14 ) ;
assign n15762 =  ( n170 ) ? ( n15759 ) : ( n15761 ) ;
assign n15763 =  ( n168 ) ? ( n15758 ) : ( n15762 ) ;
assign n15764 =  ( n166 ) ? ( n15757 ) : ( n15763 ) ;
assign n15765 =  ( n162 ) ? ( n15756 ) : ( n15764 ) ;
assign n15766 =  ( n14703 ) + ( n180 )  ;
assign n15767 =  ( n14703 ) - ( n180 )  ;
assign n15768 =  ( n14703 ) & ( n180 )  ;
assign n15769 =  ( n14703 ) | ( n180 )  ;
assign n15770 =  ( ( n14703 ) * ( n180 ))  ;
assign n15771 =  ( n172 ) ? ( n15770 ) : ( VREG_0_14 ) ;
assign n15772 =  ( n170 ) ? ( n15769 ) : ( n15771 ) ;
assign n15773 =  ( n168 ) ? ( n15768 ) : ( n15772 ) ;
assign n15774 =  ( n166 ) ? ( n15767 ) : ( n15773 ) ;
assign n15775 =  ( n162 ) ? ( n15766 ) : ( n15774 ) ;
assign n15776 =  ( n15749 ) ? ( VREG_0_14 ) : ( n15775 ) ;
assign n15777 =  ( n3051 ) ? ( n15776 ) : ( VREG_0_14 ) ;
assign n15778 =  ( n3040 ) ? ( n15765 ) : ( n15777 ) ;
assign n15779 =  ( n192 ) ? ( VREG_0_14 ) : ( VREG_0_14 ) ;
assign n15780 =  ( n157 ) ? ( n15778 ) : ( n15779 ) ;
assign n15781 =  ( n6 ) ? ( n15755 ) : ( n15780 ) ;
assign n15782 =  ( n4 ) ? ( n15781 ) : ( VREG_0_14 ) ;
assign n15783 =  ( 32'd15 ) == ( 32'd15 )  ;
assign n15784 =  ( n12 ) & ( n15783 )  ;
assign n15785 =  ( 32'd15 ) == ( 32'd14 )  ;
assign n15786 =  ( n12 ) & ( n15785 )  ;
assign n15787 =  ( 32'd15 ) == ( 32'd13 )  ;
assign n15788 =  ( n12 ) & ( n15787 )  ;
assign n15789 =  ( 32'd15 ) == ( 32'd12 )  ;
assign n15790 =  ( n12 ) & ( n15789 )  ;
assign n15791 =  ( 32'd15 ) == ( 32'd11 )  ;
assign n15792 =  ( n12 ) & ( n15791 )  ;
assign n15793 =  ( 32'd15 ) == ( 32'd10 )  ;
assign n15794 =  ( n12 ) & ( n15793 )  ;
assign n15795 =  ( 32'd15 ) == ( 32'd9 )  ;
assign n15796 =  ( n12 ) & ( n15795 )  ;
assign n15797 =  ( 32'd15 ) == ( 32'd8 )  ;
assign n15798 =  ( n12 ) & ( n15797 )  ;
assign n15799 =  ( 32'd15 ) == ( 32'd7 )  ;
assign n15800 =  ( n12 ) & ( n15799 )  ;
assign n15801 =  ( 32'd15 ) == ( 32'd6 )  ;
assign n15802 =  ( n12 ) & ( n15801 )  ;
assign n15803 =  ( 32'd15 ) == ( 32'd5 )  ;
assign n15804 =  ( n12 ) & ( n15803 )  ;
assign n15805 =  ( 32'd15 ) == ( 32'd4 )  ;
assign n15806 =  ( n12 ) & ( n15805 )  ;
assign n15807 =  ( 32'd15 ) == ( 32'd3 )  ;
assign n15808 =  ( n12 ) & ( n15807 )  ;
assign n15809 =  ( 32'd15 ) == ( 32'd2 )  ;
assign n15810 =  ( n12 ) & ( n15809 )  ;
assign n15811 =  ( 32'd15 ) == ( 32'd1 )  ;
assign n15812 =  ( n12 ) & ( n15811 )  ;
assign n15813 =  ( 32'd15 ) == ( 32'd0 )  ;
assign n15814 =  ( n12 ) & ( n15813 )  ;
assign n15815 =  ( n13 ) & ( n15783 )  ;
assign n15816 =  ( n13 ) & ( n15785 )  ;
assign n15817 =  ( n13 ) & ( n15787 )  ;
assign n15818 =  ( n13 ) & ( n15789 )  ;
assign n15819 =  ( n13 ) & ( n15791 )  ;
assign n15820 =  ( n13 ) & ( n15793 )  ;
assign n15821 =  ( n13 ) & ( n15795 )  ;
assign n15822 =  ( n13 ) & ( n15797 )  ;
assign n15823 =  ( n13 ) & ( n15799 )  ;
assign n15824 =  ( n13 ) & ( n15801 )  ;
assign n15825 =  ( n13 ) & ( n15803 )  ;
assign n15826 =  ( n13 ) & ( n15805 )  ;
assign n15827 =  ( n13 ) & ( n15807 )  ;
assign n15828 =  ( n13 ) & ( n15809 )  ;
assign n15829 =  ( n13 ) & ( n15811 )  ;
assign n15830 =  ( n13 ) & ( n15813 )  ;
assign n15831 =  ( n14 ) & ( n15783 )  ;
assign n15832 =  ( n14 ) & ( n15785 )  ;
assign n15833 =  ( n14 ) & ( n15787 )  ;
assign n15834 =  ( n14 ) & ( n15789 )  ;
assign n15835 =  ( n14 ) & ( n15791 )  ;
assign n15836 =  ( n14 ) & ( n15793 )  ;
assign n15837 =  ( n14 ) & ( n15795 )  ;
assign n15838 =  ( n14 ) & ( n15797 )  ;
assign n15839 =  ( n14 ) & ( n15799 )  ;
assign n15840 =  ( n14 ) & ( n15801 )  ;
assign n15841 =  ( n14 ) & ( n15803 )  ;
assign n15842 =  ( n14 ) & ( n15805 )  ;
assign n15843 =  ( n14 ) & ( n15807 )  ;
assign n15844 =  ( n14 ) & ( n15809 )  ;
assign n15845 =  ( n14 ) & ( n15811 )  ;
assign n15846 =  ( n14 ) & ( n15813 )  ;
assign n15847 =  ( n15 ) & ( n15783 )  ;
assign n15848 =  ( n15 ) & ( n15785 )  ;
assign n15849 =  ( n15 ) & ( n15787 )  ;
assign n15850 =  ( n15 ) & ( n15789 )  ;
assign n15851 =  ( n15 ) & ( n15791 )  ;
assign n15852 =  ( n15 ) & ( n15793 )  ;
assign n15853 =  ( n15 ) & ( n15795 )  ;
assign n15854 =  ( n15 ) & ( n15797 )  ;
assign n15855 =  ( n15 ) & ( n15799 )  ;
assign n15856 =  ( n15 ) & ( n15801 )  ;
assign n15857 =  ( n15 ) & ( n15803 )  ;
assign n15858 =  ( n15 ) & ( n15805 )  ;
assign n15859 =  ( n15 ) & ( n15807 )  ;
assign n15860 =  ( n15 ) & ( n15809 )  ;
assign n15861 =  ( n15 ) & ( n15811 )  ;
assign n15862 =  ( n15 ) & ( n15813 )  ;
assign n15863 =  ( n16 ) & ( n15783 )  ;
assign n15864 =  ( n16 ) & ( n15785 )  ;
assign n15865 =  ( n16 ) & ( n15787 )  ;
assign n15866 =  ( n16 ) & ( n15789 )  ;
assign n15867 =  ( n16 ) & ( n15791 )  ;
assign n15868 =  ( n16 ) & ( n15793 )  ;
assign n15869 =  ( n16 ) & ( n15795 )  ;
assign n15870 =  ( n16 ) & ( n15797 )  ;
assign n15871 =  ( n16 ) & ( n15799 )  ;
assign n15872 =  ( n16 ) & ( n15801 )  ;
assign n15873 =  ( n16 ) & ( n15803 )  ;
assign n15874 =  ( n16 ) & ( n15805 )  ;
assign n15875 =  ( n16 ) & ( n15807 )  ;
assign n15876 =  ( n16 ) & ( n15809 )  ;
assign n15877 =  ( n16 ) & ( n15811 )  ;
assign n15878 =  ( n16 ) & ( n15813 )  ;
assign n15879 =  ( n17 ) & ( n15783 )  ;
assign n15880 =  ( n17 ) & ( n15785 )  ;
assign n15881 =  ( n17 ) & ( n15787 )  ;
assign n15882 =  ( n17 ) & ( n15789 )  ;
assign n15883 =  ( n17 ) & ( n15791 )  ;
assign n15884 =  ( n17 ) & ( n15793 )  ;
assign n15885 =  ( n17 ) & ( n15795 )  ;
assign n15886 =  ( n17 ) & ( n15797 )  ;
assign n15887 =  ( n17 ) & ( n15799 )  ;
assign n15888 =  ( n17 ) & ( n15801 )  ;
assign n15889 =  ( n17 ) & ( n15803 )  ;
assign n15890 =  ( n17 ) & ( n15805 )  ;
assign n15891 =  ( n17 ) & ( n15807 )  ;
assign n15892 =  ( n17 ) & ( n15809 )  ;
assign n15893 =  ( n17 ) & ( n15811 )  ;
assign n15894 =  ( n17 ) & ( n15813 )  ;
assign n15895 =  ( n18 ) & ( n15783 )  ;
assign n15896 =  ( n18 ) & ( n15785 )  ;
assign n15897 =  ( n18 ) & ( n15787 )  ;
assign n15898 =  ( n18 ) & ( n15789 )  ;
assign n15899 =  ( n18 ) & ( n15791 )  ;
assign n15900 =  ( n18 ) & ( n15793 )  ;
assign n15901 =  ( n18 ) & ( n15795 )  ;
assign n15902 =  ( n18 ) & ( n15797 )  ;
assign n15903 =  ( n18 ) & ( n15799 )  ;
assign n15904 =  ( n18 ) & ( n15801 )  ;
assign n15905 =  ( n18 ) & ( n15803 )  ;
assign n15906 =  ( n18 ) & ( n15805 )  ;
assign n15907 =  ( n18 ) & ( n15807 )  ;
assign n15908 =  ( n18 ) & ( n15809 )  ;
assign n15909 =  ( n18 ) & ( n15811 )  ;
assign n15910 =  ( n18 ) & ( n15813 )  ;
assign n15911 =  ( n19 ) & ( n15783 )  ;
assign n15912 =  ( n19 ) & ( n15785 )  ;
assign n15913 =  ( n19 ) & ( n15787 )  ;
assign n15914 =  ( n19 ) & ( n15789 )  ;
assign n15915 =  ( n19 ) & ( n15791 )  ;
assign n15916 =  ( n19 ) & ( n15793 )  ;
assign n15917 =  ( n19 ) & ( n15795 )  ;
assign n15918 =  ( n19 ) & ( n15797 )  ;
assign n15919 =  ( n19 ) & ( n15799 )  ;
assign n15920 =  ( n19 ) & ( n15801 )  ;
assign n15921 =  ( n19 ) & ( n15803 )  ;
assign n15922 =  ( n19 ) & ( n15805 )  ;
assign n15923 =  ( n19 ) & ( n15807 )  ;
assign n15924 =  ( n19 ) & ( n15809 )  ;
assign n15925 =  ( n19 ) & ( n15811 )  ;
assign n15926 =  ( n19 ) & ( n15813 )  ;
assign n15927 =  ( n20 ) & ( n15783 )  ;
assign n15928 =  ( n20 ) & ( n15785 )  ;
assign n15929 =  ( n20 ) & ( n15787 )  ;
assign n15930 =  ( n20 ) & ( n15789 )  ;
assign n15931 =  ( n20 ) & ( n15791 )  ;
assign n15932 =  ( n20 ) & ( n15793 )  ;
assign n15933 =  ( n20 ) & ( n15795 )  ;
assign n15934 =  ( n20 ) & ( n15797 )  ;
assign n15935 =  ( n20 ) & ( n15799 )  ;
assign n15936 =  ( n20 ) & ( n15801 )  ;
assign n15937 =  ( n20 ) & ( n15803 )  ;
assign n15938 =  ( n20 ) & ( n15805 )  ;
assign n15939 =  ( n20 ) & ( n15807 )  ;
assign n15940 =  ( n20 ) & ( n15809 )  ;
assign n15941 =  ( n20 ) & ( n15811 )  ;
assign n15942 =  ( n20 ) & ( n15813 )  ;
assign n15943 =  ( n21 ) & ( n15783 )  ;
assign n15944 =  ( n21 ) & ( n15785 )  ;
assign n15945 =  ( n21 ) & ( n15787 )  ;
assign n15946 =  ( n21 ) & ( n15789 )  ;
assign n15947 =  ( n21 ) & ( n15791 )  ;
assign n15948 =  ( n21 ) & ( n15793 )  ;
assign n15949 =  ( n21 ) & ( n15795 )  ;
assign n15950 =  ( n21 ) & ( n15797 )  ;
assign n15951 =  ( n21 ) & ( n15799 )  ;
assign n15952 =  ( n21 ) & ( n15801 )  ;
assign n15953 =  ( n21 ) & ( n15803 )  ;
assign n15954 =  ( n21 ) & ( n15805 )  ;
assign n15955 =  ( n21 ) & ( n15807 )  ;
assign n15956 =  ( n21 ) & ( n15809 )  ;
assign n15957 =  ( n21 ) & ( n15811 )  ;
assign n15958 =  ( n21 ) & ( n15813 )  ;
assign n15959 =  ( n22 ) & ( n15783 )  ;
assign n15960 =  ( n22 ) & ( n15785 )  ;
assign n15961 =  ( n22 ) & ( n15787 )  ;
assign n15962 =  ( n22 ) & ( n15789 )  ;
assign n15963 =  ( n22 ) & ( n15791 )  ;
assign n15964 =  ( n22 ) & ( n15793 )  ;
assign n15965 =  ( n22 ) & ( n15795 )  ;
assign n15966 =  ( n22 ) & ( n15797 )  ;
assign n15967 =  ( n22 ) & ( n15799 )  ;
assign n15968 =  ( n22 ) & ( n15801 )  ;
assign n15969 =  ( n22 ) & ( n15803 )  ;
assign n15970 =  ( n22 ) & ( n15805 )  ;
assign n15971 =  ( n22 ) & ( n15807 )  ;
assign n15972 =  ( n22 ) & ( n15809 )  ;
assign n15973 =  ( n22 ) & ( n15811 )  ;
assign n15974 =  ( n22 ) & ( n15813 )  ;
assign n15975 =  ( n23 ) & ( n15783 )  ;
assign n15976 =  ( n23 ) & ( n15785 )  ;
assign n15977 =  ( n23 ) & ( n15787 )  ;
assign n15978 =  ( n23 ) & ( n15789 )  ;
assign n15979 =  ( n23 ) & ( n15791 )  ;
assign n15980 =  ( n23 ) & ( n15793 )  ;
assign n15981 =  ( n23 ) & ( n15795 )  ;
assign n15982 =  ( n23 ) & ( n15797 )  ;
assign n15983 =  ( n23 ) & ( n15799 )  ;
assign n15984 =  ( n23 ) & ( n15801 )  ;
assign n15985 =  ( n23 ) & ( n15803 )  ;
assign n15986 =  ( n23 ) & ( n15805 )  ;
assign n15987 =  ( n23 ) & ( n15807 )  ;
assign n15988 =  ( n23 ) & ( n15809 )  ;
assign n15989 =  ( n23 ) & ( n15811 )  ;
assign n15990 =  ( n23 ) & ( n15813 )  ;
assign n15991 =  ( n24 ) & ( n15783 )  ;
assign n15992 =  ( n24 ) & ( n15785 )  ;
assign n15993 =  ( n24 ) & ( n15787 )  ;
assign n15994 =  ( n24 ) & ( n15789 )  ;
assign n15995 =  ( n24 ) & ( n15791 )  ;
assign n15996 =  ( n24 ) & ( n15793 )  ;
assign n15997 =  ( n24 ) & ( n15795 )  ;
assign n15998 =  ( n24 ) & ( n15797 )  ;
assign n15999 =  ( n24 ) & ( n15799 )  ;
assign n16000 =  ( n24 ) & ( n15801 )  ;
assign n16001 =  ( n24 ) & ( n15803 )  ;
assign n16002 =  ( n24 ) & ( n15805 )  ;
assign n16003 =  ( n24 ) & ( n15807 )  ;
assign n16004 =  ( n24 ) & ( n15809 )  ;
assign n16005 =  ( n24 ) & ( n15811 )  ;
assign n16006 =  ( n24 ) & ( n15813 )  ;
assign n16007 =  ( n25 ) & ( n15783 )  ;
assign n16008 =  ( n25 ) & ( n15785 )  ;
assign n16009 =  ( n25 ) & ( n15787 )  ;
assign n16010 =  ( n25 ) & ( n15789 )  ;
assign n16011 =  ( n25 ) & ( n15791 )  ;
assign n16012 =  ( n25 ) & ( n15793 )  ;
assign n16013 =  ( n25 ) & ( n15795 )  ;
assign n16014 =  ( n25 ) & ( n15797 )  ;
assign n16015 =  ( n25 ) & ( n15799 )  ;
assign n16016 =  ( n25 ) & ( n15801 )  ;
assign n16017 =  ( n25 ) & ( n15803 )  ;
assign n16018 =  ( n25 ) & ( n15805 )  ;
assign n16019 =  ( n25 ) & ( n15807 )  ;
assign n16020 =  ( n25 ) & ( n15809 )  ;
assign n16021 =  ( n25 ) & ( n15811 )  ;
assign n16022 =  ( n25 ) & ( n15813 )  ;
assign n16023 =  ( n26 ) & ( n15783 )  ;
assign n16024 =  ( n26 ) & ( n15785 )  ;
assign n16025 =  ( n26 ) & ( n15787 )  ;
assign n16026 =  ( n26 ) & ( n15789 )  ;
assign n16027 =  ( n26 ) & ( n15791 )  ;
assign n16028 =  ( n26 ) & ( n15793 )  ;
assign n16029 =  ( n26 ) & ( n15795 )  ;
assign n16030 =  ( n26 ) & ( n15797 )  ;
assign n16031 =  ( n26 ) & ( n15799 )  ;
assign n16032 =  ( n26 ) & ( n15801 )  ;
assign n16033 =  ( n26 ) & ( n15803 )  ;
assign n16034 =  ( n26 ) & ( n15805 )  ;
assign n16035 =  ( n26 ) & ( n15807 )  ;
assign n16036 =  ( n26 ) & ( n15809 )  ;
assign n16037 =  ( n26 ) & ( n15811 )  ;
assign n16038 =  ( n26 ) & ( n15813 )  ;
assign n16039 =  ( n27 ) & ( n15783 )  ;
assign n16040 =  ( n27 ) & ( n15785 )  ;
assign n16041 =  ( n27 ) & ( n15787 )  ;
assign n16042 =  ( n27 ) & ( n15789 )  ;
assign n16043 =  ( n27 ) & ( n15791 )  ;
assign n16044 =  ( n27 ) & ( n15793 )  ;
assign n16045 =  ( n27 ) & ( n15795 )  ;
assign n16046 =  ( n27 ) & ( n15797 )  ;
assign n16047 =  ( n27 ) & ( n15799 )  ;
assign n16048 =  ( n27 ) & ( n15801 )  ;
assign n16049 =  ( n27 ) & ( n15803 )  ;
assign n16050 =  ( n27 ) & ( n15805 )  ;
assign n16051 =  ( n27 ) & ( n15807 )  ;
assign n16052 =  ( n27 ) & ( n15809 )  ;
assign n16053 =  ( n27 ) & ( n15811 )  ;
assign n16054 =  ( n27 ) & ( n15813 )  ;
assign n16055 =  ( n28 ) & ( n15783 )  ;
assign n16056 =  ( n28 ) & ( n15785 )  ;
assign n16057 =  ( n28 ) & ( n15787 )  ;
assign n16058 =  ( n28 ) & ( n15789 )  ;
assign n16059 =  ( n28 ) & ( n15791 )  ;
assign n16060 =  ( n28 ) & ( n15793 )  ;
assign n16061 =  ( n28 ) & ( n15795 )  ;
assign n16062 =  ( n28 ) & ( n15797 )  ;
assign n16063 =  ( n28 ) & ( n15799 )  ;
assign n16064 =  ( n28 ) & ( n15801 )  ;
assign n16065 =  ( n28 ) & ( n15803 )  ;
assign n16066 =  ( n28 ) & ( n15805 )  ;
assign n16067 =  ( n28 ) & ( n15807 )  ;
assign n16068 =  ( n28 ) & ( n15809 )  ;
assign n16069 =  ( n28 ) & ( n15811 )  ;
assign n16070 =  ( n28 ) & ( n15813 )  ;
assign n16071 =  ( n29 ) & ( n15783 )  ;
assign n16072 =  ( n29 ) & ( n15785 )  ;
assign n16073 =  ( n29 ) & ( n15787 )  ;
assign n16074 =  ( n29 ) & ( n15789 )  ;
assign n16075 =  ( n29 ) & ( n15791 )  ;
assign n16076 =  ( n29 ) & ( n15793 )  ;
assign n16077 =  ( n29 ) & ( n15795 )  ;
assign n16078 =  ( n29 ) & ( n15797 )  ;
assign n16079 =  ( n29 ) & ( n15799 )  ;
assign n16080 =  ( n29 ) & ( n15801 )  ;
assign n16081 =  ( n29 ) & ( n15803 )  ;
assign n16082 =  ( n29 ) & ( n15805 )  ;
assign n16083 =  ( n29 ) & ( n15807 )  ;
assign n16084 =  ( n29 ) & ( n15809 )  ;
assign n16085 =  ( n29 ) & ( n15811 )  ;
assign n16086 =  ( n29 ) & ( n15813 )  ;
assign n16087 =  ( n30 ) & ( n15783 )  ;
assign n16088 =  ( n30 ) & ( n15785 )  ;
assign n16089 =  ( n30 ) & ( n15787 )  ;
assign n16090 =  ( n30 ) & ( n15789 )  ;
assign n16091 =  ( n30 ) & ( n15791 )  ;
assign n16092 =  ( n30 ) & ( n15793 )  ;
assign n16093 =  ( n30 ) & ( n15795 )  ;
assign n16094 =  ( n30 ) & ( n15797 )  ;
assign n16095 =  ( n30 ) & ( n15799 )  ;
assign n16096 =  ( n30 ) & ( n15801 )  ;
assign n16097 =  ( n30 ) & ( n15803 )  ;
assign n16098 =  ( n30 ) & ( n15805 )  ;
assign n16099 =  ( n30 ) & ( n15807 )  ;
assign n16100 =  ( n30 ) & ( n15809 )  ;
assign n16101 =  ( n30 ) & ( n15811 )  ;
assign n16102 =  ( n30 ) & ( n15813 )  ;
assign n16103 =  ( n31 ) & ( n15783 )  ;
assign n16104 =  ( n31 ) & ( n15785 )  ;
assign n16105 =  ( n31 ) & ( n15787 )  ;
assign n16106 =  ( n31 ) & ( n15789 )  ;
assign n16107 =  ( n31 ) & ( n15791 )  ;
assign n16108 =  ( n31 ) & ( n15793 )  ;
assign n16109 =  ( n31 ) & ( n15795 )  ;
assign n16110 =  ( n31 ) & ( n15797 )  ;
assign n16111 =  ( n31 ) & ( n15799 )  ;
assign n16112 =  ( n31 ) & ( n15801 )  ;
assign n16113 =  ( n31 ) & ( n15803 )  ;
assign n16114 =  ( n31 ) & ( n15805 )  ;
assign n16115 =  ( n31 ) & ( n15807 )  ;
assign n16116 =  ( n31 ) & ( n15809 )  ;
assign n16117 =  ( n31 ) & ( n15811 )  ;
assign n16118 =  ( n31 ) & ( n15813 )  ;
assign n16119 =  ( n32 ) & ( n15783 )  ;
assign n16120 =  ( n32 ) & ( n15785 )  ;
assign n16121 =  ( n32 ) & ( n15787 )  ;
assign n16122 =  ( n32 ) & ( n15789 )  ;
assign n16123 =  ( n32 ) & ( n15791 )  ;
assign n16124 =  ( n32 ) & ( n15793 )  ;
assign n16125 =  ( n32 ) & ( n15795 )  ;
assign n16126 =  ( n32 ) & ( n15797 )  ;
assign n16127 =  ( n32 ) & ( n15799 )  ;
assign n16128 =  ( n32 ) & ( n15801 )  ;
assign n16129 =  ( n32 ) & ( n15803 )  ;
assign n16130 =  ( n32 ) & ( n15805 )  ;
assign n16131 =  ( n32 ) & ( n15807 )  ;
assign n16132 =  ( n32 ) & ( n15809 )  ;
assign n16133 =  ( n32 ) & ( n15811 )  ;
assign n16134 =  ( n32 ) & ( n15813 )  ;
assign n16135 =  ( n33 ) & ( n15783 )  ;
assign n16136 =  ( n33 ) & ( n15785 )  ;
assign n16137 =  ( n33 ) & ( n15787 )  ;
assign n16138 =  ( n33 ) & ( n15789 )  ;
assign n16139 =  ( n33 ) & ( n15791 )  ;
assign n16140 =  ( n33 ) & ( n15793 )  ;
assign n16141 =  ( n33 ) & ( n15795 )  ;
assign n16142 =  ( n33 ) & ( n15797 )  ;
assign n16143 =  ( n33 ) & ( n15799 )  ;
assign n16144 =  ( n33 ) & ( n15801 )  ;
assign n16145 =  ( n33 ) & ( n15803 )  ;
assign n16146 =  ( n33 ) & ( n15805 )  ;
assign n16147 =  ( n33 ) & ( n15807 )  ;
assign n16148 =  ( n33 ) & ( n15809 )  ;
assign n16149 =  ( n33 ) & ( n15811 )  ;
assign n16150 =  ( n33 ) & ( n15813 )  ;
assign n16151 =  ( n34 ) & ( n15783 )  ;
assign n16152 =  ( n34 ) & ( n15785 )  ;
assign n16153 =  ( n34 ) & ( n15787 )  ;
assign n16154 =  ( n34 ) & ( n15789 )  ;
assign n16155 =  ( n34 ) & ( n15791 )  ;
assign n16156 =  ( n34 ) & ( n15793 )  ;
assign n16157 =  ( n34 ) & ( n15795 )  ;
assign n16158 =  ( n34 ) & ( n15797 )  ;
assign n16159 =  ( n34 ) & ( n15799 )  ;
assign n16160 =  ( n34 ) & ( n15801 )  ;
assign n16161 =  ( n34 ) & ( n15803 )  ;
assign n16162 =  ( n34 ) & ( n15805 )  ;
assign n16163 =  ( n34 ) & ( n15807 )  ;
assign n16164 =  ( n34 ) & ( n15809 )  ;
assign n16165 =  ( n34 ) & ( n15811 )  ;
assign n16166 =  ( n34 ) & ( n15813 )  ;
assign n16167 =  ( n35 ) & ( n15783 )  ;
assign n16168 =  ( n35 ) & ( n15785 )  ;
assign n16169 =  ( n35 ) & ( n15787 )  ;
assign n16170 =  ( n35 ) & ( n15789 )  ;
assign n16171 =  ( n35 ) & ( n15791 )  ;
assign n16172 =  ( n35 ) & ( n15793 )  ;
assign n16173 =  ( n35 ) & ( n15795 )  ;
assign n16174 =  ( n35 ) & ( n15797 )  ;
assign n16175 =  ( n35 ) & ( n15799 )  ;
assign n16176 =  ( n35 ) & ( n15801 )  ;
assign n16177 =  ( n35 ) & ( n15803 )  ;
assign n16178 =  ( n35 ) & ( n15805 )  ;
assign n16179 =  ( n35 ) & ( n15807 )  ;
assign n16180 =  ( n35 ) & ( n15809 )  ;
assign n16181 =  ( n35 ) & ( n15811 )  ;
assign n16182 =  ( n35 ) & ( n15813 )  ;
assign n16183 =  ( n36 ) & ( n15783 )  ;
assign n16184 =  ( n36 ) & ( n15785 )  ;
assign n16185 =  ( n36 ) & ( n15787 )  ;
assign n16186 =  ( n36 ) & ( n15789 )  ;
assign n16187 =  ( n36 ) & ( n15791 )  ;
assign n16188 =  ( n36 ) & ( n15793 )  ;
assign n16189 =  ( n36 ) & ( n15795 )  ;
assign n16190 =  ( n36 ) & ( n15797 )  ;
assign n16191 =  ( n36 ) & ( n15799 )  ;
assign n16192 =  ( n36 ) & ( n15801 )  ;
assign n16193 =  ( n36 ) & ( n15803 )  ;
assign n16194 =  ( n36 ) & ( n15805 )  ;
assign n16195 =  ( n36 ) & ( n15807 )  ;
assign n16196 =  ( n36 ) & ( n15809 )  ;
assign n16197 =  ( n36 ) & ( n15811 )  ;
assign n16198 =  ( n36 ) & ( n15813 )  ;
assign n16199 =  ( n37 ) & ( n15783 )  ;
assign n16200 =  ( n37 ) & ( n15785 )  ;
assign n16201 =  ( n37 ) & ( n15787 )  ;
assign n16202 =  ( n37 ) & ( n15789 )  ;
assign n16203 =  ( n37 ) & ( n15791 )  ;
assign n16204 =  ( n37 ) & ( n15793 )  ;
assign n16205 =  ( n37 ) & ( n15795 )  ;
assign n16206 =  ( n37 ) & ( n15797 )  ;
assign n16207 =  ( n37 ) & ( n15799 )  ;
assign n16208 =  ( n37 ) & ( n15801 )  ;
assign n16209 =  ( n37 ) & ( n15803 )  ;
assign n16210 =  ( n37 ) & ( n15805 )  ;
assign n16211 =  ( n37 ) & ( n15807 )  ;
assign n16212 =  ( n37 ) & ( n15809 )  ;
assign n16213 =  ( n37 ) & ( n15811 )  ;
assign n16214 =  ( n37 ) & ( n15813 )  ;
assign n16215 =  ( n38 ) & ( n15783 )  ;
assign n16216 =  ( n38 ) & ( n15785 )  ;
assign n16217 =  ( n38 ) & ( n15787 )  ;
assign n16218 =  ( n38 ) & ( n15789 )  ;
assign n16219 =  ( n38 ) & ( n15791 )  ;
assign n16220 =  ( n38 ) & ( n15793 )  ;
assign n16221 =  ( n38 ) & ( n15795 )  ;
assign n16222 =  ( n38 ) & ( n15797 )  ;
assign n16223 =  ( n38 ) & ( n15799 )  ;
assign n16224 =  ( n38 ) & ( n15801 )  ;
assign n16225 =  ( n38 ) & ( n15803 )  ;
assign n16226 =  ( n38 ) & ( n15805 )  ;
assign n16227 =  ( n38 ) & ( n15807 )  ;
assign n16228 =  ( n38 ) & ( n15809 )  ;
assign n16229 =  ( n38 ) & ( n15811 )  ;
assign n16230 =  ( n38 ) & ( n15813 )  ;
assign n16231 =  ( n39 ) & ( n15783 )  ;
assign n16232 =  ( n39 ) & ( n15785 )  ;
assign n16233 =  ( n39 ) & ( n15787 )  ;
assign n16234 =  ( n39 ) & ( n15789 )  ;
assign n16235 =  ( n39 ) & ( n15791 )  ;
assign n16236 =  ( n39 ) & ( n15793 )  ;
assign n16237 =  ( n39 ) & ( n15795 )  ;
assign n16238 =  ( n39 ) & ( n15797 )  ;
assign n16239 =  ( n39 ) & ( n15799 )  ;
assign n16240 =  ( n39 ) & ( n15801 )  ;
assign n16241 =  ( n39 ) & ( n15803 )  ;
assign n16242 =  ( n39 ) & ( n15805 )  ;
assign n16243 =  ( n39 ) & ( n15807 )  ;
assign n16244 =  ( n39 ) & ( n15809 )  ;
assign n16245 =  ( n39 ) & ( n15811 )  ;
assign n16246 =  ( n39 ) & ( n15813 )  ;
assign n16247 =  ( n40 ) & ( n15783 )  ;
assign n16248 =  ( n40 ) & ( n15785 )  ;
assign n16249 =  ( n40 ) & ( n15787 )  ;
assign n16250 =  ( n40 ) & ( n15789 )  ;
assign n16251 =  ( n40 ) & ( n15791 )  ;
assign n16252 =  ( n40 ) & ( n15793 )  ;
assign n16253 =  ( n40 ) & ( n15795 )  ;
assign n16254 =  ( n40 ) & ( n15797 )  ;
assign n16255 =  ( n40 ) & ( n15799 )  ;
assign n16256 =  ( n40 ) & ( n15801 )  ;
assign n16257 =  ( n40 ) & ( n15803 )  ;
assign n16258 =  ( n40 ) & ( n15805 )  ;
assign n16259 =  ( n40 ) & ( n15807 )  ;
assign n16260 =  ( n40 ) & ( n15809 )  ;
assign n16261 =  ( n40 ) & ( n15811 )  ;
assign n16262 =  ( n40 ) & ( n15813 )  ;
assign n16263 =  ( n41 ) & ( n15783 )  ;
assign n16264 =  ( n41 ) & ( n15785 )  ;
assign n16265 =  ( n41 ) & ( n15787 )  ;
assign n16266 =  ( n41 ) & ( n15789 )  ;
assign n16267 =  ( n41 ) & ( n15791 )  ;
assign n16268 =  ( n41 ) & ( n15793 )  ;
assign n16269 =  ( n41 ) & ( n15795 )  ;
assign n16270 =  ( n41 ) & ( n15797 )  ;
assign n16271 =  ( n41 ) & ( n15799 )  ;
assign n16272 =  ( n41 ) & ( n15801 )  ;
assign n16273 =  ( n41 ) & ( n15803 )  ;
assign n16274 =  ( n41 ) & ( n15805 )  ;
assign n16275 =  ( n41 ) & ( n15807 )  ;
assign n16276 =  ( n41 ) & ( n15809 )  ;
assign n16277 =  ( n41 ) & ( n15811 )  ;
assign n16278 =  ( n41 ) & ( n15813 )  ;
assign n16279 =  ( n42 ) & ( n15783 )  ;
assign n16280 =  ( n42 ) & ( n15785 )  ;
assign n16281 =  ( n42 ) & ( n15787 )  ;
assign n16282 =  ( n42 ) & ( n15789 )  ;
assign n16283 =  ( n42 ) & ( n15791 )  ;
assign n16284 =  ( n42 ) & ( n15793 )  ;
assign n16285 =  ( n42 ) & ( n15795 )  ;
assign n16286 =  ( n42 ) & ( n15797 )  ;
assign n16287 =  ( n42 ) & ( n15799 )  ;
assign n16288 =  ( n42 ) & ( n15801 )  ;
assign n16289 =  ( n42 ) & ( n15803 )  ;
assign n16290 =  ( n42 ) & ( n15805 )  ;
assign n16291 =  ( n42 ) & ( n15807 )  ;
assign n16292 =  ( n42 ) & ( n15809 )  ;
assign n16293 =  ( n42 ) & ( n15811 )  ;
assign n16294 =  ( n42 ) & ( n15813 )  ;
assign n16295 =  ( n43 ) & ( n15783 )  ;
assign n16296 =  ( n43 ) & ( n15785 )  ;
assign n16297 =  ( n43 ) & ( n15787 )  ;
assign n16298 =  ( n43 ) & ( n15789 )  ;
assign n16299 =  ( n43 ) & ( n15791 )  ;
assign n16300 =  ( n43 ) & ( n15793 )  ;
assign n16301 =  ( n43 ) & ( n15795 )  ;
assign n16302 =  ( n43 ) & ( n15797 )  ;
assign n16303 =  ( n43 ) & ( n15799 )  ;
assign n16304 =  ( n43 ) & ( n15801 )  ;
assign n16305 =  ( n43 ) & ( n15803 )  ;
assign n16306 =  ( n43 ) & ( n15805 )  ;
assign n16307 =  ( n43 ) & ( n15807 )  ;
assign n16308 =  ( n43 ) & ( n15809 )  ;
assign n16309 =  ( n43 ) & ( n15811 )  ;
assign n16310 =  ( n43 ) & ( n15813 )  ;
assign n16311 =  ( n16310 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n16312 =  ( n16309 ) ? ( VREG_0_1 ) : ( n16311 ) ;
assign n16313 =  ( n16308 ) ? ( VREG_0_2 ) : ( n16312 ) ;
assign n16314 =  ( n16307 ) ? ( VREG_0_3 ) : ( n16313 ) ;
assign n16315 =  ( n16306 ) ? ( VREG_0_4 ) : ( n16314 ) ;
assign n16316 =  ( n16305 ) ? ( VREG_0_5 ) : ( n16315 ) ;
assign n16317 =  ( n16304 ) ? ( VREG_0_6 ) : ( n16316 ) ;
assign n16318 =  ( n16303 ) ? ( VREG_0_7 ) : ( n16317 ) ;
assign n16319 =  ( n16302 ) ? ( VREG_0_8 ) : ( n16318 ) ;
assign n16320 =  ( n16301 ) ? ( VREG_0_9 ) : ( n16319 ) ;
assign n16321 =  ( n16300 ) ? ( VREG_0_10 ) : ( n16320 ) ;
assign n16322 =  ( n16299 ) ? ( VREG_0_11 ) : ( n16321 ) ;
assign n16323 =  ( n16298 ) ? ( VREG_0_12 ) : ( n16322 ) ;
assign n16324 =  ( n16297 ) ? ( VREG_0_13 ) : ( n16323 ) ;
assign n16325 =  ( n16296 ) ? ( VREG_0_14 ) : ( n16324 ) ;
assign n16326 =  ( n16295 ) ? ( VREG_0_15 ) : ( n16325 ) ;
assign n16327 =  ( n16294 ) ? ( VREG_1_0 ) : ( n16326 ) ;
assign n16328 =  ( n16293 ) ? ( VREG_1_1 ) : ( n16327 ) ;
assign n16329 =  ( n16292 ) ? ( VREG_1_2 ) : ( n16328 ) ;
assign n16330 =  ( n16291 ) ? ( VREG_1_3 ) : ( n16329 ) ;
assign n16331 =  ( n16290 ) ? ( VREG_1_4 ) : ( n16330 ) ;
assign n16332 =  ( n16289 ) ? ( VREG_1_5 ) : ( n16331 ) ;
assign n16333 =  ( n16288 ) ? ( VREG_1_6 ) : ( n16332 ) ;
assign n16334 =  ( n16287 ) ? ( VREG_1_7 ) : ( n16333 ) ;
assign n16335 =  ( n16286 ) ? ( VREG_1_8 ) : ( n16334 ) ;
assign n16336 =  ( n16285 ) ? ( VREG_1_9 ) : ( n16335 ) ;
assign n16337 =  ( n16284 ) ? ( VREG_1_10 ) : ( n16336 ) ;
assign n16338 =  ( n16283 ) ? ( VREG_1_11 ) : ( n16337 ) ;
assign n16339 =  ( n16282 ) ? ( VREG_1_12 ) : ( n16338 ) ;
assign n16340 =  ( n16281 ) ? ( VREG_1_13 ) : ( n16339 ) ;
assign n16341 =  ( n16280 ) ? ( VREG_1_14 ) : ( n16340 ) ;
assign n16342 =  ( n16279 ) ? ( VREG_1_15 ) : ( n16341 ) ;
assign n16343 =  ( n16278 ) ? ( VREG_2_0 ) : ( n16342 ) ;
assign n16344 =  ( n16277 ) ? ( VREG_2_1 ) : ( n16343 ) ;
assign n16345 =  ( n16276 ) ? ( VREG_2_2 ) : ( n16344 ) ;
assign n16346 =  ( n16275 ) ? ( VREG_2_3 ) : ( n16345 ) ;
assign n16347 =  ( n16274 ) ? ( VREG_2_4 ) : ( n16346 ) ;
assign n16348 =  ( n16273 ) ? ( VREG_2_5 ) : ( n16347 ) ;
assign n16349 =  ( n16272 ) ? ( VREG_2_6 ) : ( n16348 ) ;
assign n16350 =  ( n16271 ) ? ( VREG_2_7 ) : ( n16349 ) ;
assign n16351 =  ( n16270 ) ? ( VREG_2_8 ) : ( n16350 ) ;
assign n16352 =  ( n16269 ) ? ( VREG_2_9 ) : ( n16351 ) ;
assign n16353 =  ( n16268 ) ? ( VREG_2_10 ) : ( n16352 ) ;
assign n16354 =  ( n16267 ) ? ( VREG_2_11 ) : ( n16353 ) ;
assign n16355 =  ( n16266 ) ? ( VREG_2_12 ) : ( n16354 ) ;
assign n16356 =  ( n16265 ) ? ( VREG_2_13 ) : ( n16355 ) ;
assign n16357 =  ( n16264 ) ? ( VREG_2_14 ) : ( n16356 ) ;
assign n16358 =  ( n16263 ) ? ( VREG_2_15 ) : ( n16357 ) ;
assign n16359 =  ( n16262 ) ? ( VREG_3_0 ) : ( n16358 ) ;
assign n16360 =  ( n16261 ) ? ( VREG_3_1 ) : ( n16359 ) ;
assign n16361 =  ( n16260 ) ? ( VREG_3_2 ) : ( n16360 ) ;
assign n16362 =  ( n16259 ) ? ( VREG_3_3 ) : ( n16361 ) ;
assign n16363 =  ( n16258 ) ? ( VREG_3_4 ) : ( n16362 ) ;
assign n16364 =  ( n16257 ) ? ( VREG_3_5 ) : ( n16363 ) ;
assign n16365 =  ( n16256 ) ? ( VREG_3_6 ) : ( n16364 ) ;
assign n16366 =  ( n16255 ) ? ( VREG_3_7 ) : ( n16365 ) ;
assign n16367 =  ( n16254 ) ? ( VREG_3_8 ) : ( n16366 ) ;
assign n16368 =  ( n16253 ) ? ( VREG_3_9 ) : ( n16367 ) ;
assign n16369 =  ( n16252 ) ? ( VREG_3_10 ) : ( n16368 ) ;
assign n16370 =  ( n16251 ) ? ( VREG_3_11 ) : ( n16369 ) ;
assign n16371 =  ( n16250 ) ? ( VREG_3_12 ) : ( n16370 ) ;
assign n16372 =  ( n16249 ) ? ( VREG_3_13 ) : ( n16371 ) ;
assign n16373 =  ( n16248 ) ? ( VREG_3_14 ) : ( n16372 ) ;
assign n16374 =  ( n16247 ) ? ( VREG_3_15 ) : ( n16373 ) ;
assign n16375 =  ( n16246 ) ? ( VREG_4_0 ) : ( n16374 ) ;
assign n16376 =  ( n16245 ) ? ( VREG_4_1 ) : ( n16375 ) ;
assign n16377 =  ( n16244 ) ? ( VREG_4_2 ) : ( n16376 ) ;
assign n16378 =  ( n16243 ) ? ( VREG_4_3 ) : ( n16377 ) ;
assign n16379 =  ( n16242 ) ? ( VREG_4_4 ) : ( n16378 ) ;
assign n16380 =  ( n16241 ) ? ( VREG_4_5 ) : ( n16379 ) ;
assign n16381 =  ( n16240 ) ? ( VREG_4_6 ) : ( n16380 ) ;
assign n16382 =  ( n16239 ) ? ( VREG_4_7 ) : ( n16381 ) ;
assign n16383 =  ( n16238 ) ? ( VREG_4_8 ) : ( n16382 ) ;
assign n16384 =  ( n16237 ) ? ( VREG_4_9 ) : ( n16383 ) ;
assign n16385 =  ( n16236 ) ? ( VREG_4_10 ) : ( n16384 ) ;
assign n16386 =  ( n16235 ) ? ( VREG_4_11 ) : ( n16385 ) ;
assign n16387 =  ( n16234 ) ? ( VREG_4_12 ) : ( n16386 ) ;
assign n16388 =  ( n16233 ) ? ( VREG_4_13 ) : ( n16387 ) ;
assign n16389 =  ( n16232 ) ? ( VREG_4_14 ) : ( n16388 ) ;
assign n16390 =  ( n16231 ) ? ( VREG_4_15 ) : ( n16389 ) ;
assign n16391 =  ( n16230 ) ? ( VREG_5_0 ) : ( n16390 ) ;
assign n16392 =  ( n16229 ) ? ( VREG_5_1 ) : ( n16391 ) ;
assign n16393 =  ( n16228 ) ? ( VREG_5_2 ) : ( n16392 ) ;
assign n16394 =  ( n16227 ) ? ( VREG_5_3 ) : ( n16393 ) ;
assign n16395 =  ( n16226 ) ? ( VREG_5_4 ) : ( n16394 ) ;
assign n16396 =  ( n16225 ) ? ( VREG_5_5 ) : ( n16395 ) ;
assign n16397 =  ( n16224 ) ? ( VREG_5_6 ) : ( n16396 ) ;
assign n16398 =  ( n16223 ) ? ( VREG_5_7 ) : ( n16397 ) ;
assign n16399 =  ( n16222 ) ? ( VREG_5_8 ) : ( n16398 ) ;
assign n16400 =  ( n16221 ) ? ( VREG_5_9 ) : ( n16399 ) ;
assign n16401 =  ( n16220 ) ? ( VREG_5_10 ) : ( n16400 ) ;
assign n16402 =  ( n16219 ) ? ( VREG_5_11 ) : ( n16401 ) ;
assign n16403 =  ( n16218 ) ? ( VREG_5_12 ) : ( n16402 ) ;
assign n16404 =  ( n16217 ) ? ( VREG_5_13 ) : ( n16403 ) ;
assign n16405 =  ( n16216 ) ? ( VREG_5_14 ) : ( n16404 ) ;
assign n16406 =  ( n16215 ) ? ( VREG_5_15 ) : ( n16405 ) ;
assign n16407 =  ( n16214 ) ? ( VREG_6_0 ) : ( n16406 ) ;
assign n16408 =  ( n16213 ) ? ( VREG_6_1 ) : ( n16407 ) ;
assign n16409 =  ( n16212 ) ? ( VREG_6_2 ) : ( n16408 ) ;
assign n16410 =  ( n16211 ) ? ( VREG_6_3 ) : ( n16409 ) ;
assign n16411 =  ( n16210 ) ? ( VREG_6_4 ) : ( n16410 ) ;
assign n16412 =  ( n16209 ) ? ( VREG_6_5 ) : ( n16411 ) ;
assign n16413 =  ( n16208 ) ? ( VREG_6_6 ) : ( n16412 ) ;
assign n16414 =  ( n16207 ) ? ( VREG_6_7 ) : ( n16413 ) ;
assign n16415 =  ( n16206 ) ? ( VREG_6_8 ) : ( n16414 ) ;
assign n16416 =  ( n16205 ) ? ( VREG_6_9 ) : ( n16415 ) ;
assign n16417 =  ( n16204 ) ? ( VREG_6_10 ) : ( n16416 ) ;
assign n16418 =  ( n16203 ) ? ( VREG_6_11 ) : ( n16417 ) ;
assign n16419 =  ( n16202 ) ? ( VREG_6_12 ) : ( n16418 ) ;
assign n16420 =  ( n16201 ) ? ( VREG_6_13 ) : ( n16419 ) ;
assign n16421 =  ( n16200 ) ? ( VREG_6_14 ) : ( n16420 ) ;
assign n16422 =  ( n16199 ) ? ( VREG_6_15 ) : ( n16421 ) ;
assign n16423 =  ( n16198 ) ? ( VREG_7_0 ) : ( n16422 ) ;
assign n16424 =  ( n16197 ) ? ( VREG_7_1 ) : ( n16423 ) ;
assign n16425 =  ( n16196 ) ? ( VREG_7_2 ) : ( n16424 ) ;
assign n16426 =  ( n16195 ) ? ( VREG_7_3 ) : ( n16425 ) ;
assign n16427 =  ( n16194 ) ? ( VREG_7_4 ) : ( n16426 ) ;
assign n16428 =  ( n16193 ) ? ( VREG_7_5 ) : ( n16427 ) ;
assign n16429 =  ( n16192 ) ? ( VREG_7_6 ) : ( n16428 ) ;
assign n16430 =  ( n16191 ) ? ( VREG_7_7 ) : ( n16429 ) ;
assign n16431 =  ( n16190 ) ? ( VREG_7_8 ) : ( n16430 ) ;
assign n16432 =  ( n16189 ) ? ( VREG_7_9 ) : ( n16431 ) ;
assign n16433 =  ( n16188 ) ? ( VREG_7_10 ) : ( n16432 ) ;
assign n16434 =  ( n16187 ) ? ( VREG_7_11 ) : ( n16433 ) ;
assign n16435 =  ( n16186 ) ? ( VREG_7_12 ) : ( n16434 ) ;
assign n16436 =  ( n16185 ) ? ( VREG_7_13 ) : ( n16435 ) ;
assign n16437 =  ( n16184 ) ? ( VREG_7_14 ) : ( n16436 ) ;
assign n16438 =  ( n16183 ) ? ( VREG_7_15 ) : ( n16437 ) ;
assign n16439 =  ( n16182 ) ? ( VREG_8_0 ) : ( n16438 ) ;
assign n16440 =  ( n16181 ) ? ( VREG_8_1 ) : ( n16439 ) ;
assign n16441 =  ( n16180 ) ? ( VREG_8_2 ) : ( n16440 ) ;
assign n16442 =  ( n16179 ) ? ( VREG_8_3 ) : ( n16441 ) ;
assign n16443 =  ( n16178 ) ? ( VREG_8_4 ) : ( n16442 ) ;
assign n16444 =  ( n16177 ) ? ( VREG_8_5 ) : ( n16443 ) ;
assign n16445 =  ( n16176 ) ? ( VREG_8_6 ) : ( n16444 ) ;
assign n16446 =  ( n16175 ) ? ( VREG_8_7 ) : ( n16445 ) ;
assign n16447 =  ( n16174 ) ? ( VREG_8_8 ) : ( n16446 ) ;
assign n16448 =  ( n16173 ) ? ( VREG_8_9 ) : ( n16447 ) ;
assign n16449 =  ( n16172 ) ? ( VREG_8_10 ) : ( n16448 ) ;
assign n16450 =  ( n16171 ) ? ( VREG_8_11 ) : ( n16449 ) ;
assign n16451 =  ( n16170 ) ? ( VREG_8_12 ) : ( n16450 ) ;
assign n16452 =  ( n16169 ) ? ( VREG_8_13 ) : ( n16451 ) ;
assign n16453 =  ( n16168 ) ? ( VREG_8_14 ) : ( n16452 ) ;
assign n16454 =  ( n16167 ) ? ( VREG_8_15 ) : ( n16453 ) ;
assign n16455 =  ( n16166 ) ? ( VREG_9_0 ) : ( n16454 ) ;
assign n16456 =  ( n16165 ) ? ( VREG_9_1 ) : ( n16455 ) ;
assign n16457 =  ( n16164 ) ? ( VREG_9_2 ) : ( n16456 ) ;
assign n16458 =  ( n16163 ) ? ( VREG_9_3 ) : ( n16457 ) ;
assign n16459 =  ( n16162 ) ? ( VREG_9_4 ) : ( n16458 ) ;
assign n16460 =  ( n16161 ) ? ( VREG_9_5 ) : ( n16459 ) ;
assign n16461 =  ( n16160 ) ? ( VREG_9_6 ) : ( n16460 ) ;
assign n16462 =  ( n16159 ) ? ( VREG_9_7 ) : ( n16461 ) ;
assign n16463 =  ( n16158 ) ? ( VREG_9_8 ) : ( n16462 ) ;
assign n16464 =  ( n16157 ) ? ( VREG_9_9 ) : ( n16463 ) ;
assign n16465 =  ( n16156 ) ? ( VREG_9_10 ) : ( n16464 ) ;
assign n16466 =  ( n16155 ) ? ( VREG_9_11 ) : ( n16465 ) ;
assign n16467 =  ( n16154 ) ? ( VREG_9_12 ) : ( n16466 ) ;
assign n16468 =  ( n16153 ) ? ( VREG_9_13 ) : ( n16467 ) ;
assign n16469 =  ( n16152 ) ? ( VREG_9_14 ) : ( n16468 ) ;
assign n16470 =  ( n16151 ) ? ( VREG_9_15 ) : ( n16469 ) ;
assign n16471 =  ( n16150 ) ? ( VREG_10_0 ) : ( n16470 ) ;
assign n16472 =  ( n16149 ) ? ( VREG_10_1 ) : ( n16471 ) ;
assign n16473 =  ( n16148 ) ? ( VREG_10_2 ) : ( n16472 ) ;
assign n16474 =  ( n16147 ) ? ( VREG_10_3 ) : ( n16473 ) ;
assign n16475 =  ( n16146 ) ? ( VREG_10_4 ) : ( n16474 ) ;
assign n16476 =  ( n16145 ) ? ( VREG_10_5 ) : ( n16475 ) ;
assign n16477 =  ( n16144 ) ? ( VREG_10_6 ) : ( n16476 ) ;
assign n16478 =  ( n16143 ) ? ( VREG_10_7 ) : ( n16477 ) ;
assign n16479 =  ( n16142 ) ? ( VREG_10_8 ) : ( n16478 ) ;
assign n16480 =  ( n16141 ) ? ( VREG_10_9 ) : ( n16479 ) ;
assign n16481 =  ( n16140 ) ? ( VREG_10_10 ) : ( n16480 ) ;
assign n16482 =  ( n16139 ) ? ( VREG_10_11 ) : ( n16481 ) ;
assign n16483 =  ( n16138 ) ? ( VREG_10_12 ) : ( n16482 ) ;
assign n16484 =  ( n16137 ) ? ( VREG_10_13 ) : ( n16483 ) ;
assign n16485 =  ( n16136 ) ? ( VREG_10_14 ) : ( n16484 ) ;
assign n16486 =  ( n16135 ) ? ( VREG_10_15 ) : ( n16485 ) ;
assign n16487 =  ( n16134 ) ? ( VREG_11_0 ) : ( n16486 ) ;
assign n16488 =  ( n16133 ) ? ( VREG_11_1 ) : ( n16487 ) ;
assign n16489 =  ( n16132 ) ? ( VREG_11_2 ) : ( n16488 ) ;
assign n16490 =  ( n16131 ) ? ( VREG_11_3 ) : ( n16489 ) ;
assign n16491 =  ( n16130 ) ? ( VREG_11_4 ) : ( n16490 ) ;
assign n16492 =  ( n16129 ) ? ( VREG_11_5 ) : ( n16491 ) ;
assign n16493 =  ( n16128 ) ? ( VREG_11_6 ) : ( n16492 ) ;
assign n16494 =  ( n16127 ) ? ( VREG_11_7 ) : ( n16493 ) ;
assign n16495 =  ( n16126 ) ? ( VREG_11_8 ) : ( n16494 ) ;
assign n16496 =  ( n16125 ) ? ( VREG_11_9 ) : ( n16495 ) ;
assign n16497 =  ( n16124 ) ? ( VREG_11_10 ) : ( n16496 ) ;
assign n16498 =  ( n16123 ) ? ( VREG_11_11 ) : ( n16497 ) ;
assign n16499 =  ( n16122 ) ? ( VREG_11_12 ) : ( n16498 ) ;
assign n16500 =  ( n16121 ) ? ( VREG_11_13 ) : ( n16499 ) ;
assign n16501 =  ( n16120 ) ? ( VREG_11_14 ) : ( n16500 ) ;
assign n16502 =  ( n16119 ) ? ( VREG_11_15 ) : ( n16501 ) ;
assign n16503 =  ( n16118 ) ? ( VREG_12_0 ) : ( n16502 ) ;
assign n16504 =  ( n16117 ) ? ( VREG_12_1 ) : ( n16503 ) ;
assign n16505 =  ( n16116 ) ? ( VREG_12_2 ) : ( n16504 ) ;
assign n16506 =  ( n16115 ) ? ( VREG_12_3 ) : ( n16505 ) ;
assign n16507 =  ( n16114 ) ? ( VREG_12_4 ) : ( n16506 ) ;
assign n16508 =  ( n16113 ) ? ( VREG_12_5 ) : ( n16507 ) ;
assign n16509 =  ( n16112 ) ? ( VREG_12_6 ) : ( n16508 ) ;
assign n16510 =  ( n16111 ) ? ( VREG_12_7 ) : ( n16509 ) ;
assign n16511 =  ( n16110 ) ? ( VREG_12_8 ) : ( n16510 ) ;
assign n16512 =  ( n16109 ) ? ( VREG_12_9 ) : ( n16511 ) ;
assign n16513 =  ( n16108 ) ? ( VREG_12_10 ) : ( n16512 ) ;
assign n16514 =  ( n16107 ) ? ( VREG_12_11 ) : ( n16513 ) ;
assign n16515 =  ( n16106 ) ? ( VREG_12_12 ) : ( n16514 ) ;
assign n16516 =  ( n16105 ) ? ( VREG_12_13 ) : ( n16515 ) ;
assign n16517 =  ( n16104 ) ? ( VREG_12_14 ) : ( n16516 ) ;
assign n16518 =  ( n16103 ) ? ( VREG_12_15 ) : ( n16517 ) ;
assign n16519 =  ( n16102 ) ? ( VREG_13_0 ) : ( n16518 ) ;
assign n16520 =  ( n16101 ) ? ( VREG_13_1 ) : ( n16519 ) ;
assign n16521 =  ( n16100 ) ? ( VREG_13_2 ) : ( n16520 ) ;
assign n16522 =  ( n16099 ) ? ( VREG_13_3 ) : ( n16521 ) ;
assign n16523 =  ( n16098 ) ? ( VREG_13_4 ) : ( n16522 ) ;
assign n16524 =  ( n16097 ) ? ( VREG_13_5 ) : ( n16523 ) ;
assign n16525 =  ( n16096 ) ? ( VREG_13_6 ) : ( n16524 ) ;
assign n16526 =  ( n16095 ) ? ( VREG_13_7 ) : ( n16525 ) ;
assign n16527 =  ( n16094 ) ? ( VREG_13_8 ) : ( n16526 ) ;
assign n16528 =  ( n16093 ) ? ( VREG_13_9 ) : ( n16527 ) ;
assign n16529 =  ( n16092 ) ? ( VREG_13_10 ) : ( n16528 ) ;
assign n16530 =  ( n16091 ) ? ( VREG_13_11 ) : ( n16529 ) ;
assign n16531 =  ( n16090 ) ? ( VREG_13_12 ) : ( n16530 ) ;
assign n16532 =  ( n16089 ) ? ( VREG_13_13 ) : ( n16531 ) ;
assign n16533 =  ( n16088 ) ? ( VREG_13_14 ) : ( n16532 ) ;
assign n16534 =  ( n16087 ) ? ( VREG_13_15 ) : ( n16533 ) ;
assign n16535 =  ( n16086 ) ? ( VREG_14_0 ) : ( n16534 ) ;
assign n16536 =  ( n16085 ) ? ( VREG_14_1 ) : ( n16535 ) ;
assign n16537 =  ( n16084 ) ? ( VREG_14_2 ) : ( n16536 ) ;
assign n16538 =  ( n16083 ) ? ( VREG_14_3 ) : ( n16537 ) ;
assign n16539 =  ( n16082 ) ? ( VREG_14_4 ) : ( n16538 ) ;
assign n16540 =  ( n16081 ) ? ( VREG_14_5 ) : ( n16539 ) ;
assign n16541 =  ( n16080 ) ? ( VREG_14_6 ) : ( n16540 ) ;
assign n16542 =  ( n16079 ) ? ( VREG_14_7 ) : ( n16541 ) ;
assign n16543 =  ( n16078 ) ? ( VREG_14_8 ) : ( n16542 ) ;
assign n16544 =  ( n16077 ) ? ( VREG_14_9 ) : ( n16543 ) ;
assign n16545 =  ( n16076 ) ? ( VREG_14_10 ) : ( n16544 ) ;
assign n16546 =  ( n16075 ) ? ( VREG_14_11 ) : ( n16545 ) ;
assign n16547 =  ( n16074 ) ? ( VREG_14_12 ) : ( n16546 ) ;
assign n16548 =  ( n16073 ) ? ( VREG_14_13 ) : ( n16547 ) ;
assign n16549 =  ( n16072 ) ? ( VREG_14_14 ) : ( n16548 ) ;
assign n16550 =  ( n16071 ) ? ( VREG_14_15 ) : ( n16549 ) ;
assign n16551 =  ( n16070 ) ? ( VREG_15_0 ) : ( n16550 ) ;
assign n16552 =  ( n16069 ) ? ( VREG_15_1 ) : ( n16551 ) ;
assign n16553 =  ( n16068 ) ? ( VREG_15_2 ) : ( n16552 ) ;
assign n16554 =  ( n16067 ) ? ( VREG_15_3 ) : ( n16553 ) ;
assign n16555 =  ( n16066 ) ? ( VREG_15_4 ) : ( n16554 ) ;
assign n16556 =  ( n16065 ) ? ( VREG_15_5 ) : ( n16555 ) ;
assign n16557 =  ( n16064 ) ? ( VREG_15_6 ) : ( n16556 ) ;
assign n16558 =  ( n16063 ) ? ( VREG_15_7 ) : ( n16557 ) ;
assign n16559 =  ( n16062 ) ? ( VREG_15_8 ) : ( n16558 ) ;
assign n16560 =  ( n16061 ) ? ( VREG_15_9 ) : ( n16559 ) ;
assign n16561 =  ( n16060 ) ? ( VREG_15_10 ) : ( n16560 ) ;
assign n16562 =  ( n16059 ) ? ( VREG_15_11 ) : ( n16561 ) ;
assign n16563 =  ( n16058 ) ? ( VREG_15_12 ) : ( n16562 ) ;
assign n16564 =  ( n16057 ) ? ( VREG_15_13 ) : ( n16563 ) ;
assign n16565 =  ( n16056 ) ? ( VREG_15_14 ) : ( n16564 ) ;
assign n16566 =  ( n16055 ) ? ( VREG_15_15 ) : ( n16565 ) ;
assign n16567 =  ( n16054 ) ? ( VREG_16_0 ) : ( n16566 ) ;
assign n16568 =  ( n16053 ) ? ( VREG_16_1 ) : ( n16567 ) ;
assign n16569 =  ( n16052 ) ? ( VREG_16_2 ) : ( n16568 ) ;
assign n16570 =  ( n16051 ) ? ( VREG_16_3 ) : ( n16569 ) ;
assign n16571 =  ( n16050 ) ? ( VREG_16_4 ) : ( n16570 ) ;
assign n16572 =  ( n16049 ) ? ( VREG_16_5 ) : ( n16571 ) ;
assign n16573 =  ( n16048 ) ? ( VREG_16_6 ) : ( n16572 ) ;
assign n16574 =  ( n16047 ) ? ( VREG_16_7 ) : ( n16573 ) ;
assign n16575 =  ( n16046 ) ? ( VREG_16_8 ) : ( n16574 ) ;
assign n16576 =  ( n16045 ) ? ( VREG_16_9 ) : ( n16575 ) ;
assign n16577 =  ( n16044 ) ? ( VREG_16_10 ) : ( n16576 ) ;
assign n16578 =  ( n16043 ) ? ( VREG_16_11 ) : ( n16577 ) ;
assign n16579 =  ( n16042 ) ? ( VREG_16_12 ) : ( n16578 ) ;
assign n16580 =  ( n16041 ) ? ( VREG_16_13 ) : ( n16579 ) ;
assign n16581 =  ( n16040 ) ? ( VREG_16_14 ) : ( n16580 ) ;
assign n16582 =  ( n16039 ) ? ( VREG_16_15 ) : ( n16581 ) ;
assign n16583 =  ( n16038 ) ? ( VREG_17_0 ) : ( n16582 ) ;
assign n16584 =  ( n16037 ) ? ( VREG_17_1 ) : ( n16583 ) ;
assign n16585 =  ( n16036 ) ? ( VREG_17_2 ) : ( n16584 ) ;
assign n16586 =  ( n16035 ) ? ( VREG_17_3 ) : ( n16585 ) ;
assign n16587 =  ( n16034 ) ? ( VREG_17_4 ) : ( n16586 ) ;
assign n16588 =  ( n16033 ) ? ( VREG_17_5 ) : ( n16587 ) ;
assign n16589 =  ( n16032 ) ? ( VREG_17_6 ) : ( n16588 ) ;
assign n16590 =  ( n16031 ) ? ( VREG_17_7 ) : ( n16589 ) ;
assign n16591 =  ( n16030 ) ? ( VREG_17_8 ) : ( n16590 ) ;
assign n16592 =  ( n16029 ) ? ( VREG_17_9 ) : ( n16591 ) ;
assign n16593 =  ( n16028 ) ? ( VREG_17_10 ) : ( n16592 ) ;
assign n16594 =  ( n16027 ) ? ( VREG_17_11 ) : ( n16593 ) ;
assign n16595 =  ( n16026 ) ? ( VREG_17_12 ) : ( n16594 ) ;
assign n16596 =  ( n16025 ) ? ( VREG_17_13 ) : ( n16595 ) ;
assign n16597 =  ( n16024 ) ? ( VREG_17_14 ) : ( n16596 ) ;
assign n16598 =  ( n16023 ) ? ( VREG_17_15 ) : ( n16597 ) ;
assign n16599 =  ( n16022 ) ? ( VREG_18_0 ) : ( n16598 ) ;
assign n16600 =  ( n16021 ) ? ( VREG_18_1 ) : ( n16599 ) ;
assign n16601 =  ( n16020 ) ? ( VREG_18_2 ) : ( n16600 ) ;
assign n16602 =  ( n16019 ) ? ( VREG_18_3 ) : ( n16601 ) ;
assign n16603 =  ( n16018 ) ? ( VREG_18_4 ) : ( n16602 ) ;
assign n16604 =  ( n16017 ) ? ( VREG_18_5 ) : ( n16603 ) ;
assign n16605 =  ( n16016 ) ? ( VREG_18_6 ) : ( n16604 ) ;
assign n16606 =  ( n16015 ) ? ( VREG_18_7 ) : ( n16605 ) ;
assign n16607 =  ( n16014 ) ? ( VREG_18_8 ) : ( n16606 ) ;
assign n16608 =  ( n16013 ) ? ( VREG_18_9 ) : ( n16607 ) ;
assign n16609 =  ( n16012 ) ? ( VREG_18_10 ) : ( n16608 ) ;
assign n16610 =  ( n16011 ) ? ( VREG_18_11 ) : ( n16609 ) ;
assign n16611 =  ( n16010 ) ? ( VREG_18_12 ) : ( n16610 ) ;
assign n16612 =  ( n16009 ) ? ( VREG_18_13 ) : ( n16611 ) ;
assign n16613 =  ( n16008 ) ? ( VREG_18_14 ) : ( n16612 ) ;
assign n16614 =  ( n16007 ) ? ( VREG_18_15 ) : ( n16613 ) ;
assign n16615 =  ( n16006 ) ? ( VREG_19_0 ) : ( n16614 ) ;
assign n16616 =  ( n16005 ) ? ( VREG_19_1 ) : ( n16615 ) ;
assign n16617 =  ( n16004 ) ? ( VREG_19_2 ) : ( n16616 ) ;
assign n16618 =  ( n16003 ) ? ( VREG_19_3 ) : ( n16617 ) ;
assign n16619 =  ( n16002 ) ? ( VREG_19_4 ) : ( n16618 ) ;
assign n16620 =  ( n16001 ) ? ( VREG_19_5 ) : ( n16619 ) ;
assign n16621 =  ( n16000 ) ? ( VREG_19_6 ) : ( n16620 ) ;
assign n16622 =  ( n15999 ) ? ( VREG_19_7 ) : ( n16621 ) ;
assign n16623 =  ( n15998 ) ? ( VREG_19_8 ) : ( n16622 ) ;
assign n16624 =  ( n15997 ) ? ( VREG_19_9 ) : ( n16623 ) ;
assign n16625 =  ( n15996 ) ? ( VREG_19_10 ) : ( n16624 ) ;
assign n16626 =  ( n15995 ) ? ( VREG_19_11 ) : ( n16625 ) ;
assign n16627 =  ( n15994 ) ? ( VREG_19_12 ) : ( n16626 ) ;
assign n16628 =  ( n15993 ) ? ( VREG_19_13 ) : ( n16627 ) ;
assign n16629 =  ( n15992 ) ? ( VREG_19_14 ) : ( n16628 ) ;
assign n16630 =  ( n15991 ) ? ( VREG_19_15 ) : ( n16629 ) ;
assign n16631 =  ( n15990 ) ? ( VREG_20_0 ) : ( n16630 ) ;
assign n16632 =  ( n15989 ) ? ( VREG_20_1 ) : ( n16631 ) ;
assign n16633 =  ( n15988 ) ? ( VREG_20_2 ) : ( n16632 ) ;
assign n16634 =  ( n15987 ) ? ( VREG_20_3 ) : ( n16633 ) ;
assign n16635 =  ( n15986 ) ? ( VREG_20_4 ) : ( n16634 ) ;
assign n16636 =  ( n15985 ) ? ( VREG_20_5 ) : ( n16635 ) ;
assign n16637 =  ( n15984 ) ? ( VREG_20_6 ) : ( n16636 ) ;
assign n16638 =  ( n15983 ) ? ( VREG_20_7 ) : ( n16637 ) ;
assign n16639 =  ( n15982 ) ? ( VREG_20_8 ) : ( n16638 ) ;
assign n16640 =  ( n15981 ) ? ( VREG_20_9 ) : ( n16639 ) ;
assign n16641 =  ( n15980 ) ? ( VREG_20_10 ) : ( n16640 ) ;
assign n16642 =  ( n15979 ) ? ( VREG_20_11 ) : ( n16641 ) ;
assign n16643 =  ( n15978 ) ? ( VREG_20_12 ) : ( n16642 ) ;
assign n16644 =  ( n15977 ) ? ( VREG_20_13 ) : ( n16643 ) ;
assign n16645 =  ( n15976 ) ? ( VREG_20_14 ) : ( n16644 ) ;
assign n16646 =  ( n15975 ) ? ( VREG_20_15 ) : ( n16645 ) ;
assign n16647 =  ( n15974 ) ? ( VREG_21_0 ) : ( n16646 ) ;
assign n16648 =  ( n15973 ) ? ( VREG_21_1 ) : ( n16647 ) ;
assign n16649 =  ( n15972 ) ? ( VREG_21_2 ) : ( n16648 ) ;
assign n16650 =  ( n15971 ) ? ( VREG_21_3 ) : ( n16649 ) ;
assign n16651 =  ( n15970 ) ? ( VREG_21_4 ) : ( n16650 ) ;
assign n16652 =  ( n15969 ) ? ( VREG_21_5 ) : ( n16651 ) ;
assign n16653 =  ( n15968 ) ? ( VREG_21_6 ) : ( n16652 ) ;
assign n16654 =  ( n15967 ) ? ( VREG_21_7 ) : ( n16653 ) ;
assign n16655 =  ( n15966 ) ? ( VREG_21_8 ) : ( n16654 ) ;
assign n16656 =  ( n15965 ) ? ( VREG_21_9 ) : ( n16655 ) ;
assign n16657 =  ( n15964 ) ? ( VREG_21_10 ) : ( n16656 ) ;
assign n16658 =  ( n15963 ) ? ( VREG_21_11 ) : ( n16657 ) ;
assign n16659 =  ( n15962 ) ? ( VREG_21_12 ) : ( n16658 ) ;
assign n16660 =  ( n15961 ) ? ( VREG_21_13 ) : ( n16659 ) ;
assign n16661 =  ( n15960 ) ? ( VREG_21_14 ) : ( n16660 ) ;
assign n16662 =  ( n15959 ) ? ( VREG_21_15 ) : ( n16661 ) ;
assign n16663 =  ( n15958 ) ? ( VREG_22_0 ) : ( n16662 ) ;
assign n16664 =  ( n15957 ) ? ( VREG_22_1 ) : ( n16663 ) ;
assign n16665 =  ( n15956 ) ? ( VREG_22_2 ) : ( n16664 ) ;
assign n16666 =  ( n15955 ) ? ( VREG_22_3 ) : ( n16665 ) ;
assign n16667 =  ( n15954 ) ? ( VREG_22_4 ) : ( n16666 ) ;
assign n16668 =  ( n15953 ) ? ( VREG_22_5 ) : ( n16667 ) ;
assign n16669 =  ( n15952 ) ? ( VREG_22_6 ) : ( n16668 ) ;
assign n16670 =  ( n15951 ) ? ( VREG_22_7 ) : ( n16669 ) ;
assign n16671 =  ( n15950 ) ? ( VREG_22_8 ) : ( n16670 ) ;
assign n16672 =  ( n15949 ) ? ( VREG_22_9 ) : ( n16671 ) ;
assign n16673 =  ( n15948 ) ? ( VREG_22_10 ) : ( n16672 ) ;
assign n16674 =  ( n15947 ) ? ( VREG_22_11 ) : ( n16673 ) ;
assign n16675 =  ( n15946 ) ? ( VREG_22_12 ) : ( n16674 ) ;
assign n16676 =  ( n15945 ) ? ( VREG_22_13 ) : ( n16675 ) ;
assign n16677 =  ( n15944 ) ? ( VREG_22_14 ) : ( n16676 ) ;
assign n16678 =  ( n15943 ) ? ( VREG_22_15 ) : ( n16677 ) ;
assign n16679 =  ( n15942 ) ? ( VREG_23_0 ) : ( n16678 ) ;
assign n16680 =  ( n15941 ) ? ( VREG_23_1 ) : ( n16679 ) ;
assign n16681 =  ( n15940 ) ? ( VREG_23_2 ) : ( n16680 ) ;
assign n16682 =  ( n15939 ) ? ( VREG_23_3 ) : ( n16681 ) ;
assign n16683 =  ( n15938 ) ? ( VREG_23_4 ) : ( n16682 ) ;
assign n16684 =  ( n15937 ) ? ( VREG_23_5 ) : ( n16683 ) ;
assign n16685 =  ( n15936 ) ? ( VREG_23_6 ) : ( n16684 ) ;
assign n16686 =  ( n15935 ) ? ( VREG_23_7 ) : ( n16685 ) ;
assign n16687 =  ( n15934 ) ? ( VREG_23_8 ) : ( n16686 ) ;
assign n16688 =  ( n15933 ) ? ( VREG_23_9 ) : ( n16687 ) ;
assign n16689 =  ( n15932 ) ? ( VREG_23_10 ) : ( n16688 ) ;
assign n16690 =  ( n15931 ) ? ( VREG_23_11 ) : ( n16689 ) ;
assign n16691 =  ( n15930 ) ? ( VREG_23_12 ) : ( n16690 ) ;
assign n16692 =  ( n15929 ) ? ( VREG_23_13 ) : ( n16691 ) ;
assign n16693 =  ( n15928 ) ? ( VREG_23_14 ) : ( n16692 ) ;
assign n16694 =  ( n15927 ) ? ( VREG_23_15 ) : ( n16693 ) ;
assign n16695 =  ( n15926 ) ? ( VREG_24_0 ) : ( n16694 ) ;
assign n16696 =  ( n15925 ) ? ( VREG_24_1 ) : ( n16695 ) ;
assign n16697 =  ( n15924 ) ? ( VREG_24_2 ) : ( n16696 ) ;
assign n16698 =  ( n15923 ) ? ( VREG_24_3 ) : ( n16697 ) ;
assign n16699 =  ( n15922 ) ? ( VREG_24_4 ) : ( n16698 ) ;
assign n16700 =  ( n15921 ) ? ( VREG_24_5 ) : ( n16699 ) ;
assign n16701 =  ( n15920 ) ? ( VREG_24_6 ) : ( n16700 ) ;
assign n16702 =  ( n15919 ) ? ( VREG_24_7 ) : ( n16701 ) ;
assign n16703 =  ( n15918 ) ? ( VREG_24_8 ) : ( n16702 ) ;
assign n16704 =  ( n15917 ) ? ( VREG_24_9 ) : ( n16703 ) ;
assign n16705 =  ( n15916 ) ? ( VREG_24_10 ) : ( n16704 ) ;
assign n16706 =  ( n15915 ) ? ( VREG_24_11 ) : ( n16705 ) ;
assign n16707 =  ( n15914 ) ? ( VREG_24_12 ) : ( n16706 ) ;
assign n16708 =  ( n15913 ) ? ( VREG_24_13 ) : ( n16707 ) ;
assign n16709 =  ( n15912 ) ? ( VREG_24_14 ) : ( n16708 ) ;
assign n16710 =  ( n15911 ) ? ( VREG_24_15 ) : ( n16709 ) ;
assign n16711 =  ( n15910 ) ? ( VREG_25_0 ) : ( n16710 ) ;
assign n16712 =  ( n15909 ) ? ( VREG_25_1 ) : ( n16711 ) ;
assign n16713 =  ( n15908 ) ? ( VREG_25_2 ) : ( n16712 ) ;
assign n16714 =  ( n15907 ) ? ( VREG_25_3 ) : ( n16713 ) ;
assign n16715 =  ( n15906 ) ? ( VREG_25_4 ) : ( n16714 ) ;
assign n16716 =  ( n15905 ) ? ( VREG_25_5 ) : ( n16715 ) ;
assign n16717 =  ( n15904 ) ? ( VREG_25_6 ) : ( n16716 ) ;
assign n16718 =  ( n15903 ) ? ( VREG_25_7 ) : ( n16717 ) ;
assign n16719 =  ( n15902 ) ? ( VREG_25_8 ) : ( n16718 ) ;
assign n16720 =  ( n15901 ) ? ( VREG_25_9 ) : ( n16719 ) ;
assign n16721 =  ( n15900 ) ? ( VREG_25_10 ) : ( n16720 ) ;
assign n16722 =  ( n15899 ) ? ( VREG_25_11 ) : ( n16721 ) ;
assign n16723 =  ( n15898 ) ? ( VREG_25_12 ) : ( n16722 ) ;
assign n16724 =  ( n15897 ) ? ( VREG_25_13 ) : ( n16723 ) ;
assign n16725 =  ( n15896 ) ? ( VREG_25_14 ) : ( n16724 ) ;
assign n16726 =  ( n15895 ) ? ( VREG_25_15 ) : ( n16725 ) ;
assign n16727 =  ( n15894 ) ? ( VREG_26_0 ) : ( n16726 ) ;
assign n16728 =  ( n15893 ) ? ( VREG_26_1 ) : ( n16727 ) ;
assign n16729 =  ( n15892 ) ? ( VREG_26_2 ) : ( n16728 ) ;
assign n16730 =  ( n15891 ) ? ( VREG_26_3 ) : ( n16729 ) ;
assign n16731 =  ( n15890 ) ? ( VREG_26_4 ) : ( n16730 ) ;
assign n16732 =  ( n15889 ) ? ( VREG_26_5 ) : ( n16731 ) ;
assign n16733 =  ( n15888 ) ? ( VREG_26_6 ) : ( n16732 ) ;
assign n16734 =  ( n15887 ) ? ( VREG_26_7 ) : ( n16733 ) ;
assign n16735 =  ( n15886 ) ? ( VREG_26_8 ) : ( n16734 ) ;
assign n16736 =  ( n15885 ) ? ( VREG_26_9 ) : ( n16735 ) ;
assign n16737 =  ( n15884 ) ? ( VREG_26_10 ) : ( n16736 ) ;
assign n16738 =  ( n15883 ) ? ( VREG_26_11 ) : ( n16737 ) ;
assign n16739 =  ( n15882 ) ? ( VREG_26_12 ) : ( n16738 ) ;
assign n16740 =  ( n15881 ) ? ( VREG_26_13 ) : ( n16739 ) ;
assign n16741 =  ( n15880 ) ? ( VREG_26_14 ) : ( n16740 ) ;
assign n16742 =  ( n15879 ) ? ( VREG_26_15 ) : ( n16741 ) ;
assign n16743 =  ( n15878 ) ? ( VREG_27_0 ) : ( n16742 ) ;
assign n16744 =  ( n15877 ) ? ( VREG_27_1 ) : ( n16743 ) ;
assign n16745 =  ( n15876 ) ? ( VREG_27_2 ) : ( n16744 ) ;
assign n16746 =  ( n15875 ) ? ( VREG_27_3 ) : ( n16745 ) ;
assign n16747 =  ( n15874 ) ? ( VREG_27_4 ) : ( n16746 ) ;
assign n16748 =  ( n15873 ) ? ( VREG_27_5 ) : ( n16747 ) ;
assign n16749 =  ( n15872 ) ? ( VREG_27_6 ) : ( n16748 ) ;
assign n16750 =  ( n15871 ) ? ( VREG_27_7 ) : ( n16749 ) ;
assign n16751 =  ( n15870 ) ? ( VREG_27_8 ) : ( n16750 ) ;
assign n16752 =  ( n15869 ) ? ( VREG_27_9 ) : ( n16751 ) ;
assign n16753 =  ( n15868 ) ? ( VREG_27_10 ) : ( n16752 ) ;
assign n16754 =  ( n15867 ) ? ( VREG_27_11 ) : ( n16753 ) ;
assign n16755 =  ( n15866 ) ? ( VREG_27_12 ) : ( n16754 ) ;
assign n16756 =  ( n15865 ) ? ( VREG_27_13 ) : ( n16755 ) ;
assign n16757 =  ( n15864 ) ? ( VREG_27_14 ) : ( n16756 ) ;
assign n16758 =  ( n15863 ) ? ( VREG_27_15 ) : ( n16757 ) ;
assign n16759 =  ( n15862 ) ? ( VREG_28_0 ) : ( n16758 ) ;
assign n16760 =  ( n15861 ) ? ( VREG_28_1 ) : ( n16759 ) ;
assign n16761 =  ( n15860 ) ? ( VREG_28_2 ) : ( n16760 ) ;
assign n16762 =  ( n15859 ) ? ( VREG_28_3 ) : ( n16761 ) ;
assign n16763 =  ( n15858 ) ? ( VREG_28_4 ) : ( n16762 ) ;
assign n16764 =  ( n15857 ) ? ( VREG_28_5 ) : ( n16763 ) ;
assign n16765 =  ( n15856 ) ? ( VREG_28_6 ) : ( n16764 ) ;
assign n16766 =  ( n15855 ) ? ( VREG_28_7 ) : ( n16765 ) ;
assign n16767 =  ( n15854 ) ? ( VREG_28_8 ) : ( n16766 ) ;
assign n16768 =  ( n15853 ) ? ( VREG_28_9 ) : ( n16767 ) ;
assign n16769 =  ( n15852 ) ? ( VREG_28_10 ) : ( n16768 ) ;
assign n16770 =  ( n15851 ) ? ( VREG_28_11 ) : ( n16769 ) ;
assign n16771 =  ( n15850 ) ? ( VREG_28_12 ) : ( n16770 ) ;
assign n16772 =  ( n15849 ) ? ( VREG_28_13 ) : ( n16771 ) ;
assign n16773 =  ( n15848 ) ? ( VREG_28_14 ) : ( n16772 ) ;
assign n16774 =  ( n15847 ) ? ( VREG_28_15 ) : ( n16773 ) ;
assign n16775 =  ( n15846 ) ? ( VREG_29_0 ) : ( n16774 ) ;
assign n16776 =  ( n15845 ) ? ( VREG_29_1 ) : ( n16775 ) ;
assign n16777 =  ( n15844 ) ? ( VREG_29_2 ) : ( n16776 ) ;
assign n16778 =  ( n15843 ) ? ( VREG_29_3 ) : ( n16777 ) ;
assign n16779 =  ( n15842 ) ? ( VREG_29_4 ) : ( n16778 ) ;
assign n16780 =  ( n15841 ) ? ( VREG_29_5 ) : ( n16779 ) ;
assign n16781 =  ( n15840 ) ? ( VREG_29_6 ) : ( n16780 ) ;
assign n16782 =  ( n15839 ) ? ( VREG_29_7 ) : ( n16781 ) ;
assign n16783 =  ( n15838 ) ? ( VREG_29_8 ) : ( n16782 ) ;
assign n16784 =  ( n15837 ) ? ( VREG_29_9 ) : ( n16783 ) ;
assign n16785 =  ( n15836 ) ? ( VREG_29_10 ) : ( n16784 ) ;
assign n16786 =  ( n15835 ) ? ( VREG_29_11 ) : ( n16785 ) ;
assign n16787 =  ( n15834 ) ? ( VREG_29_12 ) : ( n16786 ) ;
assign n16788 =  ( n15833 ) ? ( VREG_29_13 ) : ( n16787 ) ;
assign n16789 =  ( n15832 ) ? ( VREG_29_14 ) : ( n16788 ) ;
assign n16790 =  ( n15831 ) ? ( VREG_29_15 ) : ( n16789 ) ;
assign n16791 =  ( n15830 ) ? ( VREG_30_0 ) : ( n16790 ) ;
assign n16792 =  ( n15829 ) ? ( VREG_30_1 ) : ( n16791 ) ;
assign n16793 =  ( n15828 ) ? ( VREG_30_2 ) : ( n16792 ) ;
assign n16794 =  ( n15827 ) ? ( VREG_30_3 ) : ( n16793 ) ;
assign n16795 =  ( n15826 ) ? ( VREG_30_4 ) : ( n16794 ) ;
assign n16796 =  ( n15825 ) ? ( VREG_30_5 ) : ( n16795 ) ;
assign n16797 =  ( n15824 ) ? ( VREG_30_6 ) : ( n16796 ) ;
assign n16798 =  ( n15823 ) ? ( VREG_30_7 ) : ( n16797 ) ;
assign n16799 =  ( n15822 ) ? ( VREG_30_8 ) : ( n16798 ) ;
assign n16800 =  ( n15821 ) ? ( VREG_30_9 ) : ( n16799 ) ;
assign n16801 =  ( n15820 ) ? ( VREG_30_10 ) : ( n16800 ) ;
assign n16802 =  ( n15819 ) ? ( VREG_30_11 ) : ( n16801 ) ;
assign n16803 =  ( n15818 ) ? ( VREG_30_12 ) : ( n16802 ) ;
assign n16804 =  ( n15817 ) ? ( VREG_30_13 ) : ( n16803 ) ;
assign n16805 =  ( n15816 ) ? ( VREG_30_14 ) : ( n16804 ) ;
assign n16806 =  ( n15815 ) ? ( VREG_30_15 ) : ( n16805 ) ;
assign n16807 =  ( n15814 ) ? ( VREG_31_0 ) : ( n16806 ) ;
assign n16808 =  ( n15812 ) ? ( VREG_31_1 ) : ( n16807 ) ;
assign n16809 =  ( n15810 ) ? ( VREG_31_2 ) : ( n16808 ) ;
assign n16810 =  ( n15808 ) ? ( VREG_31_3 ) : ( n16809 ) ;
assign n16811 =  ( n15806 ) ? ( VREG_31_4 ) : ( n16810 ) ;
assign n16812 =  ( n15804 ) ? ( VREG_31_5 ) : ( n16811 ) ;
assign n16813 =  ( n15802 ) ? ( VREG_31_6 ) : ( n16812 ) ;
assign n16814 =  ( n15800 ) ? ( VREG_31_7 ) : ( n16813 ) ;
assign n16815 =  ( n15798 ) ? ( VREG_31_8 ) : ( n16814 ) ;
assign n16816 =  ( n15796 ) ? ( VREG_31_9 ) : ( n16815 ) ;
assign n16817 =  ( n15794 ) ? ( VREG_31_10 ) : ( n16816 ) ;
assign n16818 =  ( n15792 ) ? ( VREG_31_11 ) : ( n16817 ) ;
assign n16819 =  ( n15790 ) ? ( VREG_31_12 ) : ( n16818 ) ;
assign n16820 =  ( n15788 ) ? ( VREG_31_13 ) : ( n16819 ) ;
assign n16821 =  ( n15786 ) ? ( VREG_31_14 ) : ( n16820 ) ;
assign n16822 =  ( n15784 ) ? ( VREG_31_15 ) : ( n16821 ) ;
assign n16823 =  ( n16822 ) + ( n140 )  ;
assign n16824 =  ( n16822 ) - ( n140 )  ;
assign n16825 =  ( n16822 ) & ( n140 )  ;
assign n16826 =  ( n16822 ) | ( n140 )  ;
assign n16827 =  ( ( n16822 ) * ( n140 ))  ;
assign n16828 =  ( n148 ) ? ( n16827 ) : ( VREG_0_15 ) ;
assign n16829 =  ( n146 ) ? ( n16826 ) : ( n16828 ) ;
assign n16830 =  ( n144 ) ? ( n16825 ) : ( n16829 ) ;
assign n16831 =  ( n142 ) ? ( n16824 ) : ( n16830 ) ;
assign n16832 =  ( n10 ) ? ( n16823 ) : ( n16831 ) ;
assign n16833 =  ( n77 ) & ( n15783 )  ;
assign n16834 =  ( n77 ) & ( n15785 )  ;
assign n16835 =  ( n77 ) & ( n15787 )  ;
assign n16836 =  ( n77 ) & ( n15789 )  ;
assign n16837 =  ( n77 ) & ( n15791 )  ;
assign n16838 =  ( n77 ) & ( n15793 )  ;
assign n16839 =  ( n77 ) & ( n15795 )  ;
assign n16840 =  ( n77 ) & ( n15797 )  ;
assign n16841 =  ( n77 ) & ( n15799 )  ;
assign n16842 =  ( n77 ) & ( n15801 )  ;
assign n16843 =  ( n77 ) & ( n15803 )  ;
assign n16844 =  ( n77 ) & ( n15805 )  ;
assign n16845 =  ( n77 ) & ( n15807 )  ;
assign n16846 =  ( n77 ) & ( n15809 )  ;
assign n16847 =  ( n77 ) & ( n15811 )  ;
assign n16848 =  ( n77 ) & ( n15813 )  ;
assign n16849 =  ( n78 ) & ( n15783 )  ;
assign n16850 =  ( n78 ) & ( n15785 )  ;
assign n16851 =  ( n78 ) & ( n15787 )  ;
assign n16852 =  ( n78 ) & ( n15789 )  ;
assign n16853 =  ( n78 ) & ( n15791 )  ;
assign n16854 =  ( n78 ) & ( n15793 )  ;
assign n16855 =  ( n78 ) & ( n15795 )  ;
assign n16856 =  ( n78 ) & ( n15797 )  ;
assign n16857 =  ( n78 ) & ( n15799 )  ;
assign n16858 =  ( n78 ) & ( n15801 )  ;
assign n16859 =  ( n78 ) & ( n15803 )  ;
assign n16860 =  ( n78 ) & ( n15805 )  ;
assign n16861 =  ( n78 ) & ( n15807 )  ;
assign n16862 =  ( n78 ) & ( n15809 )  ;
assign n16863 =  ( n78 ) & ( n15811 )  ;
assign n16864 =  ( n78 ) & ( n15813 )  ;
assign n16865 =  ( n79 ) & ( n15783 )  ;
assign n16866 =  ( n79 ) & ( n15785 )  ;
assign n16867 =  ( n79 ) & ( n15787 )  ;
assign n16868 =  ( n79 ) & ( n15789 )  ;
assign n16869 =  ( n79 ) & ( n15791 )  ;
assign n16870 =  ( n79 ) & ( n15793 )  ;
assign n16871 =  ( n79 ) & ( n15795 )  ;
assign n16872 =  ( n79 ) & ( n15797 )  ;
assign n16873 =  ( n79 ) & ( n15799 )  ;
assign n16874 =  ( n79 ) & ( n15801 )  ;
assign n16875 =  ( n79 ) & ( n15803 )  ;
assign n16876 =  ( n79 ) & ( n15805 )  ;
assign n16877 =  ( n79 ) & ( n15807 )  ;
assign n16878 =  ( n79 ) & ( n15809 )  ;
assign n16879 =  ( n79 ) & ( n15811 )  ;
assign n16880 =  ( n79 ) & ( n15813 )  ;
assign n16881 =  ( n80 ) & ( n15783 )  ;
assign n16882 =  ( n80 ) & ( n15785 )  ;
assign n16883 =  ( n80 ) & ( n15787 )  ;
assign n16884 =  ( n80 ) & ( n15789 )  ;
assign n16885 =  ( n80 ) & ( n15791 )  ;
assign n16886 =  ( n80 ) & ( n15793 )  ;
assign n16887 =  ( n80 ) & ( n15795 )  ;
assign n16888 =  ( n80 ) & ( n15797 )  ;
assign n16889 =  ( n80 ) & ( n15799 )  ;
assign n16890 =  ( n80 ) & ( n15801 )  ;
assign n16891 =  ( n80 ) & ( n15803 )  ;
assign n16892 =  ( n80 ) & ( n15805 )  ;
assign n16893 =  ( n80 ) & ( n15807 )  ;
assign n16894 =  ( n80 ) & ( n15809 )  ;
assign n16895 =  ( n80 ) & ( n15811 )  ;
assign n16896 =  ( n80 ) & ( n15813 )  ;
assign n16897 =  ( n81 ) & ( n15783 )  ;
assign n16898 =  ( n81 ) & ( n15785 )  ;
assign n16899 =  ( n81 ) & ( n15787 )  ;
assign n16900 =  ( n81 ) & ( n15789 )  ;
assign n16901 =  ( n81 ) & ( n15791 )  ;
assign n16902 =  ( n81 ) & ( n15793 )  ;
assign n16903 =  ( n81 ) & ( n15795 )  ;
assign n16904 =  ( n81 ) & ( n15797 )  ;
assign n16905 =  ( n81 ) & ( n15799 )  ;
assign n16906 =  ( n81 ) & ( n15801 )  ;
assign n16907 =  ( n81 ) & ( n15803 )  ;
assign n16908 =  ( n81 ) & ( n15805 )  ;
assign n16909 =  ( n81 ) & ( n15807 )  ;
assign n16910 =  ( n81 ) & ( n15809 )  ;
assign n16911 =  ( n81 ) & ( n15811 )  ;
assign n16912 =  ( n81 ) & ( n15813 )  ;
assign n16913 =  ( n82 ) & ( n15783 )  ;
assign n16914 =  ( n82 ) & ( n15785 )  ;
assign n16915 =  ( n82 ) & ( n15787 )  ;
assign n16916 =  ( n82 ) & ( n15789 )  ;
assign n16917 =  ( n82 ) & ( n15791 )  ;
assign n16918 =  ( n82 ) & ( n15793 )  ;
assign n16919 =  ( n82 ) & ( n15795 )  ;
assign n16920 =  ( n82 ) & ( n15797 )  ;
assign n16921 =  ( n82 ) & ( n15799 )  ;
assign n16922 =  ( n82 ) & ( n15801 )  ;
assign n16923 =  ( n82 ) & ( n15803 )  ;
assign n16924 =  ( n82 ) & ( n15805 )  ;
assign n16925 =  ( n82 ) & ( n15807 )  ;
assign n16926 =  ( n82 ) & ( n15809 )  ;
assign n16927 =  ( n82 ) & ( n15811 )  ;
assign n16928 =  ( n82 ) & ( n15813 )  ;
assign n16929 =  ( n83 ) & ( n15783 )  ;
assign n16930 =  ( n83 ) & ( n15785 )  ;
assign n16931 =  ( n83 ) & ( n15787 )  ;
assign n16932 =  ( n83 ) & ( n15789 )  ;
assign n16933 =  ( n83 ) & ( n15791 )  ;
assign n16934 =  ( n83 ) & ( n15793 )  ;
assign n16935 =  ( n83 ) & ( n15795 )  ;
assign n16936 =  ( n83 ) & ( n15797 )  ;
assign n16937 =  ( n83 ) & ( n15799 )  ;
assign n16938 =  ( n83 ) & ( n15801 )  ;
assign n16939 =  ( n83 ) & ( n15803 )  ;
assign n16940 =  ( n83 ) & ( n15805 )  ;
assign n16941 =  ( n83 ) & ( n15807 )  ;
assign n16942 =  ( n83 ) & ( n15809 )  ;
assign n16943 =  ( n83 ) & ( n15811 )  ;
assign n16944 =  ( n83 ) & ( n15813 )  ;
assign n16945 =  ( n84 ) & ( n15783 )  ;
assign n16946 =  ( n84 ) & ( n15785 )  ;
assign n16947 =  ( n84 ) & ( n15787 )  ;
assign n16948 =  ( n84 ) & ( n15789 )  ;
assign n16949 =  ( n84 ) & ( n15791 )  ;
assign n16950 =  ( n84 ) & ( n15793 )  ;
assign n16951 =  ( n84 ) & ( n15795 )  ;
assign n16952 =  ( n84 ) & ( n15797 )  ;
assign n16953 =  ( n84 ) & ( n15799 )  ;
assign n16954 =  ( n84 ) & ( n15801 )  ;
assign n16955 =  ( n84 ) & ( n15803 )  ;
assign n16956 =  ( n84 ) & ( n15805 )  ;
assign n16957 =  ( n84 ) & ( n15807 )  ;
assign n16958 =  ( n84 ) & ( n15809 )  ;
assign n16959 =  ( n84 ) & ( n15811 )  ;
assign n16960 =  ( n84 ) & ( n15813 )  ;
assign n16961 =  ( n85 ) & ( n15783 )  ;
assign n16962 =  ( n85 ) & ( n15785 )  ;
assign n16963 =  ( n85 ) & ( n15787 )  ;
assign n16964 =  ( n85 ) & ( n15789 )  ;
assign n16965 =  ( n85 ) & ( n15791 )  ;
assign n16966 =  ( n85 ) & ( n15793 )  ;
assign n16967 =  ( n85 ) & ( n15795 )  ;
assign n16968 =  ( n85 ) & ( n15797 )  ;
assign n16969 =  ( n85 ) & ( n15799 )  ;
assign n16970 =  ( n85 ) & ( n15801 )  ;
assign n16971 =  ( n85 ) & ( n15803 )  ;
assign n16972 =  ( n85 ) & ( n15805 )  ;
assign n16973 =  ( n85 ) & ( n15807 )  ;
assign n16974 =  ( n85 ) & ( n15809 )  ;
assign n16975 =  ( n85 ) & ( n15811 )  ;
assign n16976 =  ( n85 ) & ( n15813 )  ;
assign n16977 =  ( n86 ) & ( n15783 )  ;
assign n16978 =  ( n86 ) & ( n15785 )  ;
assign n16979 =  ( n86 ) & ( n15787 )  ;
assign n16980 =  ( n86 ) & ( n15789 )  ;
assign n16981 =  ( n86 ) & ( n15791 )  ;
assign n16982 =  ( n86 ) & ( n15793 )  ;
assign n16983 =  ( n86 ) & ( n15795 )  ;
assign n16984 =  ( n86 ) & ( n15797 )  ;
assign n16985 =  ( n86 ) & ( n15799 )  ;
assign n16986 =  ( n86 ) & ( n15801 )  ;
assign n16987 =  ( n86 ) & ( n15803 )  ;
assign n16988 =  ( n86 ) & ( n15805 )  ;
assign n16989 =  ( n86 ) & ( n15807 )  ;
assign n16990 =  ( n86 ) & ( n15809 )  ;
assign n16991 =  ( n86 ) & ( n15811 )  ;
assign n16992 =  ( n86 ) & ( n15813 )  ;
assign n16993 =  ( n87 ) & ( n15783 )  ;
assign n16994 =  ( n87 ) & ( n15785 )  ;
assign n16995 =  ( n87 ) & ( n15787 )  ;
assign n16996 =  ( n87 ) & ( n15789 )  ;
assign n16997 =  ( n87 ) & ( n15791 )  ;
assign n16998 =  ( n87 ) & ( n15793 )  ;
assign n16999 =  ( n87 ) & ( n15795 )  ;
assign n17000 =  ( n87 ) & ( n15797 )  ;
assign n17001 =  ( n87 ) & ( n15799 )  ;
assign n17002 =  ( n87 ) & ( n15801 )  ;
assign n17003 =  ( n87 ) & ( n15803 )  ;
assign n17004 =  ( n87 ) & ( n15805 )  ;
assign n17005 =  ( n87 ) & ( n15807 )  ;
assign n17006 =  ( n87 ) & ( n15809 )  ;
assign n17007 =  ( n87 ) & ( n15811 )  ;
assign n17008 =  ( n87 ) & ( n15813 )  ;
assign n17009 =  ( n88 ) & ( n15783 )  ;
assign n17010 =  ( n88 ) & ( n15785 )  ;
assign n17011 =  ( n88 ) & ( n15787 )  ;
assign n17012 =  ( n88 ) & ( n15789 )  ;
assign n17013 =  ( n88 ) & ( n15791 )  ;
assign n17014 =  ( n88 ) & ( n15793 )  ;
assign n17015 =  ( n88 ) & ( n15795 )  ;
assign n17016 =  ( n88 ) & ( n15797 )  ;
assign n17017 =  ( n88 ) & ( n15799 )  ;
assign n17018 =  ( n88 ) & ( n15801 )  ;
assign n17019 =  ( n88 ) & ( n15803 )  ;
assign n17020 =  ( n88 ) & ( n15805 )  ;
assign n17021 =  ( n88 ) & ( n15807 )  ;
assign n17022 =  ( n88 ) & ( n15809 )  ;
assign n17023 =  ( n88 ) & ( n15811 )  ;
assign n17024 =  ( n88 ) & ( n15813 )  ;
assign n17025 =  ( n89 ) & ( n15783 )  ;
assign n17026 =  ( n89 ) & ( n15785 )  ;
assign n17027 =  ( n89 ) & ( n15787 )  ;
assign n17028 =  ( n89 ) & ( n15789 )  ;
assign n17029 =  ( n89 ) & ( n15791 )  ;
assign n17030 =  ( n89 ) & ( n15793 )  ;
assign n17031 =  ( n89 ) & ( n15795 )  ;
assign n17032 =  ( n89 ) & ( n15797 )  ;
assign n17033 =  ( n89 ) & ( n15799 )  ;
assign n17034 =  ( n89 ) & ( n15801 )  ;
assign n17035 =  ( n89 ) & ( n15803 )  ;
assign n17036 =  ( n89 ) & ( n15805 )  ;
assign n17037 =  ( n89 ) & ( n15807 )  ;
assign n17038 =  ( n89 ) & ( n15809 )  ;
assign n17039 =  ( n89 ) & ( n15811 )  ;
assign n17040 =  ( n89 ) & ( n15813 )  ;
assign n17041 =  ( n90 ) & ( n15783 )  ;
assign n17042 =  ( n90 ) & ( n15785 )  ;
assign n17043 =  ( n90 ) & ( n15787 )  ;
assign n17044 =  ( n90 ) & ( n15789 )  ;
assign n17045 =  ( n90 ) & ( n15791 )  ;
assign n17046 =  ( n90 ) & ( n15793 )  ;
assign n17047 =  ( n90 ) & ( n15795 )  ;
assign n17048 =  ( n90 ) & ( n15797 )  ;
assign n17049 =  ( n90 ) & ( n15799 )  ;
assign n17050 =  ( n90 ) & ( n15801 )  ;
assign n17051 =  ( n90 ) & ( n15803 )  ;
assign n17052 =  ( n90 ) & ( n15805 )  ;
assign n17053 =  ( n90 ) & ( n15807 )  ;
assign n17054 =  ( n90 ) & ( n15809 )  ;
assign n17055 =  ( n90 ) & ( n15811 )  ;
assign n17056 =  ( n90 ) & ( n15813 )  ;
assign n17057 =  ( n91 ) & ( n15783 )  ;
assign n17058 =  ( n91 ) & ( n15785 )  ;
assign n17059 =  ( n91 ) & ( n15787 )  ;
assign n17060 =  ( n91 ) & ( n15789 )  ;
assign n17061 =  ( n91 ) & ( n15791 )  ;
assign n17062 =  ( n91 ) & ( n15793 )  ;
assign n17063 =  ( n91 ) & ( n15795 )  ;
assign n17064 =  ( n91 ) & ( n15797 )  ;
assign n17065 =  ( n91 ) & ( n15799 )  ;
assign n17066 =  ( n91 ) & ( n15801 )  ;
assign n17067 =  ( n91 ) & ( n15803 )  ;
assign n17068 =  ( n91 ) & ( n15805 )  ;
assign n17069 =  ( n91 ) & ( n15807 )  ;
assign n17070 =  ( n91 ) & ( n15809 )  ;
assign n17071 =  ( n91 ) & ( n15811 )  ;
assign n17072 =  ( n91 ) & ( n15813 )  ;
assign n17073 =  ( n92 ) & ( n15783 )  ;
assign n17074 =  ( n92 ) & ( n15785 )  ;
assign n17075 =  ( n92 ) & ( n15787 )  ;
assign n17076 =  ( n92 ) & ( n15789 )  ;
assign n17077 =  ( n92 ) & ( n15791 )  ;
assign n17078 =  ( n92 ) & ( n15793 )  ;
assign n17079 =  ( n92 ) & ( n15795 )  ;
assign n17080 =  ( n92 ) & ( n15797 )  ;
assign n17081 =  ( n92 ) & ( n15799 )  ;
assign n17082 =  ( n92 ) & ( n15801 )  ;
assign n17083 =  ( n92 ) & ( n15803 )  ;
assign n17084 =  ( n92 ) & ( n15805 )  ;
assign n17085 =  ( n92 ) & ( n15807 )  ;
assign n17086 =  ( n92 ) & ( n15809 )  ;
assign n17087 =  ( n92 ) & ( n15811 )  ;
assign n17088 =  ( n92 ) & ( n15813 )  ;
assign n17089 =  ( n93 ) & ( n15783 )  ;
assign n17090 =  ( n93 ) & ( n15785 )  ;
assign n17091 =  ( n93 ) & ( n15787 )  ;
assign n17092 =  ( n93 ) & ( n15789 )  ;
assign n17093 =  ( n93 ) & ( n15791 )  ;
assign n17094 =  ( n93 ) & ( n15793 )  ;
assign n17095 =  ( n93 ) & ( n15795 )  ;
assign n17096 =  ( n93 ) & ( n15797 )  ;
assign n17097 =  ( n93 ) & ( n15799 )  ;
assign n17098 =  ( n93 ) & ( n15801 )  ;
assign n17099 =  ( n93 ) & ( n15803 )  ;
assign n17100 =  ( n93 ) & ( n15805 )  ;
assign n17101 =  ( n93 ) & ( n15807 )  ;
assign n17102 =  ( n93 ) & ( n15809 )  ;
assign n17103 =  ( n93 ) & ( n15811 )  ;
assign n17104 =  ( n93 ) & ( n15813 )  ;
assign n17105 =  ( n94 ) & ( n15783 )  ;
assign n17106 =  ( n94 ) & ( n15785 )  ;
assign n17107 =  ( n94 ) & ( n15787 )  ;
assign n17108 =  ( n94 ) & ( n15789 )  ;
assign n17109 =  ( n94 ) & ( n15791 )  ;
assign n17110 =  ( n94 ) & ( n15793 )  ;
assign n17111 =  ( n94 ) & ( n15795 )  ;
assign n17112 =  ( n94 ) & ( n15797 )  ;
assign n17113 =  ( n94 ) & ( n15799 )  ;
assign n17114 =  ( n94 ) & ( n15801 )  ;
assign n17115 =  ( n94 ) & ( n15803 )  ;
assign n17116 =  ( n94 ) & ( n15805 )  ;
assign n17117 =  ( n94 ) & ( n15807 )  ;
assign n17118 =  ( n94 ) & ( n15809 )  ;
assign n17119 =  ( n94 ) & ( n15811 )  ;
assign n17120 =  ( n94 ) & ( n15813 )  ;
assign n17121 =  ( n95 ) & ( n15783 )  ;
assign n17122 =  ( n95 ) & ( n15785 )  ;
assign n17123 =  ( n95 ) & ( n15787 )  ;
assign n17124 =  ( n95 ) & ( n15789 )  ;
assign n17125 =  ( n95 ) & ( n15791 )  ;
assign n17126 =  ( n95 ) & ( n15793 )  ;
assign n17127 =  ( n95 ) & ( n15795 )  ;
assign n17128 =  ( n95 ) & ( n15797 )  ;
assign n17129 =  ( n95 ) & ( n15799 )  ;
assign n17130 =  ( n95 ) & ( n15801 )  ;
assign n17131 =  ( n95 ) & ( n15803 )  ;
assign n17132 =  ( n95 ) & ( n15805 )  ;
assign n17133 =  ( n95 ) & ( n15807 )  ;
assign n17134 =  ( n95 ) & ( n15809 )  ;
assign n17135 =  ( n95 ) & ( n15811 )  ;
assign n17136 =  ( n95 ) & ( n15813 )  ;
assign n17137 =  ( n96 ) & ( n15783 )  ;
assign n17138 =  ( n96 ) & ( n15785 )  ;
assign n17139 =  ( n96 ) & ( n15787 )  ;
assign n17140 =  ( n96 ) & ( n15789 )  ;
assign n17141 =  ( n96 ) & ( n15791 )  ;
assign n17142 =  ( n96 ) & ( n15793 )  ;
assign n17143 =  ( n96 ) & ( n15795 )  ;
assign n17144 =  ( n96 ) & ( n15797 )  ;
assign n17145 =  ( n96 ) & ( n15799 )  ;
assign n17146 =  ( n96 ) & ( n15801 )  ;
assign n17147 =  ( n96 ) & ( n15803 )  ;
assign n17148 =  ( n96 ) & ( n15805 )  ;
assign n17149 =  ( n96 ) & ( n15807 )  ;
assign n17150 =  ( n96 ) & ( n15809 )  ;
assign n17151 =  ( n96 ) & ( n15811 )  ;
assign n17152 =  ( n96 ) & ( n15813 )  ;
assign n17153 =  ( n97 ) & ( n15783 )  ;
assign n17154 =  ( n97 ) & ( n15785 )  ;
assign n17155 =  ( n97 ) & ( n15787 )  ;
assign n17156 =  ( n97 ) & ( n15789 )  ;
assign n17157 =  ( n97 ) & ( n15791 )  ;
assign n17158 =  ( n97 ) & ( n15793 )  ;
assign n17159 =  ( n97 ) & ( n15795 )  ;
assign n17160 =  ( n97 ) & ( n15797 )  ;
assign n17161 =  ( n97 ) & ( n15799 )  ;
assign n17162 =  ( n97 ) & ( n15801 )  ;
assign n17163 =  ( n97 ) & ( n15803 )  ;
assign n17164 =  ( n97 ) & ( n15805 )  ;
assign n17165 =  ( n97 ) & ( n15807 )  ;
assign n17166 =  ( n97 ) & ( n15809 )  ;
assign n17167 =  ( n97 ) & ( n15811 )  ;
assign n17168 =  ( n97 ) & ( n15813 )  ;
assign n17169 =  ( n98 ) & ( n15783 )  ;
assign n17170 =  ( n98 ) & ( n15785 )  ;
assign n17171 =  ( n98 ) & ( n15787 )  ;
assign n17172 =  ( n98 ) & ( n15789 )  ;
assign n17173 =  ( n98 ) & ( n15791 )  ;
assign n17174 =  ( n98 ) & ( n15793 )  ;
assign n17175 =  ( n98 ) & ( n15795 )  ;
assign n17176 =  ( n98 ) & ( n15797 )  ;
assign n17177 =  ( n98 ) & ( n15799 )  ;
assign n17178 =  ( n98 ) & ( n15801 )  ;
assign n17179 =  ( n98 ) & ( n15803 )  ;
assign n17180 =  ( n98 ) & ( n15805 )  ;
assign n17181 =  ( n98 ) & ( n15807 )  ;
assign n17182 =  ( n98 ) & ( n15809 )  ;
assign n17183 =  ( n98 ) & ( n15811 )  ;
assign n17184 =  ( n98 ) & ( n15813 )  ;
assign n17185 =  ( n99 ) & ( n15783 )  ;
assign n17186 =  ( n99 ) & ( n15785 )  ;
assign n17187 =  ( n99 ) & ( n15787 )  ;
assign n17188 =  ( n99 ) & ( n15789 )  ;
assign n17189 =  ( n99 ) & ( n15791 )  ;
assign n17190 =  ( n99 ) & ( n15793 )  ;
assign n17191 =  ( n99 ) & ( n15795 )  ;
assign n17192 =  ( n99 ) & ( n15797 )  ;
assign n17193 =  ( n99 ) & ( n15799 )  ;
assign n17194 =  ( n99 ) & ( n15801 )  ;
assign n17195 =  ( n99 ) & ( n15803 )  ;
assign n17196 =  ( n99 ) & ( n15805 )  ;
assign n17197 =  ( n99 ) & ( n15807 )  ;
assign n17198 =  ( n99 ) & ( n15809 )  ;
assign n17199 =  ( n99 ) & ( n15811 )  ;
assign n17200 =  ( n99 ) & ( n15813 )  ;
assign n17201 =  ( n100 ) & ( n15783 )  ;
assign n17202 =  ( n100 ) & ( n15785 )  ;
assign n17203 =  ( n100 ) & ( n15787 )  ;
assign n17204 =  ( n100 ) & ( n15789 )  ;
assign n17205 =  ( n100 ) & ( n15791 )  ;
assign n17206 =  ( n100 ) & ( n15793 )  ;
assign n17207 =  ( n100 ) & ( n15795 )  ;
assign n17208 =  ( n100 ) & ( n15797 )  ;
assign n17209 =  ( n100 ) & ( n15799 )  ;
assign n17210 =  ( n100 ) & ( n15801 )  ;
assign n17211 =  ( n100 ) & ( n15803 )  ;
assign n17212 =  ( n100 ) & ( n15805 )  ;
assign n17213 =  ( n100 ) & ( n15807 )  ;
assign n17214 =  ( n100 ) & ( n15809 )  ;
assign n17215 =  ( n100 ) & ( n15811 )  ;
assign n17216 =  ( n100 ) & ( n15813 )  ;
assign n17217 =  ( n101 ) & ( n15783 )  ;
assign n17218 =  ( n101 ) & ( n15785 )  ;
assign n17219 =  ( n101 ) & ( n15787 )  ;
assign n17220 =  ( n101 ) & ( n15789 )  ;
assign n17221 =  ( n101 ) & ( n15791 )  ;
assign n17222 =  ( n101 ) & ( n15793 )  ;
assign n17223 =  ( n101 ) & ( n15795 )  ;
assign n17224 =  ( n101 ) & ( n15797 )  ;
assign n17225 =  ( n101 ) & ( n15799 )  ;
assign n17226 =  ( n101 ) & ( n15801 )  ;
assign n17227 =  ( n101 ) & ( n15803 )  ;
assign n17228 =  ( n101 ) & ( n15805 )  ;
assign n17229 =  ( n101 ) & ( n15807 )  ;
assign n17230 =  ( n101 ) & ( n15809 )  ;
assign n17231 =  ( n101 ) & ( n15811 )  ;
assign n17232 =  ( n101 ) & ( n15813 )  ;
assign n17233 =  ( n102 ) & ( n15783 )  ;
assign n17234 =  ( n102 ) & ( n15785 )  ;
assign n17235 =  ( n102 ) & ( n15787 )  ;
assign n17236 =  ( n102 ) & ( n15789 )  ;
assign n17237 =  ( n102 ) & ( n15791 )  ;
assign n17238 =  ( n102 ) & ( n15793 )  ;
assign n17239 =  ( n102 ) & ( n15795 )  ;
assign n17240 =  ( n102 ) & ( n15797 )  ;
assign n17241 =  ( n102 ) & ( n15799 )  ;
assign n17242 =  ( n102 ) & ( n15801 )  ;
assign n17243 =  ( n102 ) & ( n15803 )  ;
assign n17244 =  ( n102 ) & ( n15805 )  ;
assign n17245 =  ( n102 ) & ( n15807 )  ;
assign n17246 =  ( n102 ) & ( n15809 )  ;
assign n17247 =  ( n102 ) & ( n15811 )  ;
assign n17248 =  ( n102 ) & ( n15813 )  ;
assign n17249 =  ( n103 ) & ( n15783 )  ;
assign n17250 =  ( n103 ) & ( n15785 )  ;
assign n17251 =  ( n103 ) & ( n15787 )  ;
assign n17252 =  ( n103 ) & ( n15789 )  ;
assign n17253 =  ( n103 ) & ( n15791 )  ;
assign n17254 =  ( n103 ) & ( n15793 )  ;
assign n17255 =  ( n103 ) & ( n15795 )  ;
assign n17256 =  ( n103 ) & ( n15797 )  ;
assign n17257 =  ( n103 ) & ( n15799 )  ;
assign n17258 =  ( n103 ) & ( n15801 )  ;
assign n17259 =  ( n103 ) & ( n15803 )  ;
assign n17260 =  ( n103 ) & ( n15805 )  ;
assign n17261 =  ( n103 ) & ( n15807 )  ;
assign n17262 =  ( n103 ) & ( n15809 )  ;
assign n17263 =  ( n103 ) & ( n15811 )  ;
assign n17264 =  ( n103 ) & ( n15813 )  ;
assign n17265 =  ( n104 ) & ( n15783 )  ;
assign n17266 =  ( n104 ) & ( n15785 )  ;
assign n17267 =  ( n104 ) & ( n15787 )  ;
assign n17268 =  ( n104 ) & ( n15789 )  ;
assign n17269 =  ( n104 ) & ( n15791 )  ;
assign n17270 =  ( n104 ) & ( n15793 )  ;
assign n17271 =  ( n104 ) & ( n15795 )  ;
assign n17272 =  ( n104 ) & ( n15797 )  ;
assign n17273 =  ( n104 ) & ( n15799 )  ;
assign n17274 =  ( n104 ) & ( n15801 )  ;
assign n17275 =  ( n104 ) & ( n15803 )  ;
assign n17276 =  ( n104 ) & ( n15805 )  ;
assign n17277 =  ( n104 ) & ( n15807 )  ;
assign n17278 =  ( n104 ) & ( n15809 )  ;
assign n17279 =  ( n104 ) & ( n15811 )  ;
assign n17280 =  ( n104 ) & ( n15813 )  ;
assign n17281 =  ( n105 ) & ( n15783 )  ;
assign n17282 =  ( n105 ) & ( n15785 )  ;
assign n17283 =  ( n105 ) & ( n15787 )  ;
assign n17284 =  ( n105 ) & ( n15789 )  ;
assign n17285 =  ( n105 ) & ( n15791 )  ;
assign n17286 =  ( n105 ) & ( n15793 )  ;
assign n17287 =  ( n105 ) & ( n15795 )  ;
assign n17288 =  ( n105 ) & ( n15797 )  ;
assign n17289 =  ( n105 ) & ( n15799 )  ;
assign n17290 =  ( n105 ) & ( n15801 )  ;
assign n17291 =  ( n105 ) & ( n15803 )  ;
assign n17292 =  ( n105 ) & ( n15805 )  ;
assign n17293 =  ( n105 ) & ( n15807 )  ;
assign n17294 =  ( n105 ) & ( n15809 )  ;
assign n17295 =  ( n105 ) & ( n15811 )  ;
assign n17296 =  ( n105 ) & ( n15813 )  ;
assign n17297 =  ( n106 ) & ( n15783 )  ;
assign n17298 =  ( n106 ) & ( n15785 )  ;
assign n17299 =  ( n106 ) & ( n15787 )  ;
assign n17300 =  ( n106 ) & ( n15789 )  ;
assign n17301 =  ( n106 ) & ( n15791 )  ;
assign n17302 =  ( n106 ) & ( n15793 )  ;
assign n17303 =  ( n106 ) & ( n15795 )  ;
assign n17304 =  ( n106 ) & ( n15797 )  ;
assign n17305 =  ( n106 ) & ( n15799 )  ;
assign n17306 =  ( n106 ) & ( n15801 )  ;
assign n17307 =  ( n106 ) & ( n15803 )  ;
assign n17308 =  ( n106 ) & ( n15805 )  ;
assign n17309 =  ( n106 ) & ( n15807 )  ;
assign n17310 =  ( n106 ) & ( n15809 )  ;
assign n17311 =  ( n106 ) & ( n15811 )  ;
assign n17312 =  ( n106 ) & ( n15813 )  ;
assign n17313 =  ( n107 ) & ( n15783 )  ;
assign n17314 =  ( n107 ) & ( n15785 )  ;
assign n17315 =  ( n107 ) & ( n15787 )  ;
assign n17316 =  ( n107 ) & ( n15789 )  ;
assign n17317 =  ( n107 ) & ( n15791 )  ;
assign n17318 =  ( n107 ) & ( n15793 )  ;
assign n17319 =  ( n107 ) & ( n15795 )  ;
assign n17320 =  ( n107 ) & ( n15797 )  ;
assign n17321 =  ( n107 ) & ( n15799 )  ;
assign n17322 =  ( n107 ) & ( n15801 )  ;
assign n17323 =  ( n107 ) & ( n15803 )  ;
assign n17324 =  ( n107 ) & ( n15805 )  ;
assign n17325 =  ( n107 ) & ( n15807 )  ;
assign n17326 =  ( n107 ) & ( n15809 )  ;
assign n17327 =  ( n107 ) & ( n15811 )  ;
assign n17328 =  ( n107 ) & ( n15813 )  ;
assign n17329 =  ( n108 ) & ( n15783 )  ;
assign n17330 =  ( n108 ) & ( n15785 )  ;
assign n17331 =  ( n108 ) & ( n15787 )  ;
assign n17332 =  ( n108 ) & ( n15789 )  ;
assign n17333 =  ( n108 ) & ( n15791 )  ;
assign n17334 =  ( n108 ) & ( n15793 )  ;
assign n17335 =  ( n108 ) & ( n15795 )  ;
assign n17336 =  ( n108 ) & ( n15797 )  ;
assign n17337 =  ( n108 ) & ( n15799 )  ;
assign n17338 =  ( n108 ) & ( n15801 )  ;
assign n17339 =  ( n108 ) & ( n15803 )  ;
assign n17340 =  ( n108 ) & ( n15805 )  ;
assign n17341 =  ( n108 ) & ( n15807 )  ;
assign n17342 =  ( n108 ) & ( n15809 )  ;
assign n17343 =  ( n108 ) & ( n15811 )  ;
assign n17344 =  ( n108 ) & ( n15813 )  ;
assign n17345 =  ( n17344 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n17346 =  ( n17343 ) ? ( VREG_0_1 ) : ( n17345 ) ;
assign n17347 =  ( n17342 ) ? ( VREG_0_2 ) : ( n17346 ) ;
assign n17348 =  ( n17341 ) ? ( VREG_0_3 ) : ( n17347 ) ;
assign n17349 =  ( n17340 ) ? ( VREG_0_4 ) : ( n17348 ) ;
assign n17350 =  ( n17339 ) ? ( VREG_0_5 ) : ( n17349 ) ;
assign n17351 =  ( n17338 ) ? ( VREG_0_6 ) : ( n17350 ) ;
assign n17352 =  ( n17337 ) ? ( VREG_0_7 ) : ( n17351 ) ;
assign n17353 =  ( n17336 ) ? ( VREG_0_8 ) : ( n17352 ) ;
assign n17354 =  ( n17335 ) ? ( VREG_0_9 ) : ( n17353 ) ;
assign n17355 =  ( n17334 ) ? ( VREG_0_10 ) : ( n17354 ) ;
assign n17356 =  ( n17333 ) ? ( VREG_0_11 ) : ( n17355 ) ;
assign n17357 =  ( n17332 ) ? ( VREG_0_12 ) : ( n17356 ) ;
assign n17358 =  ( n17331 ) ? ( VREG_0_13 ) : ( n17357 ) ;
assign n17359 =  ( n17330 ) ? ( VREG_0_14 ) : ( n17358 ) ;
assign n17360 =  ( n17329 ) ? ( VREG_0_15 ) : ( n17359 ) ;
assign n17361 =  ( n17328 ) ? ( VREG_1_0 ) : ( n17360 ) ;
assign n17362 =  ( n17327 ) ? ( VREG_1_1 ) : ( n17361 ) ;
assign n17363 =  ( n17326 ) ? ( VREG_1_2 ) : ( n17362 ) ;
assign n17364 =  ( n17325 ) ? ( VREG_1_3 ) : ( n17363 ) ;
assign n17365 =  ( n17324 ) ? ( VREG_1_4 ) : ( n17364 ) ;
assign n17366 =  ( n17323 ) ? ( VREG_1_5 ) : ( n17365 ) ;
assign n17367 =  ( n17322 ) ? ( VREG_1_6 ) : ( n17366 ) ;
assign n17368 =  ( n17321 ) ? ( VREG_1_7 ) : ( n17367 ) ;
assign n17369 =  ( n17320 ) ? ( VREG_1_8 ) : ( n17368 ) ;
assign n17370 =  ( n17319 ) ? ( VREG_1_9 ) : ( n17369 ) ;
assign n17371 =  ( n17318 ) ? ( VREG_1_10 ) : ( n17370 ) ;
assign n17372 =  ( n17317 ) ? ( VREG_1_11 ) : ( n17371 ) ;
assign n17373 =  ( n17316 ) ? ( VREG_1_12 ) : ( n17372 ) ;
assign n17374 =  ( n17315 ) ? ( VREG_1_13 ) : ( n17373 ) ;
assign n17375 =  ( n17314 ) ? ( VREG_1_14 ) : ( n17374 ) ;
assign n17376 =  ( n17313 ) ? ( VREG_1_15 ) : ( n17375 ) ;
assign n17377 =  ( n17312 ) ? ( VREG_2_0 ) : ( n17376 ) ;
assign n17378 =  ( n17311 ) ? ( VREG_2_1 ) : ( n17377 ) ;
assign n17379 =  ( n17310 ) ? ( VREG_2_2 ) : ( n17378 ) ;
assign n17380 =  ( n17309 ) ? ( VREG_2_3 ) : ( n17379 ) ;
assign n17381 =  ( n17308 ) ? ( VREG_2_4 ) : ( n17380 ) ;
assign n17382 =  ( n17307 ) ? ( VREG_2_5 ) : ( n17381 ) ;
assign n17383 =  ( n17306 ) ? ( VREG_2_6 ) : ( n17382 ) ;
assign n17384 =  ( n17305 ) ? ( VREG_2_7 ) : ( n17383 ) ;
assign n17385 =  ( n17304 ) ? ( VREG_2_8 ) : ( n17384 ) ;
assign n17386 =  ( n17303 ) ? ( VREG_2_9 ) : ( n17385 ) ;
assign n17387 =  ( n17302 ) ? ( VREG_2_10 ) : ( n17386 ) ;
assign n17388 =  ( n17301 ) ? ( VREG_2_11 ) : ( n17387 ) ;
assign n17389 =  ( n17300 ) ? ( VREG_2_12 ) : ( n17388 ) ;
assign n17390 =  ( n17299 ) ? ( VREG_2_13 ) : ( n17389 ) ;
assign n17391 =  ( n17298 ) ? ( VREG_2_14 ) : ( n17390 ) ;
assign n17392 =  ( n17297 ) ? ( VREG_2_15 ) : ( n17391 ) ;
assign n17393 =  ( n17296 ) ? ( VREG_3_0 ) : ( n17392 ) ;
assign n17394 =  ( n17295 ) ? ( VREG_3_1 ) : ( n17393 ) ;
assign n17395 =  ( n17294 ) ? ( VREG_3_2 ) : ( n17394 ) ;
assign n17396 =  ( n17293 ) ? ( VREG_3_3 ) : ( n17395 ) ;
assign n17397 =  ( n17292 ) ? ( VREG_3_4 ) : ( n17396 ) ;
assign n17398 =  ( n17291 ) ? ( VREG_3_5 ) : ( n17397 ) ;
assign n17399 =  ( n17290 ) ? ( VREG_3_6 ) : ( n17398 ) ;
assign n17400 =  ( n17289 ) ? ( VREG_3_7 ) : ( n17399 ) ;
assign n17401 =  ( n17288 ) ? ( VREG_3_8 ) : ( n17400 ) ;
assign n17402 =  ( n17287 ) ? ( VREG_3_9 ) : ( n17401 ) ;
assign n17403 =  ( n17286 ) ? ( VREG_3_10 ) : ( n17402 ) ;
assign n17404 =  ( n17285 ) ? ( VREG_3_11 ) : ( n17403 ) ;
assign n17405 =  ( n17284 ) ? ( VREG_3_12 ) : ( n17404 ) ;
assign n17406 =  ( n17283 ) ? ( VREG_3_13 ) : ( n17405 ) ;
assign n17407 =  ( n17282 ) ? ( VREG_3_14 ) : ( n17406 ) ;
assign n17408 =  ( n17281 ) ? ( VREG_3_15 ) : ( n17407 ) ;
assign n17409 =  ( n17280 ) ? ( VREG_4_0 ) : ( n17408 ) ;
assign n17410 =  ( n17279 ) ? ( VREG_4_1 ) : ( n17409 ) ;
assign n17411 =  ( n17278 ) ? ( VREG_4_2 ) : ( n17410 ) ;
assign n17412 =  ( n17277 ) ? ( VREG_4_3 ) : ( n17411 ) ;
assign n17413 =  ( n17276 ) ? ( VREG_4_4 ) : ( n17412 ) ;
assign n17414 =  ( n17275 ) ? ( VREG_4_5 ) : ( n17413 ) ;
assign n17415 =  ( n17274 ) ? ( VREG_4_6 ) : ( n17414 ) ;
assign n17416 =  ( n17273 ) ? ( VREG_4_7 ) : ( n17415 ) ;
assign n17417 =  ( n17272 ) ? ( VREG_4_8 ) : ( n17416 ) ;
assign n17418 =  ( n17271 ) ? ( VREG_4_9 ) : ( n17417 ) ;
assign n17419 =  ( n17270 ) ? ( VREG_4_10 ) : ( n17418 ) ;
assign n17420 =  ( n17269 ) ? ( VREG_4_11 ) : ( n17419 ) ;
assign n17421 =  ( n17268 ) ? ( VREG_4_12 ) : ( n17420 ) ;
assign n17422 =  ( n17267 ) ? ( VREG_4_13 ) : ( n17421 ) ;
assign n17423 =  ( n17266 ) ? ( VREG_4_14 ) : ( n17422 ) ;
assign n17424 =  ( n17265 ) ? ( VREG_4_15 ) : ( n17423 ) ;
assign n17425 =  ( n17264 ) ? ( VREG_5_0 ) : ( n17424 ) ;
assign n17426 =  ( n17263 ) ? ( VREG_5_1 ) : ( n17425 ) ;
assign n17427 =  ( n17262 ) ? ( VREG_5_2 ) : ( n17426 ) ;
assign n17428 =  ( n17261 ) ? ( VREG_5_3 ) : ( n17427 ) ;
assign n17429 =  ( n17260 ) ? ( VREG_5_4 ) : ( n17428 ) ;
assign n17430 =  ( n17259 ) ? ( VREG_5_5 ) : ( n17429 ) ;
assign n17431 =  ( n17258 ) ? ( VREG_5_6 ) : ( n17430 ) ;
assign n17432 =  ( n17257 ) ? ( VREG_5_7 ) : ( n17431 ) ;
assign n17433 =  ( n17256 ) ? ( VREG_5_8 ) : ( n17432 ) ;
assign n17434 =  ( n17255 ) ? ( VREG_5_9 ) : ( n17433 ) ;
assign n17435 =  ( n17254 ) ? ( VREG_5_10 ) : ( n17434 ) ;
assign n17436 =  ( n17253 ) ? ( VREG_5_11 ) : ( n17435 ) ;
assign n17437 =  ( n17252 ) ? ( VREG_5_12 ) : ( n17436 ) ;
assign n17438 =  ( n17251 ) ? ( VREG_5_13 ) : ( n17437 ) ;
assign n17439 =  ( n17250 ) ? ( VREG_5_14 ) : ( n17438 ) ;
assign n17440 =  ( n17249 ) ? ( VREG_5_15 ) : ( n17439 ) ;
assign n17441 =  ( n17248 ) ? ( VREG_6_0 ) : ( n17440 ) ;
assign n17442 =  ( n17247 ) ? ( VREG_6_1 ) : ( n17441 ) ;
assign n17443 =  ( n17246 ) ? ( VREG_6_2 ) : ( n17442 ) ;
assign n17444 =  ( n17245 ) ? ( VREG_6_3 ) : ( n17443 ) ;
assign n17445 =  ( n17244 ) ? ( VREG_6_4 ) : ( n17444 ) ;
assign n17446 =  ( n17243 ) ? ( VREG_6_5 ) : ( n17445 ) ;
assign n17447 =  ( n17242 ) ? ( VREG_6_6 ) : ( n17446 ) ;
assign n17448 =  ( n17241 ) ? ( VREG_6_7 ) : ( n17447 ) ;
assign n17449 =  ( n17240 ) ? ( VREG_6_8 ) : ( n17448 ) ;
assign n17450 =  ( n17239 ) ? ( VREG_6_9 ) : ( n17449 ) ;
assign n17451 =  ( n17238 ) ? ( VREG_6_10 ) : ( n17450 ) ;
assign n17452 =  ( n17237 ) ? ( VREG_6_11 ) : ( n17451 ) ;
assign n17453 =  ( n17236 ) ? ( VREG_6_12 ) : ( n17452 ) ;
assign n17454 =  ( n17235 ) ? ( VREG_6_13 ) : ( n17453 ) ;
assign n17455 =  ( n17234 ) ? ( VREG_6_14 ) : ( n17454 ) ;
assign n17456 =  ( n17233 ) ? ( VREG_6_15 ) : ( n17455 ) ;
assign n17457 =  ( n17232 ) ? ( VREG_7_0 ) : ( n17456 ) ;
assign n17458 =  ( n17231 ) ? ( VREG_7_1 ) : ( n17457 ) ;
assign n17459 =  ( n17230 ) ? ( VREG_7_2 ) : ( n17458 ) ;
assign n17460 =  ( n17229 ) ? ( VREG_7_3 ) : ( n17459 ) ;
assign n17461 =  ( n17228 ) ? ( VREG_7_4 ) : ( n17460 ) ;
assign n17462 =  ( n17227 ) ? ( VREG_7_5 ) : ( n17461 ) ;
assign n17463 =  ( n17226 ) ? ( VREG_7_6 ) : ( n17462 ) ;
assign n17464 =  ( n17225 ) ? ( VREG_7_7 ) : ( n17463 ) ;
assign n17465 =  ( n17224 ) ? ( VREG_7_8 ) : ( n17464 ) ;
assign n17466 =  ( n17223 ) ? ( VREG_7_9 ) : ( n17465 ) ;
assign n17467 =  ( n17222 ) ? ( VREG_7_10 ) : ( n17466 ) ;
assign n17468 =  ( n17221 ) ? ( VREG_7_11 ) : ( n17467 ) ;
assign n17469 =  ( n17220 ) ? ( VREG_7_12 ) : ( n17468 ) ;
assign n17470 =  ( n17219 ) ? ( VREG_7_13 ) : ( n17469 ) ;
assign n17471 =  ( n17218 ) ? ( VREG_7_14 ) : ( n17470 ) ;
assign n17472 =  ( n17217 ) ? ( VREG_7_15 ) : ( n17471 ) ;
assign n17473 =  ( n17216 ) ? ( VREG_8_0 ) : ( n17472 ) ;
assign n17474 =  ( n17215 ) ? ( VREG_8_1 ) : ( n17473 ) ;
assign n17475 =  ( n17214 ) ? ( VREG_8_2 ) : ( n17474 ) ;
assign n17476 =  ( n17213 ) ? ( VREG_8_3 ) : ( n17475 ) ;
assign n17477 =  ( n17212 ) ? ( VREG_8_4 ) : ( n17476 ) ;
assign n17478 =  ( n17211 ) ? ( VREG_8_5 ) : ( n17477 ) ;
assign n17479 =  ( n17210 ) ? ( VREG_8_6 ) : ( n17478 ) ;
assign n17480 =  ( n17209 ) ? ( VREG_8_7 ) : ( n17479 ) ;
assign n17481 =  ( n17208 ) ? ( VREG_8_8 ) : ( n17480 ) ;
assign n17482 =  ( n17207 ) ? ( VREG_8_9 ) : ( n17481 ) ;
assign n17483 =  ( n17206 ) ? ( VREG_8_10 ) : ( n17482 ) ;
assign n17484 =  ( n17205 ) ? ( VREG_8_11 ) : ( n17483 ) ;
assign n17485 =  ( n17204 ) ? ( VREG_8_12 ) : ( n17484 ) ;
assign n17486 =  ( n17203 ) ? ( VREG_8_13 ) : ( n17485 ) ;
assign n17487 =  ( n17202 ) ? ( VREG_8_14 ) : ( n17486 ) ;
assign n17488 =  ( n17201 ) ? ( VREG_8_15 ) : ( n17487 ) ;
assign n17489 =  ( n17200 ) ? ( VREG_9_0 ) : ( n17488 ) ;
assign n17490 =  ( n17199 ) ? ( VREG_9_1 ) : ( n17489 ) ;
assign n17491 =  ( n17198 ) ? ( VREG_9_2 ) : ( n17490 ) ;
assign n17492 =  ( n17197 ) ? ( VREG_9_3 ) : ( n17491 ) ;
assign n17493 =  ( n17196 ) ? ( VREG_9_4 ) : ( n17492 ) ;
assign n17494 =  ( n17195 ) ? ( VREG_9_5 ) : ( n17493 ) ;
assign n17495 =  ( n17194 ) ? ( VREG_9_6 ) : ( n17494 ) ;
assign n17496 =  ( n17193 ) ? ( VREG_9_7 ) : ( n17495 ) ;
assign n17497 =  ( n17192 ) ? ( VREG_9_8 ) : ( n17496 ) ;
assign n17498 =  ( n17191 ) ? ( VREG_9_9 ) : ( n17497 ) ;
assign n17499 =  ( n17190 ) ? ( VREG_9_10 ) : ( n17498 ) ;
assign n17500 =  ( n17189 ) ? ( VREG_9_11 ) : ( n17499 ) ;
assign n17501 =  ( n17188 ) ? ( VREG_9_12 ) : ( n17500 ) ;
assign n17502 =  ( n17187 ) ? ( VREG_9_13 ) : ( n17501 ) ;
assign n17503 =  ( n17186 ) ? ( VREG_9_14 ) : ( n17502 ) ;
assign n17504 =  ( n17185 ) ? ( VREG_9_15 ) : ( n17503 ) ;
assign n17505 =  ( n17184 ) ? ( VREG_10_0 ) : ( n17504 ) ;
assign n17506 =  ( n17183 ) ? ( VREG_10_1 ) : ( n17505 ) ;
assign n17507 =  ( n17182 ) ? ( VREG_10_2 ) : ( n17506 ) ;
assign n17508 =  ( n17181 ) ? ( VREG_10_3 ) : ( n17507 ) ;
assign n17509 =  ( n17180 ) ? ( VREG_10_4 ) : ( n17508 ) ;
assign n17510 =  ( n17179 ) ? ( VREG_10_5 ) : ( n17509 ) ;
assign n17511 =  ( n17178 ) ? ( VREG_10_6 ) : ( n17510 ) ;
assign n17512 =  ( n17177 ) ? ( VREG_10_7 ) : ( n17511 ) ;
assign n17513 =  ( n17176 ) ? ( VREG_10_8 ) : ( n17512 ) ;
assign n17514 =  ( n17175 ) ? ( VREG_10_9 ) : ( n17513 ) ;
assign n17515 =  ( n17174 ) ? ( VREG_10_10 ) : ( n17514 ) ;
assign n17516 =  ( n17173 ) ? ( VREG_10_11 ) : ( n17515 ) ;
assign n17517 =  ( n17172 ) ? ( VREG_10_12 ) : ( n17516 ) ;
assign n17518 =  ( n17171 ) ? ( VREG_10_13 ) : ( n17517 ) ;
assign n17519 =  ( n17170 ) ? ( VREG_10_14 ) : ( n17518 ) ;
assign n17520 =  ( n17169 ) ? ( VREG_10_15 ) : ( n17519 ) ;
assign n17521 =  ( n17168 ) ? ( VREG_11_0 ) : ( n17520 ) ;
assign n17522 =  ( n17167 ) ? ( VREG_11_1 ) : ( n17521 ) ;
assign n17523 =  ( n17166 ) ? ( VREG_11_2 ) : ( n17522 ) ;
assign n17524 =  ( n17165 ) ? ( VREG_11_3 ) : ( n17523 ) ;
assign n17525 =  ( n17164 ) ? ( VREG_11_4 ) : ( n17524 ) ;
assign n17526 =  ( n17163 ) ? ( VREG_11_5 ) : ( n17525 ) ;
assign n17527 =  ( n17162 ) ? ( VREG_11_6 ) : ( n17526 ) ;
assign n17528 =  ( n17161 ) ? ( VREG_11_7 ) : ( n17527 ) ;
assign n17529 =  ( n17160 ) ? ( VREG_11_8 ) : ( n17528 ) ;
assign n17530 =  ( n17159 ) ? ( VREG_11_9 ) : ( n17529 ) ;
assign n17531 =  ( n17158 ) ? ( VREG_11_10 ) : ( n17530 ) ;
assign n17532 =  ( n17157 ) ? ( VREG_11_11 ) : ( n17531 ) ;
assign n17533 =  ( n17156 ) ? ( VREG_11_12 ) : ( n17532 ) ;
assign n17534 =  ( n17155 ) ? ( VREG_11_13 ) : ( n17533 ) ;
assign n17535 =  ( n17154 ) ? ( VREG_11_14 ) : ( n17534 ) ;
assign n17536 =  ( n17153 ) ? ( VREG_11_15 ) : ( n17535 ) ;
assign n17537 =  ( n17152 ) ? ( VREG_12_0 ) : ( n17536 ) ;
assign n17538 =  ( n17151 ) ? ( VREG_12_1 ) : ( n17537 ) ;
assign n17539 =  ( n17150 ) ? ( VREG_12_2 ) : ( n17538 ) ;
assign n17540 =  ( n17149 ) ? ( VREG_12_3 ) : ( n17539 ) ;
assign n17541 =  ( n17148 ) ? ( VREG_12_4 ) : ( n17540 ) ;
assign n17542 =  ( n17147 ) ? ( VREG_12_5 ) : ( n17541 ) ;
assign n17543 =  ( n17146 ) ? ( VREG_12_6 ) : ( n17542 ) ;
assign n17544 =  ( n17145 ) ? ( VREG_12_7 ) : ( n17543 ) ;
assign n17545 =  ( n17144 ) ? ( VREG_12_8 ) : ( n17544 ) ;
assign n17546 =  ( n17143 ) ? ( VREG_12_9 ) : ( n17545 ) ;
assign n17547 =  ( n17142 ) ? ( VREG_12_10 ) : ( n17546 ) ;
assign n17548 =  ( n17141 ) ? ( VREG_12_11 ) : ( n17547 ) ;
assign n17549 =  ( n17140 ) ? ( VREG_12_12 ) : ( n17548 ) ;
assign n17550 =  ( n17139 ) ? ( VREG_12_13 ) : ( n17549 ) ;
assign n17551 =  ( n17138 ) ? ( VREG_12_14 ) : ( n17550 ) ;
assign n17552 =  ( n17137 ) ? ( VREG_12_15 ) : ( n17551 ) ;
assign n17553 =  ( n17136 ) ? ( VREG_13_0 ) : ( n17552 ) ;
assign n17554 =  ( n17135 ) ? ( VREG_13_1 ) : ( n17553 ) ;
assign n17555 =  ( n17134 ) ? ( VREG_13_2 ) : ( n17554 ) ;
assign n17556 =  ( n17133 ) ? ( VREG_13_3 ) : ( n17555 ) ;
assign n17557 =  ( n17132 ) ? ( VREG_13_4 ) : ( n17556 ) ;
assign n17558 =  ( n17131 ) ? ( VREG_13_5 ) : ( n17557 ) ;
assign n17559 =  ( n17130 ) ? ( VREG_13_6 ) : ( n17558 ) ;
assign n17560 =  ( n17129 ) ? ( VREG_13_7 ) : ( n17559 ) ;
assign n17561 =  ( n17128 ) ? ( VREG_13_8 ) : ( n17560 ) ;
assign n17562 =  ( n17127 ) ? ( VREG_13_9 ) : ( n17561 ) ;
assign n17563 =  ( n17126 ) ? ( VREG_13_10 ) : ( n17562 ) ;
assign n17564 =  ( n17125 ) ? ( VREG_13_11 ) : ( n17563 ) ;
assign n17565 =  ( n17124 ) ? ( VREG_13_12 ) : ( n17564 ) ;
assign n17566 =  ( n17123 ) ? ( VREG_13_13 ) : ( n17565 ) ;
assign n17567 =  ( n17122 ) ? ( VREG_13_14 ) : ( n17566 ) ;
assign n17568 =  ( n17121 ) ? ( VREG_13_15 ) : ( n17567 ) ;
assign n17569 =  ( n17120 ) ? ( VREG_14_0 ) : ( n17568 ) ;
assign n17570 =  ( n17119 ) ? ( VREG_14_1 ) : ( n17569 ) ;
assign n17571 =  ( n17118 ) ? ( VREG_14_2 ) : ( n17570 ) ;
assign n17572 =  ( n17117 ) ? ( VREG_14_3 ) : ( n17571 ) ;
assign n17573 =  ( n17116 ) ? ( VREG_14_4 ) : ( n17572 ) ;
assign n17574 =  ( n17115 ) ? ( VREG_14_5 ) : ( n17573 ) ;
assign n17575 =  ( n17114 ) ? ( VREG_14_6 ) : ( n17574 ) ;
assign n17576 =  ( n17113 ) ? ( VREG_14_7 ) : ( n17575 ) ;
assign n17577 =  ( n17112 ) ? ( VREG_14_8 ) : ( n17576 ) ;
assign n17578 =  ( n17111 ) ? ( VREG_14_9 ) : ( n17577 ) ;
assign n17579 =  ( n17110 ) ? ( VREG_14_10 ) : ( n17578 ) ;
assign n17580 =  ( n17109 ) ? ( VREG_14_11 ) : ( n17579 ) ;
assign n17581 =  ( n17108 ) ? ( VREG_14_12 ) : ( n17580 ) ;
assign n17582 =  ( n17107 ) ? ( VREG_14_13 ) : ( n17581 ) ;
assign n17583 =  ( n17106 ) ? ( VREG_14_14 ) : ( n17582 ) ;
assign n17584 =  ( n17105 ) ? ( VREG_14_15 ) : ( n17583 ) ;
assign n17585 =  ( n17104 ) ? ( VREG_15_0 ) : ( n17584 ) ;
assign n17586 =  ( n17103 ) ? ( VREG_15_1 ) : ( n17585 ) ;
assign n17587 =  ( n17102 ) ? ( VREG_15_2 ) : ( n17586 ) ;
assign n17588 =  ( n17101 ) ? ( VREG_15_3 ) : ( n17587 ) ;
assign n17589 =  ( n17100 ) ? ( VREG_15_4 ) : ( n17588 ) ;
assign n17590 =  ( n17099 ) ? ( VREG_15_5 ) : ( n17589 ) ;
assign n17591 =  ( n17098 ) ? ( VREG_15_6 ) : ( n17590 ) ;
assign n17592 =  ( n17097 ) ? ( VREG_15_7 ) : ( n17591 ) ;
assign n17593 =  ( n17096 ) ? ( VREG_15_8 ) : ( n17592 ) ;
assign n17594 =  ( n17095 ) ? ( VREG_15_9 ) : ( n17593 ) ;
assign n17595 =  ( n17094 ) ? ( VREG_15_10 ) : ( n17594 ) ;
assign n17596 =  ( n17093 ) ? ( VREG_15_11 ) : ( n17595 ) ;
assign n17597 =  ( n17092 ) ? ( VREG_15_12 ) : ( n17596 ) ;
assign n17598 =  ( n17091 ) ? ( VREG_15_13 ) : ( n17597 ) ;
assign n17599 =  ( n17090 ) ? ( VREG_15_14 ) : ( n17598 ) ;
assign n17600 =  ( n17089 ) ? ( VREG_15_15 ) : ( n17599 ) ;
assign n17601 =  ( n17088 ) ? ( VREG_16_0 ) : ( n17600 ) ;
assign n17602 =  ( n17087 ) ? ( VREG_16_1 ) : ( n17601 ) ;
assign n17603 =  ( n17086 ) ? ( VREG_16_2 ) : ( n17602 ) ;
assign n17604 =  ( n17085 ) ? ( VREG_16_3 ) : ( n17603 ) ;
assign n17605 =  ( n17084 ) ? ( VREG_16_4 ) : ( n17604 ) ;
assign n17606 =  ( n17083 ) ? ( VREG_16_5 ) : ( n17605 ) ;
assign n17607 =  ( n17082 ) ? ( VREG_16_6 ) : ( n17606 ) ;
assign n17608 =  ( n17081 ) ? ( VREG_16_7 ) : ( n17607 ) ;
assign n17609 =  ( n17080 ) ? ( VREG_16_8 ) : ( n17608 ) ;
assign n17610 =  ( n17079 ) ? ( VREG_16_9 ) : ( n17609 ) ;
assign n17611 =  ( n17078 ) ? ( VREG_16_10 ) : ( n17610 ) ;
assign n17612 =  ( n17077 ) ? ( VREG_16_11 ) : ( n17611 ) ;
assign n17613 =  ( n17076 ) ? ( VREG_16_12 ) : ( n17612 ) ;
assign n17614 =  ( n17075 ) ? ( VREG_16_13 ) : ( n17613 ) ;
assign n17615 =  ( n17074 ) ? ( VREG_16_14 ) : ( n17614 ) ;
assign n17616 =  ( n17073 ) ? ( VREG_16_15 ) : ( n17615 ) ;
assign n17617 =  ( n17072 ) ? ( VREG_17_0 ) : ( n17616 ) ;
assign n17618 =  ( n17071 ) ? ( VREG_17_1 ) : ( n17617 ) ;
assign n17619 =  ( n17070 ) ? ( VREG_17_2 ) : ( n17618 ) ;
assign n17620 =  ( n17069 ) ? ( VREG_17_3 ) : ( n17619 ) ;
assign n17621 =  ( n17068 ) ? ( VREG_17_4 ) : ( n17620 ) ;
assign n17622 =  ( n17067 ) ? ( VREG_17_5 ) : ( n17621 ) ;
assign n17623 =  ( n17066 ) ? ( VREG_17_6 ) : ( n17622 ) ;
assign n17624 =  ( n17065 ) ? ( VREG_17_7 ) : ( n17623 ) ;
assign n17625 =  ( n17064 ) ? ( VREG_17_8 ) : ( n17624 ) ;
assign n17626 =  ( n17063 ) ? ( VREG_17_9 ) : ( n17625 ) ;
assign n17627 =  ( n17062 ) ? ( VREG_17_10 ) : ( n17626 ) ;
assign n17628 =  ( n17061 ) ? ( VREG_17_11 ) : ( n17627 ) ;
assign n17629 =  ( n17060 ) ? ( VREG_17_12 ) : ( n17628 ) ;
assign n17630 =  ( n17059 ) ? ( VREG_17_13 ) : ( n17629 ) ;
assign n17631 =  ( n17058 ) ? ( VREG_17_14 ) : ( n17630 ) ;
assign n17632 =  ( n17057 ) ? ( VREG_17_15 ) : ( n17631 ) ;
assign n17633 =  ( n17056 ) ? ( VREG_18_0 ) : ( n17632 ) ;
assign n17634 =  ( n17055 ) ? ( VREG_18_1 ) : ( n17633 ) ;
assign n17635 =  ( n17054 ) ? ( VREG_18_2 ) : ( n17634 ) ;
assign n17636 =  ( n17053 ) ? ( VREG_18_3 ) : ( n17635 ) ;
assign n17637 =  ( n17052 ) ? ( VREG_18_4 ) : ( n17636 ) ;
assign n17638 =  ( n17051 ) ? ( VREG_18_5 ) : ( n17637 ) ;
assign n17639 =  ( n17050 ) ? ( VREG_18_6 ) : ( n17638 ) ;
assign n17640 =  ( n17049 ) ? ( VREG_18_7 ) : ( n17639 ) ;
assign n17641 =  ( n17048 ) ? ( VREG_18_8 ) : ( n17640 ) ;
assign n17642 =  ( n17047 ) ? ( VREG_18_9 ) : ( n17641 ) ;
assign n17643 =  ( n17046 ) ? ( VREG_18_10 ) : ( n17642 ) ;
assign n17644 =  ( n17045 ) ? ( VREG_18_11 ) : ( n17643 ) ;
assign n17645 =  ( n17044 ) ? ( VREG_18_12 ) : ( n17644 ) ;
assign n17646 =  ( n17043 ) ? ( VREG_18_13 ) : ( n17645 ) ;
assign n17647 =  ( n17042 ) ? ( VREG_18_14 ) : ( n17646 ) ;
assign n17648 =  ( n17041 ) ? ( VREG_18_15 ) : ( n17647 ) ;
assign n17649 =  ( n17040 ) ? ( VREG_19_0 ) : ( n17648 ) ;
assign n17650 =  ( n17039 ) ? ( VREG_19_1 ) : ( n17649 ) ;
assign n17651 =  ( n17038 ) ? ( VREG_19_2 ) : ( n17650 ) ;
assign n17652 =  ( n17037 ) ? ( VREG_19_3 ) : ( n17651 ) ;
assign n17653 =  ( n17036 ) ? ( VREG_19_4 ) : ( n17652 ) ;
assign n17654 =  ( n17035 ) ? ( VREG_19_5 ) : ( n17653 ) ;
assign n17655 =  ( n17034 ) ? ( VREG_19_6 ) : ( n17654 ) ;
assign n17656 =  ( n17033 ) ? ( VREG_19_7 ) : ( n17655 ) ;
assign n17657 =  ( n17032 ) ? ( VREG_19_8 ) : ( n17656 ) ;
assign n17658 =  ( n17031 ) ? ( VREG_19_9 ) : ( n17657 ) ;
assign n17659 =  ( n17030 ) ? ( VREG_19_10 ) : ( n17658 ) ;
assign n17660 =  ( n17029 ) ? ( VREG_19_11 ) : ( n17659 ) ;
assign n17661 =  ( n17028 ) ? ( VREG_19_12 ) : ( n17660 ) ;
assign n17662 =  ( n17027 ) ? ( VREG_19_13 ) : ( n17661 ) ;
assign n17663 =  ( n17026 ) ? ( VREG_19_14 ) : ( n17662 ) ;
assign n17664 =  ( n17025 ) ? ( VREG_19_15 ) : ( n17663 ) ;
assign n17665 =  ( n17024 ) ? ( VREG_20_0 ) : ( n17664 ) ;
assign n17666 =  ( n17023 ) ? ( VREG_20_1 ) : ( n17665 ) ;
assign n17667 =  ( n17022 ) ? ( VREG_20_2 ) : ( n17666 ) ;
assign n17668 =  ( n17021 ) ? ( VREG_20_3 ) : ( n17667 ) ;
assign n17669 =  ( n17020 ) ? ( VREG_20_4 ) : ( n17668 ) ;
assign n17670 =  ( n17019 ) ? ( VREG_20_5 ) : ( n17669 ) ;
assign n17671 =  ( n17018 ) ? ( VREG_20_6 ) : ( n17670 ) ;
assign n17672 =  ( n17017 ) ? ( VREG_20_7 ) : ( n17671 ) ;
assign n17673 =  ( n17016 ) ? ( VREG_20_8 ) : ( n17672 ) ;
assign n17674 =  ( n17015 ) ? ( VREG_20_9 ) : ( n17673 ) ;
assign n17675 =  ( n17014 ) ? ( VREG_20_10 ) : ( n17674 ) ;
assign n17676 =  ( n17013 ) ? ( VREG_20_11 ) : ( n17675 ) ;
assign n17677 =  ( n17012 ) ? ( VREG_20_12 ) : ( n17676 ) ;
assign n17678 =  ( n17011 ) ? ( VREG_20_13 ) : ( n17677 ) ;
assign n17679 =  ( n17010 ) ? ( VREG_20_14 ) : ( n17678 ) ;
assign n17680 =  ( n17009 ) ? ( VREG_20_15 ) : ( n17679 ) ;
assign n17681 =  ( n17008 ) ? ( VREG_21_0 ) : ( n17680 ) ;
assign n17682 =  ( n17007 ) ? ( VREG_21_1 ) : ( n17681 ) ;
assign n17683 =  ( n17006 ) ? ( VREG_21_2 ) : ( n17682 ) ;
assign n17684 =  ( n17005 ) ? ( VREG_21_3 ) : ( n17683 ) ;
assign n17685 =  ( n17004 ) ? ( VREG_21_4 ) : ( n17684 ) ;
assign n17686 =  ( n17003 ) ? ( VREG_21_5 ) : ( n17685 ) ;
assign n17687 =  ( n17002 ) ? ( VREG_21_6 ) : ( n17686 ) ;
assign n17688 =  ( n17001 ) ? ( VREG_21_7 ) : ( n17687 ) ;
assign n17689 =  ( n17000 ) ? ( VREG_21_8 ) : ( n17688 ) ;
assign n17690 =  ( n16999 ) ? ( VREG_21_9 ) : ( n17689 ) ;
assign n17691 =  ( n16998 ) ? ( VREG_21_10 ) : ( n17690 ) ;
assign n17692 =  ( n16997 ) ? ( VREG_21_11 ) : ( n17691 ) ;
assign n17693 =  ( n16996 ) ? ( VREG_21_12 ) : ( n17692 ) ;
assign n17694 =  ( n16995 ) ? ( VREG_21_13 ) : ( n17693 ) ;
assign n17695 =  ( n16994 ) ? ( VREG_21_14 ) : ( n17694 ) ;
assign n17696 =  ( n16993 ) ? ( VREG_21_15 ) : ( n17695 ) ;
assign n17697 =  ( n16992 ) ? ( VREG_22_0 ) : ( n17696 ) ;
assign n17698 =  ( n16991 ) ? ( VREG_22_1 ) : ( n17697 ) ;
assign n17699 =  ( n16990 ) ? ( VREG_22_2 ) : ( n17698 ) ;
assign n17700 =  ( n16989 ) ? ( VREG_22_3 ) : ( n17699 ) ;
assign n17701 =  ( n16988 ) ? ( VREG_22_4 ) : ( n17700 ) ;
assign n17702 =  ( n16987 ) ? ( VREG_22_5 ) : ( n17701 ) ;
assign n17703 =  ( n16986 ) ? ( VREG_22_6 ) : ( n17702 ) ;
assign n17704 =  ( n16985 ) ? ( VREG_22_7 ) : ( n17703 ) ;
assign n17705 =  ( n16984 ) ? ( VREG_22_8 ) : ( n17704 ) ;
assign n17706 =  ( n16983 ) ? ( VREG_22_9 ) : ( n17705 ) ;
assign n17707 =  ( n16982 ) ? ( VREG_22_10 ) : ( n17706 ) ;
assign n17708 =  ( n16981 ) ? ( VREG_22_11 ) : ( n17707 ) ;
assign n17709 =  ( n16980 ) ? ( VREG_22_12 ) : ( n17708 ) ;
assign n17710 =  ( n16979 ) ? ( VREG_22_13 ) : ( n17709 ) ;
assign n17711 =  ( n16978 ) ? ( VREG_22_14 ) : ( n17710 ) ;
assign n17712 =  ( n16977 ) ? ( VREG_22_15 ) : ( n17711 ) ;
assign n17713 =  ( n16976 ) ? ( VREG_23_0 ) : ( n17712 ) ;
assign n17714 =  ( n16975 ) ? ( VREG_23_1 ) : ( n17713 ) ;
assign n17715 =  ( n16974 ) ? ( VREG_23_2 ) : ( n17714 ) ;
assign n17716 =  ( n16973 ) ? ( VREG_23_3 ) : ( n17715 ) ;
assign n17717 =  ( n16972 ) ? ( VREG_23_4 ) : ( n17716 ) ;
assign n17718 =  ( n16971 ) ? ( VREG_23_5 ) : ( n17717 ) ;
assign n17719 =  ( n16970 ) ? ( VREG_23_6 ) : ( n17718 ) ;
assign n17720 =  ( n16969 ) ? ( VREG_23_7 ) : ( n17719 ) ;
assign n17721 =  ( n16968 ) ? ( VREG_23_8 ) : ( n17720 ) ;
assign n17722 =  ( n16967 ) ? ( VREG_23_9 ) : ( n17721 ) ;
assign n17723 =  ( n16966 ) ? ( VREG_23_10 ) : ( n17722 ) ;
assign n17724 =  ( n16965 ) ? ( VREG_23_11 ) : ( n17723 ) ;
assign n17725 =  ( n16964 ) ? ( VREG_23_12 ) : ( n17724 ) ;
assign n17726 =  ( n16963 ) ? ( VREG_23_13 ) : ( n17725 ) ;
assign n17727 =  ( n16962 ) ? ( VREG_23_14 ) : ( n17726 ) ;
assign n17728 =  ( n16961 ) ? ( VREG_23_15 ) : ( n17727 ) ;
assign n17729 =  ( n16960 ) ? ( VREG_24_0 ) : ( n17728 ) ;
assign n17730 =  ( n16959 ) ? ( VREG_24_1 ) : ( n17729 ) ;
assign n17731 =  ( n16958 ) ? ( VREG_24_2 ) : ( n17730 ) ;
assign n17732 =  ( n16957 ) ? ( VREG_24_3 ) : ( n17731 ) ;
assign n17733 =  ( n16956 ) ? ( VREG_24_4 ) : ( n17732 ) ;
assign n17734 =  ( n16955 ) ? ( VREG_24_5 ) : ( n17733 ) ;
assign n17735 =  ( n16954 ) ? ( VREG_24_6 ) : ( n17734 ) ;
assign n17736 =  ( n16953 ) ? ( VREG_24_7 ) : ( n17735 ) ;
assign n17737 =  ( n16952 ) ? ( VREG_24_8 ) : ( n17736 ) ;
assign n17738 =  ( n16951 ) ? ( VREG_24_9 ) : ( n17737 ) ;
assign n17739 =  ( n16950 ) ? ( VREG_24_10 ) : ( n17738 ) ;
assign n17740 =  ( n16949 ) ? ( VREG_24_11 ) : ( n17739 ) ;
assign n17741 =  ( n16948 ) ? ( VREG_24_12 ) : ( n17740 ) ;
assign n17742 =  ( n16947 ) ? ( VREG_24_13 ) : ( n17741 ) ;
assign n17743 =  ( n16946 ) ? ( VREG_24_14 ) : ( n17742 ) ;
assign n17744 =  ( n16945 ) ? ( VREG_24_15 ) : ( n17743 ) ;
assign n17745 =  ( n16944 ) ? ( VREG_25_0 ) : ( n17744 ) ;
assign n17746 =  ( n16943 ) ? ( VREG_25_1 ) : ( n17745 ) ;
assign n17747 =  ( n16942 ) ? ( VREG_25_2 ) : ( n17746 ) ;
assign n17748 =  ( n16941 ) ? ( VREG_25_3 ) : ( n17747 ) ;
assign n17749 =  ( n16940 ) ? ( VREG_25_4 ) : ( n17748 ) ;
assign n17750 =  ( n16939 ) ? ( VREG_25_5 ) : ( n17749 ) ;
assign n17751 =  ( n16938 ) ? ( VREG_25_6 ) : ( n17750 ) ;
assign n17752 =  ( n16937 ) ? ( VREG_25_7 ) : ( n17751 ) ;
assign n17753 =  ( n16936 ) ? ( VREG_25_8 ) : ( n17752 ) ;
assign n17754 =  ( n16935 ) ? ( VREG_25_9 ) : ( n17753 ) ;
assign n17755 =  ( n16934 ) ? ( VREG_25_10 ) : ( n17754 ) ;
assign n17756 =  ( n16933 ) ? ( VREG_25_11 ) : ( n17755 ) ;
assign n17757 =  ( n16932 ) ? ( VREG_25_12 ) : ( n17756 ) ;
assign n17758 =  ( n16931 ) ? ( VREG_25_13 ) : ( n17757 ) ;
assign n17759 =  ( n16930 ) ? ( VREG_25_14 ) : ( n17758 ) ;
assign n17760 =  ( n16929 ) ? ( VREG_25_15 ) : ( n17759 ) ;
assign n17761 =  ( n16928 ) ? ( VREG_26_0 ) : ( n17760 ) ;
assign n17762 =  ( n16927 ) ? ( VREG_26_1 ) : ( n17761 ) ;
assign n17763 =  ( n16926 ) ? ( VREG_26_2 ) : ( n17762 ) ;
assign n17764 =  ( n16925 ) ? ( VREG_26_3 ) : ( n17763 ) ;
assign n17765 =  ( n16924 ) ? ( VREG_26_4 ) : ( n17764 ) ;
assign n17766 =  ( n16923 ) ? ( VREG_26_5 ) : ( n17765 ) ;
assign n17767 =  ( n16922 ) ? ( VREG_26_6 ) : ( n17766 ) ;
assign n17768 =  ( n16921 ) ? ( VREG_26_7 ) : ( n17767 ) ;
assign n17769 =  ( n16920 ) ? ( VREG_26_8 ) : ( n17768 ) ;
assign n17770 =  ( n16919 ) ? ( VREG_26_9 ) : ( n17769 ) ;
assign n17771 =  ( n16918 ) ? ( VREG_26_10 ) : ( n17770 ) ;
assign n17772 =  ( n16917 ) ? ( VREG_26_11 ) : ( n17771 ) ;
assign n17773 =  ( n16916 ) ? ( VREG_26_12 ) : ( n17772 ) ;
assign n17774 =  ( n16915 ) ? ( VREG_26_13 ) : ( n17773 ) ;
assign n17775 =  ( n16914 ) ? ( VREG_26_14 ) : ( n17774 ) ;
assign n17776 =  ( n16913 ) ? ( VREG_26_15 ) : ( n17775 ) ;
assign n17777 =  ( n16912 ) ? ( VREG_27_0 ) : ( n17776 ) ;
assign n17778 =  ( n16911 ) ? ( VREG_27_1 ) : ( n17777 ) ;
assign n17779 =  ( n16910 ) ? ( VREG_27_2 ) : ( n17778 ) ;
assign n17780 =  ( n16909 ) ? ( VREG_27_3 ) : ( n17779 ) ;
assign n17781 =  ( n16908 ) ? ( VREG_27_4 ) : ( n17780 ) ;
assign n17782 =  ( n16907 ) ? ( VREG_27_5 ) : ( n17781 ) ;
assign n17783 =  ( n16906 ) ? ( VREG_27_6 ) : ( n17782 ) ;
assign n17784 =  ( n16905 ) ? ( VREG_27_7 ) : ( n17783 ) ;
assign n17785 =  ( n16904 ) ? ( VREG_27_8 ) : ( n17784 ) ;
assign n17786 =  ( n16903 ) ? ( VREG_27_9 ) : ( n17785 ) ;
assign n17787 =  ( n16902 ) ? ( VREG_27_10 ) : ( n17786 ) ;
assign n17788 =  ( n16901 ) ? ( VREG_27_11 ) : ( n17787 ) ;
assign n17789 =  ( n16900 ) ? ( VREG_27_12 ) : ( n17788 ) ;
assign n17790 =  ( n16899 ) ? ( VREG_27_13 ) : ( n17789 ) ;
assign n17791 =  ( n16898 ) ? ( VREG_27_14 ) : ( n17790 ) ;
assign n17792 =  ( n16897 ) ? ( VREG_27_15 ) : ( n17791 ) ;
assign n17793 =  ( n16896 ) ? ( VREG_28_0 ) : ( n17792 ) ;
assign n17794 =  ( n16895 ) ? ( VREG_28_1 ) : ( n17793 ) ;
assign n17795 =  ( n16894 ) ? ( VREG_28_2 ) : ( n17794 ) ;
assign n17796 =  ( n16893 ) ? ( VREG_28_3 ) : ( n17795 ) ;
assign n17797 =  ( n16892 ) ? ( VREG_28_4 ) : ( n17796 ) ;
assign n17798 =  ( n16891 ) ? ( VREG_28_5 ) : ( n17797 ) ;
assign n17799 =  ( n16890 ) ? ( VREG_28_6 ) : ( n17798 ) ;
assign n17800 =  ( n16889 ) ? ( VREG_28_7 ) : ( n17799 ) ;
assign n17801 =  ( n16888 ) ? ( VREG_28_8 ) : ( n17800 ) ;
assign n17802 =  ( n16887 ) ? ( VREG_28_9 ) : ( n17801 ) ;
assign n17803 =  ( n16886 ) ? ( VREG_28_10 ) : ( n17802 ) ;
assign n17804 =  ( n16885 ) ? ( VREG_28_11 ) : ( n17803 ) ;
assign n17805 =  ( n16884 ) ? ( VREG_28_12 ) : ( n17804 ) ;
assign n17806 =  ( n16883 ) ? ( VREG_28_13 ) : ( n17805 ) ;
assign n17807 =  ( n16882 ) ? ( VREG_28_14 ) : ( n17806 ) ;
assign n17808 =  ( n16881 ) ? ( VREG_28_15 ) : ( n17807 ) ;
assign n17809 =  ( n16880 ) ? ( VREG_29_0 ) : ( n17808 ) ;
assign n17810 =  ( n16879 ) ? ( VREG_29_1 ) : ( n17809 ) ;
assign n17811 =  ( n16878 ) ? ( VREG_29_2 ) : ( n17810 ) ;
assign n17812 =  ( n16877 ) ? ( VREG_29_3 ) : ( n17811 ) ;
assign n17813 =  ( n16876 ) ? ( VREG_29_4 ) : ( n17812 ) ;
assign n17814 =  ( n16875 ) ? ( VREG_29_5 ) : ( n17813 ) ;
assign n17815 =  ( n16874 ) ? ( VREG_29_6 ) : ( n17814 ) ;
assign n17816 =  ( n16873 ) ? ( VREG_29_7 ) : ( n17815 ) ;
assign n17817 =  ( n16872 ) ? ( VREG_29_8 ) : ( n17816 ) ;
assign n17818 =  ( n16871 ) ? ( VREG_29_9 ) : ( n17817 ) ;
assign n17819 =  ( n16870 ) ? ( VREG_29_10 ) : ( n17818 ) ;
assign n17820 =  ( n16869 ) ? ( VREG_29_11 ) : ( n17819 ) ;
assign n17821 =  ( n16868 ) ? ( VREG_29_12 ) : ( n17820 ) ;
assign n17822 =  ( n16867 ) ? ( VREG_29_13 ) : ( n17821 ) ;
assign n17823 =  ( n16866 ) ? ( VREG_29_14 ) : ( n17822 ) ;
assign n17824 =  ( n16865 ) ? ( VREG_29_15 ) : ( n17823 ) ;
assign n17825 =  ( n16864 ) ? ( VREG_30_0 ) : ( n17824 ) ;
assign n17826 =  ( n16863 ) ? ( VREG_30_1 ) : ( n17825 ) ;
assign n17827 =  ( n16862 ) ? ( VREG_30_2 ) : ( n17826 ) ;
assign n17828 =  ( n16861 ) ? ( VREG_30_3 ) : ( n17827 ) ;
assign n17829 =  ( n16860 ) ? ( VREG_30_4 ) : ( n17828 ) ;
assign n17830 =  ( n16859 ) ? ( VREG_30_5 ) : ( n17829 ) ;
assign n17831 =  ( n16858 ) ? ( VREG_30_6 ) : ( n17830 ) ;
assign n17832 =  ( n16857 ) ? ( VREG_30_7 ) : ( n17831 ) ;
assign n17833 =  ( n16856 ) ? ( VREG_30_8 ) : ( n17832 ) ;
assign n17834 =  ( n16855 ) ? ( VREG_30_9 ) : ( n17833 ) ;
assign n17835 =  ( n16854 ) ? ( VREG_30_10 ) : ( n17834 ) ;
assign n17836 =  ( n16853 ) ? ( VREG_30_11 ) : ( n17835 ) ;
assign n17837 =  ( n16852 ) ? ( VREG_30_12 ) : ( n17836 ) ;
assign n17838 =  ( n16851 ) ? ( VREG_30_13 ) : ( n17837 ) ;
assign n17839 =  ( n16850 ) ? ( VREG_30_14 ) : ( n17838 ) ;
assign n17840 =  ( n16849 ) ? ( VREG_30_15 ) : ( n17839 ) ;
assign n17841 =  ( n16848 ) ? ( VREG_31_0 ) : ( n17840 ) ;
assign n17842 =  ( n16847 ) ? ( VREG_31_1 ) : ( n17841 ) ;
assign n17843 =  ( n16846 ) ? ( VREG_31_2 ) : ( n17842 ) ;
assign n17844 =  ( n16845 ) ? ( VREG_31_3 ) : ( n17843 ) ;
assign n17845 =  ( n16844 ) ? ( VREG_31_4 ) : ( n17844 ) ;
assign n17846 =  ( n16843 ) ? ( VREG_31_5 ) : ( n17845 ) ;
assign n17847 =  ( n16842 ) ? ( VREG_31_6 ) : ( n17846 ) ;
assign n17848 =  ( n16841 ) ? ( VREG_31_7 ) : ( n17847 ) ;
assign n17849 =  ( n16840 ) ? ( VREG_31_8 ) : ( n17848 ) ;
assign n17850 =  ( n16839 ) ? ( VREG_31_9 ) : ( n17849 ) ;
assign n17851 =  ( n16838 ) ? ( VREG_31_10 ) : ( n17850 ) ;
assign n17852 =  ( n16837 ) ? ( VREG_31_11 ) : ( n17851 ) ;
assign n17853 =  ( n16836 ) ? ( VREG_31_12 ) : ( n17852 ) ;
assign n17854 =  ( n16835 ) ? ( VREG_31_13 ) : ( n17853 ) ;
assign n17855 =  ( n16834 ) ? ( VREG_31_14 ) : ( n17854 ) ;
assign n17856 =  ( n16833 ) ? ( VREG_31_15 ) : ( n17855 ) ;
assign n17857 =  ( n16822 ) + ( n17856 )  ;
assign n17858 =  ( n16822 ) - ( n17856 )  ;
assign n17859 =  ( n16822 ) & ( n17856 )  ;
assign n17860 =  ( n16822 ) | ( n17856 )  ;
assign n17861 =  ( ( n16822 ) * ( n17856 ))  ;
assign n17862 =  ( n148 ) ? ( n17861 ) : ( VREG_0_15 ) ;
assign n17863 =  ( n146 ) ? ( n17860 ) : ( n17862 ) ;
assign n17864 =  ( n144 ) ? ( n17859 ) : ( n17863 ) ;
assign n17865 =  ( n142 ) ? ( n17858 ) : ( n17864 ) ;
assign n17866 =  ( n10 ) ? ( n17857 ) : ( n17865 ) ;
assign n17867 = n3030[15:15] ;
assign n17868 =  ( n17867 ) == ( 1'd0 )  ;
assign n17869 =  ( n17868 ) ? ( VREG_0_15 ) : ( n16832 ) ;
assign n17870 =  ( n17868 ) ? ( VREG_0_15 ) : ( n17866 ) ;
assign n17871 =  ( n3034 ) ? ( n17870 ) : ( VREG_0_15 ) ;
assign n17872 =  ( n2965 ) ? ( n17869 ) : ( n17871 ) ;
assign n17873 =  ( n1930 ) ? ( n17866 ) : ( n17872 ) ;
assign n17874 =  ( n879 ) ? ( n16832 ) : ( n17873 ) ;
assign n17875 =  ( n16822 ) + ( n164 )  ;
assign n17876 =  ( n16822 ) - ( n164 )  ;
assign n17877 =  ( n16822 ) & ( n164 )  ;
assign n17878 =  ( n16822 ) | ( n164 )  ;
assign n17879 =  ( ( n16822 ) * ( n164 ))  ;
assign n17880 =  ( n172 ) ? ( n17879 ) : ( VREG_0_15 ) ;
assign n17881 =  ( n170 ) ? ( n17878 ) : ( n17880 ) ;
assign n17882 =  ( n168 ) ? ( n17877 ) : ( n17881 ) ;
assign n17883 =  ( n166 ) ? ( n17876 ) : ( n17882 ) ;
assign n17884 =  ( n162 ) ? ( n17875 ) : ( n17883 ) ;
assign n17885 =  ( n16822 ) + ( n180 )  ;
assign n17886 =  ( n16822 ) - ( n180 )  ;
assign n17887 =  ( n16822 ) & ( n180 )  ;
assign n17888 =  ( n16822 ) | ( n180 )  ;
assign n17889 =  ( ( n16822 ) * ( n180 ))  ;
assign n17890 =  ( n172 ) ? ( n17889 ) : ( VREG_0_15 ) ;
assign n17891 =  ( n170 ) ? ( n17888 ) : ( n17890 ) ;
assign n17892 =  ( n168 ) ? ( n17887 ) : ( n17891 ) ;
assign n17893 =  ( n166 ) ? ( n17886 ) : ( n17892 ) ;
assign n17894 =  ( n162 ) ? ( n17885 ) : ( n17893 ) ;
assign n17895 =  ( n17868 ) ? ( VREG_0_15 ) : ( n17894 ) ;
assign n17896 =  ( n3051 ) ? ( n17895 ) : ( VREG_0_15 ) ;
assign n17897 =  ( n3040 ) ? ( n17884 ) : ( n17896 ) ;
assign n17898 =  ( n192 ) ? ( VREG_0_15 ) : ( VREG_0_15 ) ;
assign n17899 =  ( n157 ) ? ( n17897 ) : ( n17898 ) ;
assign n17900 =  ( n6 ) ? ( n17874 ) : ( n17899 ) ;
assign n17901 =  ( n4 ) ? ( n17900 ) : ( VREG_0_15 ) ;
assign n17902 =  ( 32'd2 ) == ( 32'd15 )  ;
assign n17903 =  ( n12 ) & ( n17902 )  ;
assign n17904 =  ( 32'd2 ) == ( 32'd14 )  ;
assign n17905 =  ( n12 ) & ( n17904 )  ;
assign n17906 =  ( 32'd2 ) == ( 32'd13 )  ;
assign n17907 =  ( n12 ) & ( n17906 )  ;
assign n17908 =  ( 32'd2 ) == ( 32'd12 )  ;
assign n17909 =  ( n12 ) & ( n17908 )  ;
assign n17910 =  ( 32'd2 ) == ( 32'd11 )  ;
assign n17911 =  ( n12 ) & ( n17910 )  ;
assign n17912 =  ( 32'd2 ) == ( 32'd10 )  ;
assign n17913 =  ( n12 ) & ( n17912 )  ;
assign n17914 =  ( 32'd2 ) == ( 32'd9 )  ;
assign n17915 =  ( n12 ) & ( n17914 )  ;
assign n17916 =  ( 32'd2 ) == ( 32'd8 )  ;
assign n17917 =  ( n12 ) & ( n17916 )  ;
assign n17918 =  ( 32'd2 ) == ( 32'd7 )  ;
assign n17919 =  ( n12 ) & ( n17918 )  ;
assign n17920 =  ( 32'd2 ) == ( 32'd6 )  ;
assign n17921 =  ( n12 ) & ( n17920 )  ;
assign n17922 =  ( 32'd2 ) == ( 32'd5 )  ;
assign n17923 =  ( n12 ) & ( n17922 )  ;
assign n17924 =  ( 32'd2 ) == ( 32'd4 )  ;
assign n17925 =  ( n12 ) & ( n17924 )  ;
assign n17926 =  ( 32'd2 ) == ( 32'd3 )  ;
assign n17927 =  ( n12 ) & ( n17926 )  ;
assign n17928 =  ( 32'd2 ) == ( 32'd2 )  ;
assign n17929 =  ( n12 ) & ( n17928 )  ;
assign n17930 =  ( 32'd2 ) == ( 32'd1 )  ;
assign n17931 =  ( n12 ) & ( n17930 )  ;
assign n17932 =  ( 32'd2 ) == ( 32'd0 )  ;
assign n17933 =  ( n12 ) & ( n17932 )  ;
assign n17934 =  ( n13 ) & ( n17902 )  ;
assign n17935 =  ( n13 ) & ( n17904 )  ;
assign n17936 =  ( n13 ) & ( n17906 )  ;
assign n17937 =  ( n13 ) & ( n17908 )  ;
assign n17938 =  ( n13 ) & ( n17910 )  ;
assign n17939 =  ( n13 ) & ( n17912 )  ;
assign n17940 =  ( n13 ) & ( n17914 )  ;
assign n17941 =  ( n13 ) & ( n17916 )  ;
assign n17942 =  ( n13 ) & ( n17918 )  ;
assign n17943 =  ( n13 ) & ( n17920 )  ;
assign n17944 =  ( n13 ) & ( n17922 )  ;
assign n17945 =  ( n13 ) & ( n17924 )  ;
assign n17946 =  ( n13 ) & ( n17926 )  ;
assign n17947 =  ( n13 ) & ( n17928 )  ;
assign n17948 =  ( n13 ) & ( n17930 )  ;
assign n17949 =  ( n13 ) & ( n17932 )  ;
assign n17950 =  ( n14 ) & ( n17902 )  ;
assign n17951 =  ( n14 ) & ( n17904 )  ;
assign n17952 =  ( n14 ) & ( n17906 )  ;
assign n17953 =  ( n14 ) & ( n17908 )  ;
assign n17954 =  ( n14 ) & ( n17910 )  ;
assign n17955 =  ( n14 ) & ( n17912 )  ;
assign n17956 =  ( n14 ) & ( n17914 )  ;
assign n17957 =  ( n14 ) & ( n17916 )  ;
assign n17958 =  ( n14 ) & ( n17918 )  ;
assign n17959 =  ( n14 ) & ( n17920 )  ;
assign n17960 =  ( n14 ) & ( n17922 )  ;
assign n17961 =  ( n14 ) & ( n17924 )  ;
assign n17962 =  ( n14 ) & ( n17926 )  ;
assign n17963 =  ( n14 ) & ( n17928 )  ;
assign n17964 =  ( n14 ) & ( n17930 )  ;
assign n17965 =  ( n14 ) & ( n17932 )  ;
assign n17966 =  ( n15 ) & ( n17902 )  ;
assign n17967 =  ( n15 ) & ( n17904 )  ;
assign n17968 =  ( n15 ) & ( n17906 )  ;
assign n17969 =  ( n15 ) & ( n17908 )  ;
assign n17970 =  ( n15 ) & ( n17910 )  ;
assign n17971 =  ( n15 ) & ( n17912 )  ;
assign n17972 =  ( n15 ) & ( n17914 )  ;
assign n17973 =  ( n15 ) & ( n17916 )  ;
assign n17974 =  ( n15 ) & ( n17918 )  ;
assign n17975 =  ( n15 ) & ( n17920 )  ;
assign n17976 =  ( n15 ) & ( n17922 )  ;
assign n17977 =  ( n15 ) & ( n17924 )  ;
assign n17978 =  ( n15 ) & ( n17926 )  ;
assign n17979 =  ( n15 ) & ( n17928 )  ;
assign n17980 =  ( n15 ) & ( n17930 )  ;
assign n17981 =  ( n15 ) & ( n17932 )  ;
assign n17982 =  ( n16 ) & ( n17902 )  ;
assign n17983 =  ( n16 ) & ( n17904 )  ;
assign n17984 =  ( n16 ) & ( n17906 )  ;
assign n17985 =  ( n16 ) & ( n17908 )  ;
assign n17986 =  ( n16 ) & ( n17910 )  ;
assign n17987 =  ( n16 ) & ( n17912 )  ;
assign n17988 =  ( n16 ) & ( n17914 )  ;
assign n17989 =  ( n16 ) & ( n17916 )  ;
assign n17990 =  ( n16 ) & ( n17918 )  ;
assign n17991 =  ( n16 ) & ( n17920 )  ;
assign n17992 =  ( n16 ) & ( n17922 )  ;
assign n17993 =  ( n16 ) & ( n17924 )  ;
assign n17994 =  ( n16 ) & ( n17926 )  ;
assign n17995 =  ( n16 ) & ( n17928 )  ;
assign n17996 =  ( n16 ) & ( n17930 )  ;
assign n17997 =  ( n16 ) & ( n17932 )  ;
assign n17998 =  ( n17 ) & ( n17902 )  ;
assign n17999 =  ( n17 ) & ( n17904 )  ;
assign n18000 =  ( n17 ) & ( n17906 )  ;
assign n18001 =  ( n17 ) & ( n17908 )  ;
assign n18002 =  ( n17 ) & ( n17910 )  ;
assign n18003 =  ( n17 ) & ( n17912 )  ;
assign n18004 =  ( n17 ) & ( n17914 )  ;
assign n18005 =  ( n17 ) & ( n17916 )  ;
assign n18006 =  ( n17 ) & ( n17918 )  ;
assign n18007 =  ( n17 ) & ( n17920 )  ;
assign n18008 =  ( n17 ) & ( n17922 )  ;
assign n18009 =  ( n17 ) & ( n17924 )  ;
assign n18010 =  ( n17 ) & ( n17926 )  ;
assign n18011 =  ( n17 ) & ( n17928 )  ;
assign n18012 =  ( n17 ) & ( n17930 )  ;
assign n18013 =  ( n17 ) & ( n17932 )  ;
assign n18014 =  ( n18 ) & ( n17902 )  ;
assign n18015 =  ( n18 ) & ( n17904 )  ;
assign n18016 =  ( n18 ) & ( n17906 )  ;
assign n18017 =  ( n18 ) & ( n17908 )  ;
assign n18018 =  ( n18 ) & ( n17910 )  ;
assign n18019 =  ( n18 ) & ( n17912 )  ;
assign n18020 =  ( n18 ) & ( n17914 )  ;
assign n18021 =  ( n18 ) & ( n17916 )  ;
assign n18022 =  ( n18 ) & ( n17918 )  ;
assign n18023 =  ( n18 ) & ( n17920 )  ;
assign n18024 =  ( n18 ) & ( n17922 )  ;
assign n18025 =  ( n18 ) & ( n17924 )  ;
assign n18026 =  ( n18 ) & ( n17926 )  ;
assign n18027 =  ( n18 ) & ( n17928 )  ;
assign n18028 =  ( n18 ) & ( n17930 )  ;
assign n18029 =  ( n18 ) & ( n17932 )  ;
assign n18030 =  ( n19 ) & ( n17902 )  ;
assign n18031 =  ( n19 ) & ( n17904 )  ;
assign n18032 =  ( n19 ) & ( n17906 )  ;
assign n18033 =  ( n19 ) & ( n17908 )  ;
assign n18034 =  ( n19 ) & ( n17910 )  ;
assign n18035 =  ( n19 ) & ( n17912 )  ;
assign n18036 =  ( n19 ) & ( n17914 )  ;
assign n18037 =  ( n19 ) & ( n17916 )  ;
assign n18038 =  ( n19 ) & ( n17918 )  ;
assign n18039 =  ( n19 ) & ( n17920 )  ;
assign n18040 =  ( n19 ) & ( n17922 )  ;
assign n18041 =  ( n19 ) & ( n17924 )  ;
assign n18042 =  ( n19 ) & ( n17926 )  ;
assign n18043 =  ( n19 ) & ( n17928 )  ;
assign n18044 =  ( n19 ) & ( n17930 )  ;
assign n18045 =  ( n19 ) & ( n17932 )  ;
assign n18046 =  ( n20 ) & ( n17902 )  ;
assign n18047 =  ( n20 ) & ( n17904 )  ;
assign n18048 =  ( n20 ) & ( n17906 )  ;
assign n18049 =  ( n20 ) & ( n17908 )  ;
assign n18050 =  ( n20 ) & ( n17910 )  ;
assign n18051 =  ( n20 ) & ( n17912 )  ;
assign n18052 =  ( n20 ) & ( n17914 )  ;
assign n18053 =  ( n20 ) & ( n17916 )  ;
assign n18054 =  ( n20 ) & ( n17918 )  ;
assign n18055 =  ( n20 ) & ( n17920 )  ;
assign n18056 =  ( n20 ) & ( n17922 )  ;
assign n18057 =  ( n20 ) & ( n17924 )  ;
assign n18058 =  ( n20 ) & ( n17926 )  ;
assign n18059 =  ( n20 ) & ( n17928 )  ;
assign n18060 =  ( n20 ) & ( n17930 )  ;
assign n18061 =  ( n20 ) & ( n17932 )  ;
assign n18062 =  ( n21 ) & ( n17902 )  ;
assign n18063 =  ( n21 ) & ( n17904 )  ;
assign n18064 =  ( n21 ) & ( n17906 )  ;
assign n18065 =  ( n21 ) & ( n17908 )  ;
assign n18066 =  ( n21 ) & ( n17910 )  ;
assign n18067 =  ( n21 ) & ( n17912 )  ;
assign n18068 =  ( n21 ) & ( n17914 )  ;
assign n18069 =  ( n21 ) & ( n17916 )  ;
assign n18070 =  ( n21 ) & ( n17918 )  ;
assign n18071 =  ( n21 ) & ( n17920 )  ;
assign n18072 =  ( n21 ) & ( n17922 )  ;
assign n18073 =  ( n21 ) & ( n17924 )  ;
assign n18074 =  ( n21 ) & ( n17926 )  ;
assign n18075 =  ( n21 ) & ( n17928 )  ;
assign n18076 =  ( n21 ) & ( n17930 )  ;
assign n18077 =  ( n21 ) & ( n17932 )  ;
assign n18078 =  ( n22 ) & ( n17902 )  ;
assign n18079 =  ( n22 ) & ( n17904 )  ;
assign n18080 =  ( n22 ) & ( n17906 )  ;
assign n18081 =  ( n22 ) & ( n17908 )  ;
assign n18082 =  ( n22 ) & ( n17910 )  ;
assign n18083 =  ( n22 ) & ( n17912 )  ;
assign n18084 =  ( n22 ) & ( n17914 )  ;
assign n18085 =  ( n22 ) & ( n17916 )  ;
assign n18086 =  ( n22 ) & ( n17918 )  ;
assign n18087 =  ( n22 ) & ( n17920 )  ;
assign n18088 =  ( n22 ) & ( n17922 )  ;
assign n18089 =  ( n22 ) & ( n17924 )  ;
assign n18090 =  ( n22 ) & ( n17926 )  ;
assign n18091 =  ( n22 ) & ( n17928 )  ;
assign n18092 =  ( n22 ) & ( n17930 )  ;
assign n18093 =  ( n22 ) & ( n17932 )  ;
assign n18094 =  ( n23 ) & ( n17902 )  ;
assign n18095 =  ( n23 ) & ( n17904 )  ;
assign n18096 =  ( n23 ) & ( n17906 )  ;
assign n18097 =  ( n23 ) & ( n17908 )  ;
assign n18098 =  ( n23 ) & ( n17910 )  ;
assign n18099 =  ( n23 ) & ( n17912 )  ;
assign n18100 =  ( n23 ) & ( n17914 )  ;
assign n18101 =  ( n23 ) & ( n17916 )  ;
assign n18102 =  ( n23 ) & ( n17918 )  ;
assign n18103 =  ( n23 ) & ( n17920 )  ;
assign n18104 =  ( n23 ) & ( n17922 )  ;
assign n18105 =  ( n23 ) & ( n17924 )  ;
assign n18106 =  ( n23 ) & ( n17926 )  ;
assign n18107 =  ( n23 ) & ( n17928 )  ;
assign n18108 =  ( n23 ) & ( n17930 )  ;
assign n18109 =  ( n23 ) & ( n17932 )  ;
assign n18110 =  ( n24 ) & ( n17902 )  ;
assign n18111 =  ( n24 ) & ( n17904 )  ;
assign n18112 =  ( n24 ) & ( n17906 )  ;
assign n18113 =  ( n24 ) & ( n17908 )  ;
assign n18114 =  ( n24 ) & ( n17910 )  ;
assign n18115 =  ( n24 ) & ( n17912 )  ;
assign n18116 =  ( n24 ) & ( n17914 )  ;
assign n18117 =  ( n24 ) & ( n17916 )  ;
assign n18118 =  ( n24 ) & ( n17918 )  ;
assign n18119 =  ( n24 ) & ( n17920 )  ;
assign n18120 =  ( n24 ) & ( n17922 )  ;
assign n18121 =  ( n24 ) & ( n17924 )  ;
assign n18122 =  ( n24 ) & ( n17926 )  ;
assign n18123 =  ( n24 ) & ( n17928 )  ;
assign n18124 =  ( n24 ) & ( n17930 )  ;
assign n18125 =  ( n24 ) & ( n17932 )  ;
assign n18126 =  ( n25 ) & ( n17902 )  ;
assign n18127 =  ( n25 ) & ( n17904 )  ;
assign n18128 =  ( n25 ) & ( n17906 )  ;
assign n18129 =  ( n25 ) & ( n17908 )  ;
assign n18130 =  ( n25 ) & ( n17910 )  ;
assign n18131 =  ( n25 ) & ( n17912 )  ;
assign n18132 =  ( n25 ) & ( n17914 )  ;
assign n18133 =  ( n25 ) & ( n17916 )  ;
assign n18134 =  ( n25 ) & ( n17918 )  ;
assign n18135 =  ( n25 ) & ( n17920 )  ;
assign n18136 =  ( n25 ) & ( n17922 )  ;
assign n18137 =  ( n25 ) & ( n17924 )  ;
assign n18138 =  ( n25 ) & ( n17926 )  ;
assign n18139 =  ( n25 ) & ( n17928 )  ;
assign n18140 =  ( n25 ) & ( n17930 )  ;
assign n18141 =  ( n25 ) & ( n17932 )  ;
assign n18142 =  ( n26 ) & ( n17902 )  ;
assign n18143 =  ( n26 ) & ( n17904 )  ;
assign n18144 =  ( n26 ) & ( n17906 )  ;
assign n18145 =  ( n26 ) & ( n17908 )  ;
assign n18146 =  ( n26 ) & ( n17910 )  ;
assign n18147 =  ( n26 ) & ( n17912 )  ;
assign n18148 =  ( n26 ) & ( n17914 )  ;
assign n18149 =  ( n26 ) & ( n17916 )  ;
assign n18150 =  ( n26 ) & ( n17918 )  ;
assign n18151 =  ( n26 ) & ( n17920 )  ;
assign n18152 =  ( n26 ) & ( n17922 )  ;
assign n18153 =  ( n26 ) & ( n17924 )  ;
assign n18154 =  ( n26 ) & ( n17926 )  ;
assign n18155 =  ( n26 ) & ( n17928 )  ;
assign n18156 =  ( n26 ) & ( n17930 )  ;
assign n18157 =  ( n26 ) & ( n17932 )  ;
assign n18158 =  ( n27 ) & ( n17902 )  ;
assign n18159 =  ( n27 ) & ( n17904 )  ;
assign n18160 =  ( n27 ) & ( n17906 )  ;
assign n18161 =  ( n27 ) & ( n17908 )  ;
assign n18162 =  ( n27 ) & ( n17910 )  ;
assign n18163 =  ( n27 ) & ( n17912 )  ;
assign n18164 =  ( n27 ) & ( n17914 )  ;
assign n18165 =  ( n27 ) & ( n17916 )  ;
assign n18166 =  ( n27 ) & ( n17918 )  ;
assign n18167 =  ( n27 ) & ( n17920 )  ;
assign n18168 =  ( n27 ) & ( n17922 )  ;
assign n18169 =  ( n27 ) & ( n17924 )  ;
assign n18170 =  ( n27 ) & ( n17926 )  ;
assign n18171 =  ( n27 ) & ( n17928 )  ;
assign n18172 =  ( n27 ) & ( n17930 )  ;
assign n18173 =  ( n27 ) & ( n17932 )  ;
assign n18174 =  ( n28 ) & ( n17902 )  ;
assign n18175 =  ( n28 ) & ( n17904 )  ;
assign n18176 =  ( n28 ) & ( n17906 )  ;
assign n18177 =  ( n28 ) & ( n17908 )  ;
assign n18178 =  ( n28 ) & ( n17910 )  ;
assign n18179 =  ( n28 ) & ( n17912 )  ;
assign n18180 =  ( n28 ) & ( n17914 )  ;
assign n18181 =  ( n28 ) & ( n17916 )  ;
assign n18182 =  ( n28 ) & ( n17918 )  ;
assign n18183 =  ( n28 ) & ( n17920 )  ;
assign n18184 =  ( n28 ) & ( n17922 )  ;
assign n18185 =  ( n28 ) & ( n17924 )  ;
assign n18186 =  ( n28 ) & ( n17926 )  ;
assign n18187 =  ( n28 ) & ( n17928 )  ;
assign n18188 =  ( n28 ) & ( n17930 )  ;
assign n18189 =  ( n28 ) & ( n17932 )  ;
assign n18190 =  ( n29 ) & ( n17902 )  ;
assign n18191 =  ( n29 ) & ( n17904 )  ;
assign n18192 =  ( n29 ) & ( n17906 )  ;
assign n18193 =  ( n29 ) & ( n17908 )  ;
assign n18194 =  ( n29 ) & ( n17910 )  ;
assign n18195 =  ( n29 ) & ( n17912 )  ;
assign n18196 =  ( n29 ) & ( n17914 )  ;
assign n18197 =  ( n29 ) & ( n17916 )  ;
assign n18198 =  ( n29 ) & ( n17918 )  ;
assign n18199 =  ( n29 ) & ( n17920 )  ;
assign n18200 =  ( n29 ) & ( n17922 )  ;
assign n18201 =  ( n29 ) & ( n17924 )  ;
assign n18202 =  ( n29 ) & ( n17926 )  ;
assign n18203 =  ( n29 ) & ( n17928 )  ;
assign n18204 =  ( n29 ) & ( n17930 )  ;
assign n18205 =  ( n29 ) & ( n17932 )  ;
assign n18206 =  ( n30 ) & ( n17902 )  ;
assign n18207 =  ( n30 ) & ( n17904 )  ;
assign n18208 =  ( n30 ) & ( n17906 )  ;
assign n18209 =  ( n30 ) & ( n17908 )  ;
assign n18210 =  ( n30 ) & ( n17910 )  ;
assign n18211 =  ( n30 ) & ( n17912 )  ;
assign n18212 =  ( n30 ) & ( n17914 )  ;
assign n18213 =  ( n30 ) & ( n17916 )  ;
assign n18214 =  ( n30 ) & ( n17918 )  ;
assign n18215 =  ( n30 ) & ( n17920 )  ;
assign n18216 =  ( n30 ) & ( n17922 )  ;
assign n18217 =  ( n30 ) & ( n17924 )  ;
assign n18218 =  ( n30 ) & ( n17926 )  ;
assign n18219 =  ( n30 ) & ( n17928 )  ;
assign n18220 =  ( n30 ) & ( n17930 )  ;
assign n18221 =  ( n30 ) & ( n17932 )  ;
assign n18222 =  ( n31 ) & ( n17902 )  ;
assign n18223 =  ( n31 ) & ( n17904 )  ;
assign n18224 =  ( n31 ) & ( n17906 )  ;
assign n18225 =  ( n31 ) & ( n17908 )  ;
assign n18226 =  ( n31 ) & ( n17910 )  ;
assign n18227 =  ( n31 ) & ( n17912 )  ;
assign n18228 =  ( n31 ) & ( n17914 )  ;
assign n18229 =  ( n31 ) & ( n17916 )  ;
assign n18230 =  ( n31 ) & ( n17918 )  ;
assign n18231 =  ( n31 ) & ( n17920 )  ;
assign n18232 =  ( n31 ) & ( n17922 )  ;
assign n18233 =  ( n31 ) & ( n17924 )  ;
assign n18234 =  ( n31 ) & ( n17926 )  ;
assign n18235 =  ( n31 ) & ( n17928 )  ;
assign n18236 =  ( n31 ) & ( n17930 )  ;
assign n18237 =  ( n31 ) & ( n17932 )  ;
assign n18238 =  ( n32 ) & ( n17902 )  ;
assign n18239 =  ( n32 ) & ( n17904 )  ;
assign n18240 =  ( n32 ) & ( n17906 )  ;
assign n18241 =  ( n32 ) & ( n17908 )  ;
assign n18242 =  ( n32 ) & ( n17910 )  ;
assign n18243 =  ( n32 ) & ( n17912 )  ;
assign n18244 =  ( n32 ) & ( n17914 )  ;
assign n18245 =  ( n32 ) & ( n17916 )  ;
assign n18246 =  ( n32 ) & ( n17918 )  ;
assign n18247 =  ( n32 ) & ( n17920 )  ;
assign n18248 =  ( n32 ) & ( n17922 )  ;
assign n18249 =  ( n32 ) & ( n17924 )  ;
assign n18250 =  ( n32 ) & ( n17926 )  ;
assign n18251 =  ( n32 ) & ( n17928 )  ;
assign n18252 =  ( n32 ) & ( n17930 )  ;
assign n18253 =  ( n32 ) & ( n17932 )  ;
assign n18254 =  ( n33 ) & ( n17902 )  ;
assign n18255 =  ( n33 ) & ( n17904 )  ;
assign n18256 =  ( n33 ) & ( n17906 )  ;
assign n18257 =  ( n33 ) & ( n17908 )  ;
assign n18258 =  ( n33 ) & ( n17910 )  ;
assign n18259 =  ( n33 ) & ( n17912 )  ;
assign n18260 =  ( n33 ) & ( n17914 )  ;
assign n18261 =  ( n33 ) & ( n17916 )  ;
assign n18262 =  ( n33 ) & ( n17918 )  ;
assign n18263 =  ( n33 ) & ( n17920 )  ;
assign n18264 =  ( n33 ) & ( n17922 )  ;
assign n18265 =  ( n33 ) & ( n17924 )  ;
assign n18266 =  ( n33 ) & ( n17926 )  ;
assign n18267 =  ( n33 ) & ( n17928 )  ;
assign n18268 =  ( n33 ) & ( n17930 )  ;
assign n18269 =  ( n33 ) & ( n17932 )  ;
assign n18270 =  ( n34 ) & ( n17902 )  ;
assign n18271 =  ( n34 ) & ( n17904 )  ;
assign n18272 =  ( n34 ) & ( n17906 )  ;
assign n18273 =  ( n34 ) & ( n17908 )  ;
assign n18274 =  ( n34 ) & ( n17910 )  ;
assign n18275 =  ( n34 ) & ( n17912 )  ;
assign n18276 =  ( n34 ) & ( n17914 )  ;
assign n18277 =  ( n34 ) & ( n17916 )  ;
assign n18278 =  ( n34 ) & ( n17918 )  ;
assign n18279 =  ( n34 ) & ( n17920 )  ;
assign n18280 =  ( n34 ) & ( n17922 )  ;
assign n18281 =  ( n34 ) & ( n17924 )  ;
assign n18282 =  ( n34 ) & ( n17926 )  ;
assign n18283 =  ( n34 ) & ( n17928 )  ;
assign n18284 =  ( n34 ) & ( n17930 )  ;
assign n18285 =  ( n34 ) & ( n17932 )  ;
assign n18286 =  ( n35 ) & ( n17902 )  ;
assign n18287 =  ( n35 ) & ( n17904 )  ;
assign n18288 =  ( n35 ) & ( n17906 )  ;
assign n18289 =  ( n35 ) & ( n17908 )  ;
assign n18290 =  ( n35 ) & ( n17910 )  ;
assign n18291 =  ( n35 ) & ( n17912 )  ;
assign n18292 =  ( n35 ) & ( n17914 )  ;
assign n18293 =  ( n35 ) & ( n17916 )  ;
assign n18294 =  ( n35 ) & ( n17918 )  ;
assign n18295 =  ( n35 ) & ( n17920 )  ;
assign n18296 =  ( n35 ) & ( n17922 )  ;
assign n18297 =  ( n35 ) & ( n17924 )  ;
assign n18298 =  ( n35 ) & ( n17926 )  ;
assign n18299 =  ( n35 ) & ( n17928 )  ;
assign n18300 =  ( n35 ) & ( n17930 )  ;
assign n18301 =  ( n35 ) & ( n17932 )  ;
assign n18302 =  ( n36 ) & ( n17902 )  ;
assign n18303 =  ( n36 ) & ( n17904 )  ;
assign n18304 =  ( n36 ) & ( n17906 )  ;
assign n18305 =  ( n36 ) & ( n17908 )  ;
assign n18306 =  ( n36 ) & ( n17910 )  ;
assign n18307 =  ( n36 ) & ( n17912 )  ;
assign n18308 =  ( n36 ) & ( n17914 )  ;
assign n18309 =  ( n36 ) & ( n17916 )  ;
assign n18310 =  ( n36 ) & ( n17918 )  ;
assign n18311 =  ( n36 ) & ( n17920 )  ;
assign n18312 =  ( n36 ) & ( n17922 )  ;
assign n18313 =  ( n36 ) & ( n17924 )  ;
assign n18314 =  ( n36 ) & ( n17926 )  ;
assign n18315 =  ( n36 ) & ( n17928 )  ;
assign n18316 =  ( n36 ) & ( n17930 )  ;
assign n18317 =  ( n36 ) & ( n17932 )  ;
assign n18318 =  ( n37 ) & ( n17902 )  ;
assign n18319 =  ( n37 ) & ( n17904 )  ;
assign n18320 =  ( n37 ) & ( n17906 )  ;
assign n18321 =  ( n37 ) & ( n17908 )  ;
assign n18322 =  ( n37 ) & ( n17910 )  ;
assign n18323 =  ( n37 ) & ( n17912 )  ;
assign n18324 =  ( n37 ) & ( n17914 )  ;
assign n18325 =  ( n37 ) & ( n17916 )  ;
assign n18326 =  ( n37 ) & ( n17918 )  ;
assign n18327 =  ( n37 ) & ( n17920 )  ;
assign n18328 =  ( n37 ) & ( n17922 )  ;
assign n18329 =  ( n37 ) & ( n17924 )  ;
assign n18330 =  ( n37 ) & ( n17926 )  ;
assign n18331 =  ( n37 ) & ( n17928 )  ;
assign n18332 =  ( n37 ) & ( n17930 )  ;
assign n18333 =  ( n37 ) & ( n17932 )  ;
assign n18334 =  ( n38 ) & ( n17902 )  ;
assign n18335 =  ( n38 ) & ( n17904 )  ;
assign n18336 =  ( n38 ) & ( n17906 )  ;
assign n18337 =  ( n38 ) & ( n17908 )  ;
assign n18338 =  ( n38 ) & ( n17910 )  ;
assign n18339 =  ( n38 ) & ( n17912 )  ;
assign n18340 =  ( n38 ) & ( n17914 )  ;
assign n18341 =  ( n38 ) & ( n17916 )  ;
assign n18342 =  ( n38 ) & ( n17918 )  ;
assign n18343 =  ( n38 ) & ( n17920 )  ;
assign n18344 =  ( n38 ) & ( n17922 )  ;
assign n18345 =  ( n38 ) & ( n17924 )  ;
assign n18346 =  ( n38 ) & ( n17926 )  ;
assign n18347 =  ( n38 ) & ( n17928 )  ;
assign n18348 =  ( n38 ) & ( n17930 )  ;
assign n18349 =  ( n38 ) & ( n17932 )  ;
assign n18350 =  ( n39 ) & ( n17902 )  ;
assign n18351 =  ( n39 ) & ( n17904 )  ;
assign n18352 =  ( n39 ) & ( n17906 )  ;
assign n18353 =  ( n39 ) & ( n17908 )  ;
assign n18354 =  ( n39 ) & ( n17910 )  ;
assign n18355 =  ( n39 ) & ( n17912 )  ;
assign n18356 =  ( n39 ) & ( n17914 )  ;
assign n18357 =  ( n39 ) & ( n17916 )  ;
assign n18358 =  ( n39 ) & ( n17918 )  ;
assign n18359 =  ( n39 ) & ( n17920 )  ;
assign n18360 =  ( n39 ) & ( n17922 )  ;
assign n18361 =  ( n39 ) & ( n17924 )  ;
assign n18362 =  ( n39 ) & ( n17926 )  ;
assign n18363 =  ( n39 ) & ( n17928 )  ;
assign n18364 =  ( n39 ) & ( n17930 )  ;
assign n18365 =  ( n39 ) & ( n17932 )  ;
assign n18366 =  ( n40 ) & ( n17902 )  ;
assign n18367 =  ( n40 ) & ( n17904 )  ;
assign n18368 =  ( n40 ) & ( n17906 )  ;
assign n18369 =  ( n40 ) & ( n17908 )  ;
assign n18370 =  ( n40 ) & ( n17910 )  ;
assign n18371 =  ( n40 ) & ( n17912 )  ;
assign n18372 =  ( n40 ) & ( n17914 )  ;
assign n18373 =  ( n40 ) & ( n17916 )  ;
assign n18374 =  ( n40 ) & ( n17918 )  ;
assign n18375 =  ( n40 ) & ( n17920 )  ;
assign n18376 =  ( n40 ) & ( n17922 )  ;
assign n18377 =  ( n40 ) & ( n17924 )  ;
assign n18378 =  ( n40 ) & ( n17926 )  ;
assign n18379 =  ( n40 ) & ( n17928 )  ;
assign n18380 =  ( n40 ) & ( n17930 )  ;
assign n18381 =  ( n40 ) & ( n17932 )  ;
assign n18382 =  ( n41 ) & ( n17902 )  ;
assign n18383 =  ( n41 ) & ( n17904 )  ;
assign n18384 =  ( n41 ) & ( n17906 )  ;
assign n18385 =  ( n41 ) & ( n17908 )  ;
assign n18386 =  ( n41 ) & ( n17910 )  ;
assign n18387 =  ( n41 ) & ( n17912 )  ;
assign n18388 =  ( n41 ) & ( n17914 )  ;
assign n18389 =  ( n41 ) & ( n17916 )  ;
assign n18390 =  ( n41 ) & ( n17918 )  ;
assign n18391 =  ( n41 ) & ( n17920 )  ;
assign n18392 =  ( n41 ) & ( n17922 )  ;
assign n18393 =  ( n41 ) & ( n17924 )  ;
assign n18394 =  ( n41 ) & ( n17926 )  ;
assign n18395 =  ( n41 ) & ( n17928 )  ;
assign n18396 =  ( n41 ) & ( n17930 )  ;
assign n18397 =  ( n41 ) & ( n17932 )  ;
assign n18398 =  ( n42 ) & ( n17902 )  ;
assign n18399 =  ( n42 ) & ( n17904 )  ;
assign n18400 =  ( n42 ) & ( n17906 )  ;
assign n18401 =  ( n42 ) & ( n17908 )  ;
assign n18402 =  ( n42 ) & ( n17910 )  ;
assign n18403 =  ( n42 ) & ( n17912 )  ;
assign n18404 =  ( n42 ) & ( n17914 )  ;
assign n18405 =  ( n42 ) & ( n17916 )  ;
assign n18406 =  ( n42 ) & ( n17918 )  ;
assign n18407 =  ( n42 ) & ( n17920 )  ;
assign n18408 =  ( n42 ) & ( n17922 )  ;
assign n18409 =  ( n42 ) & ( n17924 )  ;
assign n18410 =  ( n42 ) & ( n17926 )  ;
assign n18411 =  ( n42 ) & ( n17928 )  ;
assign n18412 =  ( n42 ) & ( n17930 )  ;
assign n18413 =  ( n42 ) & ( n17932 )  ;
assign n18414 =  ( n43 ) & ( n17902 )  ;
assign n18415 =  ( n43 ) & ( n17904 )  ;
assign n18416 =  ( n43 ) & ( n17906 )  ;
assign n18417 =  ( n43 ) & ( n17908 )  ;
assign n18418 =  ( n43 ) & ( n17910 )  ;
assign n18419 =  ( n43 ) & ( n17912 )  ;
assign n18420 =  ( n43 ) & ( n17914 )  ;
assign n18421 =  ( n43 ) & ( n17916 )  ;
assign n18422 =  ( n43 ) & ( n17918 )  ;
assign n18423 =  ( n43 ) & ( n17920 )  ;
assign n18424 =  ( n43 ) & ( n17922 )  ;
assign n18425 =  ( n43 ) & ( n17924 )  ;
assign n18426 =  ( n43 ) & ( n17926 )  ;
assign n18427 =  ( n43 ) & ( n17928 )  ;
assign n18428 =  ( n43 ) & ( n17930 )  ;
assign n18429 =  ( n43 ) & ( n17932 )  ;
assign n18430 =  ( n18429 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n18431 =  ( n18428 ) ? ( VREG_0_1 ) : ( n18430 ) ;
assign n18432 =  ( n18427 ) ? ( VREG_0_2 ) : ( n18431 ) ;
assign n18433 =  ( n18426 ) ? ( VREG_0_3 ) : ( n18432 ) ;
assign n18434 =  ( n18425 ) ? ( VREG_0_4 ) : ( n18433 ) ;
assign n18435 =  ( n18424 ) ? ( VREG_0_5 ) : ( n18434 ) ;
assign n18436 =  ( n18423 ) ? ( VREG_0_6 ) : ( n18435 ) ;
assign n18437 =  ( n18422 ) ? ( VREG_0_7 ) : ( n18436 ) ;
assign n18438 =  ( n18421 ) ? ( VREG_0_8 ) : ( n18437 ) ;
assign n18439 =  ( n18420 ) ? ( VREG_0_9 ) : ( n18438 ) ;
assign n18440 =  ( n18419 ) ? ( VREG_0_10 ) : ( n18439 ) ;
assign n18441 =  ( n18418 ) ? ( VREG_0_11 ) : ( n18440 ) ;
assign n18442 =  ( n18417 ) ? ( VREG_0_12 ) : ( n18441 ) ;
assign n18443 =  ( n18416 ) ? ( VREG_0_13 ) : ( n18442 ) ;
assign n18444 =  ( n18415 ) ? ( VREG_0_14 ) : ( n18443 ) ;
assign n18445 =  ( n18414 ) ? ( VREG_0_15 ) : ( n18444 ) ;
assign n18446 =  ( n18413 ) ? ( VREG_1_0 ) : ( n18445 ) ;
assign n18447 =  ( n18412 ) ? ( VREG_1_1 ) : ( n18446 ) ;
assign n18448 =  ( n18411 ) ? ( VREG_1_2 ) : ( n18447 ) ;
assign n18449 =  ( n18410 ) ? ( VREG_1_3 ) : ( n18448 ) ;
assign n18450 =  ( n18409 ) ? ( VREG_1_4 ) : ( n18449 ) ;
assign n18451 =  ( n18408 ) ? ( VREG_1_5 ) : ( n18450 ) ;
assign n18452 =  ( n18407 ) ? ( VREG_1_6 ) : ( n18451 ) ;
assign n18453 =  ( n18406 ) ? ( VREG_1_7 ) : ( n18452 ) ;
assign n18454 =  ( n18405 ) ? ( VREG_1_8 ) : ( n18453 ) ;
assign n18455 =  ( n18404 ) ? ( VREG_1_9 ) : ( n18454 ) ;
assign n18456 =  ( n18403 ) ? ( VREG_1_10 ) : ( n18455 ) ;
assign n18457 =  ( n18402 ) ? ( VREG_1_11 ) : ( n18456 ) ;
assign n18458 =  ( n18401 ) ? ( VREG_1_12 ) : ( n18457 ) ;
assign n18459 =  ( n18400 ) ? ( VREG_1_13 ) : ( n18458 ) ;
assign n18460 =  ( n18399 ) ? ( VREG_1_14 ) : ( n18459 ) ;
assign n18461 =  ( n18398 ) ? ( VREG_1_15 ) : ( n18460 ) ;
assign n18462 =  ( n18397 ) ? ( VREG_2_0 ) : ( n18461 ) ;
assign n18463 =  ( n18396 ) ? ( VREG_2_1 ) : ( n18462 ) ;
assign n18464 =  ( n18395 ) ? ( VREG_2_2 ) : ( n18463 ) ;
assign n18465 =  ( n18394 ) ? ( VREG_2_3 ) : ( n18464 ) ;
assign n18466 =  ( n18393 ) ? ( VREG_2_4 ) : ( n18465 ) ;
assign n18467 =  ( n18392 ) ? ( VREG_2_5 ) : ( n18466 ) ;
assign n18468 =  ( n18391 ) ? ( VREG_2_6 ) : ( n18467 ) ;
assign n18469 =  ( n18390 ) ? ( VREG_2_7 ) : ( n18468 ) ;
assign n18470 =  ( n18389 ) ? ( VREG_2_8 ) : ( n18469 ) ;
assign n18471 =  ( n18388 ) ? ( VREG_2_9 ) : ( n18470 ) ;
assign n18472 =  ( n18387 ) ? ( VREG_2_10 ) : ( n18471 ) ;
assign n18473 =  ( n18386 ) ? ( VREG_2_11 ) : ( n18472 ) ;
assign n18474 =  ( n18385 ) ? ( VREG_2_12 ) : ( n18473 ) ;
assign n18475 =  ( n18384 ) ? ( VREG_2_13 ) : ( n18474 ) ;
assign n18476 =  ( n18383 ) ? ( VREG_2_14 ) : ( n18475 ) ;
assign n18477 =  ( n18382 ) ? ( VREG_2_15 ) : ( n18476 ) ;
assign n18478 =  ( n18381 ) ? ( VREG_3_0 ) : ( n18477 ) ;
assign n18479 =  ( n18380 ) ? ( VREG_3_1 ) : ( n18478 ) ;
assign n18480 =  ( n18379 ) ? ( VREG_3_2 ) : ( n18479 ) ;
assign n18481 =  ( n18378 ) ? ( VREG_3_3 ) : ( n18480 ) ;
assign n18482 =  ( n18377 ) ? ( VREG_3_4 ) : ( n18481 ) ;
assign n18483 =  ( n18376 ) ? ( VREG_3_5 ) : ( n18482 ) ;
assign n18484 =  ( n18375 ) ? ( VREG_3_6 ) : ( n18483 ) ;
assign n18485 =  ( n18374 ) ? ( VREG_3_7 ) : ( n18484 ) ;
assign n18486 =  ( n18373 ) ? ( VREG_3_8 ) : ( n18485 ) ;
assign n18487 =  ( n18372 ) ? ( VREG_3_9 ) : ( n18486 ) ;
assign n18488 =  ( n18371 ) ? ( VREG_3_10 ) : ( n18487 ) ;
assign n18489 =  ( n18370 ) ? ( VREG_3_11 ) : ( n18488 ) ;
assign n18490 =  ( n18369 ) ? ( VREG_3_12 ) : ( n18489 ) ;
assign n18491 =  ( n18368 ) ? ( VREG_3_13 ) : ( n18490 ) ;
assign n18492 =  ( n18367 ) ? ( VREG_3_14 ) : ( n18491 ) ;
assign n18493 =  ( n18366 ) ? ( VREG_3_15 ) : ( n18492 ) ;
assign n18494 =  ( n18365 ) ? ( VREG_4_0 ) : ( n18493 ) ;
assign n18495 =  ( n18364 ) ? ( VREG_4_1 ) : ( n18494 ) ;
assign n18496 =  ( n18363 ) ? ( VREG_4_2 ) : ( n18495 ) ;
assign n18497 =  ( n18362 ) ? ( VREG_4_3 ) : ( n18496 ) ;
assign n18498 =  ( n18361 ) ? ( VREG_4_4 ) : ( n18497 ) ;
assign n18499 =  ( n18360 ) ? ( VREG_4_5 ) : ( n18498 ) ;
assign n18500 =  ( n18359 ) ? ( VREG_4_6 ) : ( n18499 ) ;
assign n18501 =  ( n18358 ) ? ( VREG_4_7 ) : ( n18500 ) ;
assign n18502 =  ( n18357 ) ? ( VREG_4_8 ) : ( n18501 ) ;
assign n18503 =  ( n18356 ) ? ( VREG_4_9 ) : ( n18502 ) ;
assign n18504 =  ( n18355 ) ? ( VREG_4_10 ) : ( n18503 ) ;
assign n18505 =  ( n18354 ) ? ( VREG_4_11 ) : ( n18504 ) ;
assign n18506 =  ( n18353 ) ? ( VREG_4_12 ) : ( n18505 ) ;
assign n18507 =  ( n18352 ) ? ( VREG_4_13 ) : ( n18506 ) ;
assign n18508 =  ( n18351 ) ? ( VREG_4_14 ) : ( n18507 ) ;
assign n18509 =  ( n18350 ) ? ( VREG_4_15 ) : ( n18508 ) ;
assign n18510 =  ( n18349 ) ? ( VREG_5_0 ) : ( n18509 ) ;
assign n18511 =  ( n18348 ) ? ( VREG_5_1 ) : ( n18510 ) ;
assign n18512 =  ( n18347 ) ? ( VREG_5_2 ) : ( n18511 ) ;
assign n18513 =  ( n18346 ) ? ( VREG_5_3 ) : ( n18512 ) ;
assign n18514 =  ( n18345 ) ? ( VREG_5_4 ) : ( n18513 ) ;
assign n18515 =  ( n18344 ) ? ( VREG_5_5 ) : ( n18514 ) ;
assign n18516 =  ( n18343 ) ? ( VREG_5_6 ) : ( n18515 ) ;
assign n18517 =  ( n18342 ) ? ( VREG_5_7 ) : ( n18516 ) ;
assign n18518 =  ( n18341 ) ? ( VREG_5_8 ) : ( n18517 ) ;
assign n18519 =  ( n18340 ) ? ( VREG_5_9 ) : ( n18518 ) ;
assign n18520 =  ( n18339 ) ? ( VREG_5_10 ) : ( n18519 ) ;
assign n18521 =  ( n18338 ) ? ( VREG_5_11 ) : ( n18520 ) ;
assign n18522 =  ( n18337 ) ? ( VREG_5_12 ) : ( n18521 ) ;
assign n18523 =  ( n18336 ) ? ( VREG_5_13 ) : ( n18522 ) ;
assign n18524 =  ( n18335 ) ? ( VREG_5_14 ) : ( n18523 ) ;
assign n18525 =  ( n18334 ) ? ( VREG_5_15 ) : ( n18524 ) ;
assign n18526 =  ( n18333 ) ? ( VREG_6_0 ) : ( n18525 ) ;
assign n18527 =  ( n18332 ) ? ( VREG_6_1 ) : ( n18526 ) ;
assign n18528 =  ( n18331 ) ? ( VREG_6_2 ) : ( n18527 ) ;
assign n18529 =  ( n18330 ) ? ( VREG_6_3 ) : ( n18528 ) ;
assign n18530 =  ( n18329 ) ? ( VREG_6_4 ) : ( n18529 ) ;
assign n18531 =  ( n18328 ) ? ( VREG_6_5 ) : ( n18530 ) ;
assign n18532 =  ( n18327 ) ? ( VREG_6_6 ) : ( n18531 ) ;
assign n18533 =  ( n18326 ) ? ( VREG_6_7 ) : ( n18532 ) ;
assign n18534 =  ( n18325 ) ? ( VREG_6_8 ) : ( n18533 ) ;
assign n18535 =  ( n18324 ) ? ( VREG_6_9 ) : ( n18534 ) ;
assign n18536 =  ( n18323 ) ? ( VREG_6_10 ) : ( n18535 ) ;
assign n18537 =  ( n18322 ) ? ( VREG_6_11 ) : ( n18536 ) ;
assign n18538 =  ( n18321 ) ? ( VREG_6_12 ) : ( n18537 ) ;
assign n18539 =  ( n18320 ) ? ( VREG_6_13 ) : ( n18538 ) ;
assign n18540 =  ( n18319 ) ? ( VREG_6_14 ) : ( n18539 ) ;
assign n18541 =  ( n18318 ) ? ( VREG_6_15 ) : ( n18540 ) ;
assign n18542 =  ( n18317 ) ? ( VREG_7_0 ) : ( n18541 ) ;
assign n18543 =  ( n18316 ) ? ( VREG_7_1 ) : ( n18542 ) ;
assign n18544 =  ( n18315 ) ? ( VREG_7_2 ) : ( n18543 ) ;
assign n18545 =  ( n18314 ) ? ( VREG_7_3 ) : ( n18544 ) ;
assign n18546 =  ( n18313 ) ? ( VREG_7_4 ) : ( n18545 ) ;
assign n18547 =  ( n18312 ) ? ( VREG_7_5 ) : ( n18546 ) ;
assign n18548 =  ( n18311 ) ? ( VREG_7_6 ) : ( n18547 ) ;
assign n18549 =  ( n18310 ) ? ( VREG_7_7 ) : ( n18548 ) ;
assign n18550 =  ( n18309 ) ? ( VREG_7_8 ) : ( n18549 ) ;
assign n18551 =  ( n18308 ) ? ( VREG_7_9 ) : ( n18550 ) ;
assign n18552 =  ( n18307 ) ? ( VREG_7_10 ) : ( n18551 ) ;
assign n18553 =  ( n18306 ) ? ( VREG_7_11 ) : ( n18552 ) ;
assign n18554 =  ( n18305 ) ? ( VREG_7_12 ) : ( n18553 ) ;
assign n18555 =  ( n18304 ) ? ( VREG_7_13 ) : ( n18554 ) ;
assign n18556 =  ( n18303 ) ? ( VREG_7_14 ) : ( n18555 ) ;
assign n18557 =  ( n18302 ) ? ( VREG_7_15 ) : ( n18556 ) ;
assign n18558 =  ( n18301 ) ? ( VREG_8_0 ) : ( n18557 ) ;
assign n18559 =  ( n18300 ) ? ( VREG_8_1 ) : ( n18558 ) ;
assign n18560 =  ( n18299 ) ? ( VREG_8_2 ) : ( n18559 ) ;
assign n18561 =  ( n18298 ) ? ( VREG_8_3 ) : ( n18560 ) ;
assign n18562 =  ( n18297 ) ? ( VREG_8_4 ) : ( n18561 ) ;
assign n18563 =  ( n18296 ) ? ( VREG_8_5 ) : ( n18562 ) ;
assign n18564 =  ( n18295 ) ? ( VREG_8_6 ) : ( n18563 ) ;
assign n18565 =  ( n18294 ) ? ( VREG_8_7 ) : ( n18564 ) ;
assign n18566 =  ( n18293 ) ? ( VREG_8_8 ) : ( n18565 ) ;
assign n18567 =  ( n18292 ) ? ( VREG_8_9 ) : ( n18566 ) ;
assign n18568 =  ( n18291 ) ? ( VREG_8_10 ) : ( n18567 ) ;
assign n18569 =  ( n18290 ) ? ( VREG_8_11 ) : ( n18568 ) ;
assign n18570 =  ( n18289 ) ? ( VREG_8_12 ) : ( n18569 ) ;
assign n18571 =  ( n18288 ) ? ( VREG_8_13 ) : ( n18570 ) ;
assign n18572 =  ( n18287 ) ? ( VREG_8_14 ) : ( n18571 ) ;
assign n18573 =  ( n18286 ) ? ( VREG_8_15 ) : ( n18572 ) ;
assign n18574 =  ( n18285 ) ? ( VREG_9_0 ) : ( n18573 ) ;
assign n18575 =  ( n18284 ) ? ( VREG_9_1 ) : ( n18574 ) ;
assign n18576 =  ( n18283 ) ? ( VREG_9_2 ) : ( n18575 ) ;
assign n18577 =  ( n18282 ) ? ( VREG_9_3 ) : ( n18576 ) ;
assign n18578 =  ( n18281 ) ? ( VREG_9_4 ) : ( n18577 ) ;
assign n18579 =  ( n18280 ) ? ( VREG_9_5 ) : ( n18578 ) ;
assign n18580 =  ( n18279 ) ? ( VREG_9_6 ) : ( n18579 ) ;
assign n18581 =  ( n18278 ) ? ( VREG_9_7 ) : ( n18580 ) ;
assign n18582 =  ( n18277 ) ? ( VREG_9_8 ) : ( n18581 ) ;
assign n18583 =  ( n18276 ) ? ( VREG_9_9 ) : ( n18582 ) ;
assign n18584 =  ( n18275 ) ? ( VREG_9_10 ) : ( n18583 ) ;
assign n18585 =  ( n18274 ) ? ( VREG_9_11 ) : ( n18584 ) ;
assign n18586 =  ( n18273 ) ? ( VREG_9_12 ) : ( n18585 ) ;
assign n18587 =  ( n18272 ) ? ( VREG_9_13 ) : ( n18586 ) ;
assign n18588 =  ( n18271 ) ? ( VREG_9_14 ) : ( n18587 ) ;
assign n18589 =  ( n18270 ) ? ( VREG_9_15 ) : ( n18588 ) ;
assign n18590 =  ( n18269 ) ? ( VREG_10_0 ) : ( n18589 ) ;
assign n18591 =  ( n18268 ) ? ( VREG_10_1 ) : ( n18590 ) ;
assign n18592 =  ( n18267 ) ? ( VREG_10_2 ) : ( n18591 ) ;
assign n18593 =  ( n18266 ) ? ( VREG_10_3 ) : ( n18592 ) ;
assign n18594 =  ( n18265 ) ? ( VREG_10_4 ) : ( n18593 ) ;
assign n18595 =  ( n18264 ) ? ( VREG_10_5 ) : ( n18594 ) ;
assign n18596 =  ( n18263 ) ? ( VREG_10_6 ) : ( n18595 ) ;
assign n18597 =  ( n18262 ) ? ( VREG_10_7 ) : ( n18596 ) ;
assign n18598 =  ( n18261 ) ? ( VREG_10_8 ) : ( n18597 ) ;
assign n18599 =  ( n18260 ) ? ( VREG_10_9 ) : ( n18598 ) ;
assign n18600 =  ( n18259 ) ? ( VREG_10_10 ) : ( n18599 ) ;
assign n18601 =  ( n18258 ) ? ( VREG_10_11 ) : ( n18600 ) ;
assign n18602 =  ( n18257 ) ? ( VREG_10_12 ) : ( n18601 ) ;
assign n18603 =  ( n18256 ) ? ( VREG_10_13 ) : ( n18602 ) ;
assign n18604 =  ( n18255 ) ? ( VREG_10_14 ) : ( n18603 ) ;
assign n18605 =  ( n18254 ) ? ( VREG_10_15 ) : ( n18604 ) ;
assign n18606 =  ( n18253 ) ? ( VREG_11_0 ) : ( n18605 ) ;
assign n18607 =  ( n18252 ) ? ( VREG_11_1 ) : ( n18606 ) ;
assign n18608 =  ( n18251 ) ? ( VREG_11_2 ) : ( n18607 ) ;
assign n18609 =  ( n18250 ) ? ( VREG_11_3 ) : ( n18608 ) ;
assign n18610 =  ( n18249 ) ? ( VREG_11_4 ) : ( n18609 ) ;
assign n18611 =  ( n18248 ) ? ( VREG_11_5 ) : ( n18610 ) ;
assign n18612 =  ( n18247 ) ? ( VREG_11_6 ) : ( n18611 ) ;
assign n18613 =  ( n18246 ) ? ( VREG_11_7 ) : ( n18612 ) ;
assign n18614 =  ( n18245 ) ? ( VREG_11_8 ) : ( n18613 ) ;
assign n18615 =  ( n18244 ) ? ( VREG_11_9 ) : ( n18614 ) ;
assign n18616 =  ( n18243 ) ? ( VREG_11_10 ) : ( n18615 ) ;
assign n18617 =  ( n18242 ) ? ( VREG_11_11 ) : ( n18616 ) ;
assign n18618 =  ( n18241 ) ? ( VREG_11_12 ) : ( n18617 ) ;
assign n18619 =  ( n18240 ) ? ( VREG_11_13 ) : ( n18618 ) ;
assign n18620 =  ( n18239 ) ? ( VREG_11_14 ) : ( n18619 ) ;
assign n18621 =  ( n18238 ) ? ( VREG_11_15 ) : ( n18620 ) ;
assign n18622 =  ( n18237 ) ? ( VREG_12_0 ) : ( n18621 ) ;
assign n18623 =  ( n18236 ) ? ( VREG_12_1 ) : ( n18622 ) ;
assign n18624 =  ( n18235 ) ? ( VREG_12_2 ) : ( n18623 ) ;
assign n18625 =  ( n18234 ) ? ( VREG_12_3 ) : ( n18624 ) ;
assign n18626 =  ( n18233 ) ? ( VREG_12_4 ) : ( n18625 ) ;
assign n18627 =  ( n18232 ) ? ( VREG_12_5 ) : ( n18626 ) ;
assign n18628 =  ( n18231 ) ? ( VREG_12_6 ) : ( n18627 ) ;
assign n18629 =  ( n18230 ) ? ( VREG_12_7 ) : ( n18628 ) ;
assign n18630 =  ( n18229 ) ? ( VREG_12_8 ) : ( n18629 ) ;
assign n18631 =  ( n18228 ) ? ( VREG_12_9 ) : ( n18630 ) ;
assign n18632 =  ( n18227 ) ? ( VREG_12_10 ) : ( n18631 ) ;
assign n18633 =  ( n18226 ) ? ( VREG_12_11 ) : ( n18632 ) ;
assign n18634 =  ( n18225 ) ? ( VREG_12_12 ) : ( n18633 ) ;
assign n18635 =  ( n18224 ) ? ( VREG_12_13 ) : ( n18634 ) ;
assign n18636 =  ( n18223 ) ? ( VREG_12_14 ) : ( n18635 ) ;
assign n18637 =  ( n18222 ) ? ( VREG_12_15 ) : ( n18636 ) ;
assign n18638 =  ( n18221 ) ? ( VREG_13_0 ) : ( n18637 ) ;
assign n18639 =  ( n18220 ) ? ( VREG_13_1 ) : ( n18638 ) ;
assign n18640 =  ( n18219 ) ? ( VREG_13_2 ) : ( n18639 ) ;
assign n18641 =  ( n18218 ) ? ( VREG_13_3 ) : ( n18640 ) ;
assign n18642 =  ( n18217 ) ? ( VREG_13_4 ) : ( n18641 ) ;
assign n18643 =  ( n18216 ) ? ( VREG_13_5 ) : ( n18642 ) ;
assign n18644 =  ( n18215 ) ? ( VREG_13_6 ) : ( n18643 ) ;
assign n18645 =  ( n18214 ) ? ( VREG_13_7 ) : ( n18644 ) ;
assign n18646 =  ( n18213 ) ? ( VREG_13_8 ) : ( n18645 ) ;
assign n18647 =  ( n18212 ) ? ( VREG_13_9 ) : ( n18646 ) ;
assign n18648 =  ( n18211 ) ? ( VREG_13_10 ) : ( n18647 ) ;
assign n18649 =  ( n18210 ) ? ( VREG_13_11 ) : ( n18648 ) ;
assign n18650 =  ( n18209 ) ? ( VREG_13_12 ) : ( n18649 ) ;
assign n18651 =  ( n18208 ) ? ( VREG_13_13 ) : ( n18650 ) ;
assign n18652 =  ( n18207 ) ? ( VREG_13_14 ) : ( n18651 ) ;
assign n18653 =  ( n18206 ) ? ( VREG_13_15 ) : ( n18652 ) ;
assign n18654 =  ( n18205 ) ? ( VREG_14_0 ) : ( n18653 ) ;
assign n18655 =  ( n18204 ) ? ( VREG_14_1 ) : ( n18654 ) ;
assign n18656 =  ( n18203 ) ? ( VREG_14_2 ) : ( n18655 ) ;
assign n18657 =  ( n18202 ) ? ( VREG_14_3 ) : ( n18656 ) ;
assign n18658 =  ( n18201 ) ? ( VREG_14_4 ) : ( n18657 ) ;
assign n18659 =  ( n18200 ) ? ( VREG_14_5 ) : ( n18658 ) ;
assign n18660 =  ( n18199 ) ? ( VREG_14_6 ) : ( n18659 ) ;
assign n18661 =  ( n18198 ) ? ( VREG_14_7 ) : ( n18660 ) ;
assign n18662 =  ( n18197 ) ? ( VREG_14_8 ) : ( n18661 ) ;
assign n18663 =  ( n18196 ) ? ( VREG_14_9 ) : ( n18662 ) ;
assign n18664 =  ( n18195 ) ? ( VREG_14_10 ) : ( n18663 ) ;
assign n18665 =  ( n18194 ) ? ( VREG_14_11 ) : ( n18664 ) ;
assign n18666 =  ( n18193 ) ? ( VREG_14_12 ) : ( n18665 ) ;
assign n18667 =  ( n18192 ) ? ( VREG_14_13 ) : ( n18666 ) ;
assign n18668 =  ( n18191 ) ? ( VREG_14_14 ) : ( n18667 ) ;
assign n18669 =  ( n18190 ) ? ( VREG_14_15 ) : ( n18668 ) ;
assign n18670 =  ( n18189 ) ? ( VREG_15_0 ) : ( n18669 ) ;
assign n18671 =  ( n18188 ) ? ( VREG_15_1 ) : ( n18670 ) ;
assign n18672 =  ( n18187 ) ? ( VREG_15_2 ) : ( n18671 ) ;
assign n18673 =  ( n18186 ) ? ( VREG_15_3 ) : ( n18672 ) ;
assign n18674 =  ( n18185 ) ? ( VREG_15_4 ) : ( n18673 ) ;
assign n18675 =  ( n18184 ) ? ( VREG_15_5 ) : ( n18674 ) ;
assign n18676 =  ( n18183 ) ? ( VREG_15_6 ) : ( n18675 ) ;
assign n18677 =  ( n18182 ) ? ( VREG_15_7 ) : ( n18676 ) ;
assign n18678 =  ( n18181 ) ? ( VREG_15_8 ) : ( n18677 ) ;
assign n18679 =  ( n18180 ) ? ( VREG_15_9 ) : ( n18678 ) ;
assign n18680 =  ( n18179 ) ? ( VREG_15_10 ) : ( n18679 ) ;
assign n18681 =  ( n18178 ) ? ( VREG_15_11 ) : ( n18680 ) ;
assign n18682 =  ( n18177 ) ? ( VREG_15_12 ) : ( n18681 ) ;
assign n18683 =  ( n18176 ) ? ( VREG_15_13 ) : ( n18682 ) ;
assign n18684 =  ( n18175 ) ? ( VREG_15_14 ) : ( n18683 ) ;
assign n18685 =  ( n18174 ) ? ( VREG_15_15 ) : ( n18684 ) ;
assign n18686 =  ( n18173 ) ? ( VREG_16_0 ) : ( n18685 ) ;
assign n18687 =  ( n18172 ) ? ( VREG_16_1 ) : ( n18686 ) ;
assign n18688 =  ( n18171 ) ? ( VREG_16_2 ) : ( n18687 ) ;
assign n18689 =  ( n18170 ) ? ( VREG_16_3 ) : ( n18688 ) ;
assign n18690 =  ( n18169 ) ? ( VREG_16_4 ) : ( n18689 ) ;
assign n18691 =  ( n18168 ) ? ( VREG_16_5 ) : ( n18690 ) ;
assign n18692 =  ( n18167 ) ? ( VREG_16_6 ) : ( n18691 ) ;
assign n18693 =  ( n18166 ) ? ( VREG_16_7 ) : ( n18692 ) ;
assign n18694 =  ( n18165 ) ? ( VREG_16_8 ) : ( n18693 ) ;
assign n18695 =  ( n18164 ) ? ( VREG_16_9 ) : ( n18694 ) ;
assign n18696 =  ( n18163 ) ? ( VREG_16_10 ) : ( n18695 ) ;
assign n18697 =  ( n18162 ) ? ( VREG_16_11 ) : ( n18696 ) ;
assign n18698 =  ( n18161 ) ? ( VREG_16_12 ) : ( n18697 ) ;
assign n18699 =  ( n18160 ) ? ( VREG_16_13 ) : ( n18698 ) ;
assign n18700 =  ( n18159 ) ? ( VREG_16_14 ) : ( n18699 ) ;
assign n18701 =  ( n18158 ) ? ( VREG_16_15 ) : ( n18700 ) ;
assign n18702 =  ( n18157 ) ? ( VREG_17_0 ) : ( n18701 ) ;
assign n18703 =  ( n18156 ) ? ( VREG_17_1 ) : ( n18702 ) ;
assign n18704 =  ( n18155 ) ? ( VREG_17_2 ) : ( n18703 ) ;
assign n18705 =  ( n18154 ) ? ( VREG_17_3 ) : ( n18704 ) ;
assign n18706 =  ( n18153 ) ? ( VREG_17_4 ) : ( n18705 ) ;
assign n18707 =  ( n18152 ) ? ( VREG_17_5 ) : ( n18706 ) ;
assign n18708 =  ( n18151 ) ? ( VREG_17_6 ) : ( n18707 ) ;
assign n18709 =  ( n18150 ) ? ( VREG_17_7 ) : ( n18708 ) ;
assign n18710 =  ( n18149 ) ? ( VREG_17_8 ) : ( n18709 ) ;
assign n18711 =  ( n18148 ) ? ( VREG_17_9 ) : ( n18710 ) ;
assign n18712 =  ( n18147 ) ? ( VREG_17_10 ) : ( n18711 ) ;
assign n18713 =  ( n18146 ) ? ( VREG_17_11 ) : ( n18712 ) ;
assign n18714 =  ( n18145 ) ? ( VREG_17_12 ) : ( n18713 ) ;
assign n18715 =  ( n18144 ) ? ( VREG_17_13 ) : ( n18714 ) ;
assign n18716 =  ( n18143 ) ? ( VREG_17_14 ) : ( n18715 ) ;
assign n18717 =  ( n18142 ) ? ( VREG_17_15 ) : ( n18716 ) ;
assign n18718 =  ( n18141 ) ? ( VREG_18_0 ) : ( n18717 ) ;
assign n18719 =  ( n18140 ) ? ( VREG_18_1 ) : ( n18718 ) ;
assign n18720 =  ( n18139 ) ? ( VREG_18_2 ) : ( n18719 ) ;
assign n18721 =  ( n18138 ) ? ( VREG_18_3 ) : ( n18720 ) ;
assign n18722 =  ( n18137 ) ? ( VREG_18_4 ) : ( n18721 ) ;
assign n18723 =  ( n18136 ) ? ( VREG_18_5 ) : ( n18722 ) ;
assign n18724 =  ( n18135 ) ? ( VREG_18_6 ) : ( n18723 ) ;
assign n18725 =  ( n18134 ) ? ( VREG_18_7 ) : ( n18724 ) ;
assign n18726 =  ( n18133 ) ? ( VREG_18_8 ) : ( n18725 ) ;
assign n18727 =  ( n18132 ) ? ( VREG_18_9 ) : ( n18726 ) ;
assign n18728 =  ( n18131 ) ? ( VREG_18_10 ) : ( n18727 ) ;
assign n18729 =  ( n18130 ) ? ( VREG_18_11 ) : ( n18728 ) ;
assign n18730 =  ( n18129 ) ? ( VREG_18_12 ) : ( n18729 ) ;
assign n18731 =  ( n18128 ) ? ( VREG_18_13 ) : ( n18730 ) ;
assign n18732 =  ( n18127 ) ? ( VREG_18_14 ) : ( n18731 ) ;
assign n18733 =  ( n18126 ) ? ( VREG_18_15 ) : ( n18732 ) ;
assign n18734 =  ( n18125 ) ? ( VREG_19_0 ) : ( n18733 ) ;
assign n18735 =  ( n18124 ) ? ( VREG_19_1 ) : ( n18734 ) ;
assign n18736 =  ( n18123 ) ? ( VREG_19_2 ) : ( n18735 ) ;
assign n18737 =  ( n18122 ) ? ( VREG_19_3 ) : ( n18736 ) ;
assign n18738 =  ( n18121 ) ? ( VREG_19_4 ) : ( n18737 ) ;
assign n18739 =  ( n18120 ) ? ( VREG_19_5 ) : ( n18738 ) ;
assign n18740 =  ( n18119 ) ? ( VREG_19_6 ) : ( n18739 ) ;
assign n18741 =  ( n18118 ) ? ( VREG_19_7 ) : ( n18740 ) ;
assign n18742 =  ( n18117 ) ? ( VREG_19_8 ) : ( n18741 ) ;
assign n18743 =  ( n18116 ) ? ( VREG_19_9 ) : ( n18742 ) ;
assign n18744 =  ( n18115 ) ? ( VREG_19_10 ) : ( n18743 ) ;
assign n18745 =  ( n18114 ) ? ( VREG_19_11 ) : ( n18744 ) ;
assign n18746 =  ( n18113 ) ? ( VREG_19_12 ) : ( n18745 ) ;
assign n18747 =  ( n18112 ) ? ( VREG_19_13 ) : ( n18746 ) ;
assign n18748 =  ( n18111 ) ? ( VREG_19_14 ) : ( n18747 ) ;
assign n18749 =  ( n18110 ) ? ( VREG_19_15 ) : ( n18748 ) ;
assign n18750 =  ( n18109 ) ? ( VREG_20_0 ) : ( n18749 ) ;
assign n18751 =  ( n18108 ) ? ( VREG_20_1 ) : ( n18750 ) ;
assign n18752 =  ( n18107 ) ? ( VREG_20_2 ) : ( n18751 ) ;
assign n18753 =  ( n18106 ) ? ( VREG_20_3 ) : ( n18752 ) ;
assign n18754 =  ( n18105 ) ? ( VREG_20_4 ) : ( n18753 ) ;
assign n18755 =  ( n18104 ) ? ( VREG_20_5 ) : ( n18754 ) ;
assign n18756 =  ( n18103 ) ? ( VREG_20_6 ) : ( n18755 ) ;
assign n18757 =  ( n18102 ) ? ( VREG_20_7 ) : ( n18756 ) ;
assign n18758 =  ( n18101 ) ? ( VREG_20_8 ) : ( n18757 ) ;
assign n18759 =  ( n18100 ) ? ( VREG_20_9 ) : ( n18758 ) ;
assign n18760 =  ( n18099 ) ? ( VREG_20_10 ) : ( n18759 ) ;
assign n18761 =  ( n18098 ) ? ( VREG_20_11 ) : ( n18760 ) ;
assign n18762 =  ( n18097 ) ? ( VREG_20_12 ) : ( n18761 ) ;
assign n18763 =  ( n18096 ) ? ( VREG_20_13 ) : ( n18762 ) ;
assign n18764 =  ( n18095 ) ? ( VREG_20_14 ) : ( n18763 ) ;
assign n18765 =  ( n18094 ) ? ( VREG_20_15 ) : ( n18764 ) ;
assign n18766 =  ( n18093 ) ? ( VREG_21_0 ) : ( n18765 ) ;
assign n18767 =  ( n18092 ) ? ( VREG_21_1 ) : ( n18766 ) ;
assign n18768 =  ( n18091 ) ? ( VREG_21_2 ) : ( n18767 ) ;
assign n18769 =  ( n18090 ) ? ( VREG_21_3 ) : ( n18768 ) ;
assign n18770 =  ( n18089 ) ? ( VREG_21_4 ) : ( n18769 ) ;
assign n18771 =  ( n18088 ) ? ( VREG_21_5 ) : ( n18770 ) ;
assign n18772 =  ( n18087 ) ? ( VREG_21_6 ) : ( n18771 ) ;
assign n18773 =  ( n18086 ) ? ( VREG_21_7 ) : ( n18772 ) ;
assign n18774 =  ( n18085 ) ? ( VREG_21_8 ) : ( n18773 ) ;
assign n18775 =  ( n18084 ) ? ( VREG_21_9 ) : ( n18774 ) ;
assign n18776 =  ( n18083 ) ? ( VREG_21_10 ) : ( n18775 ) ;
assign n18777 =  ( n18082 ) ? ( VREG_21_11 ) : ( n18776 ) ;
assign n18778 =  ( n18081 ) ? ( VREG_21_12 ) : ( n18777 ) ;
assign n18779 =  ( n18080 ) ? ( VREG_21_13 ) : ( n18778 ) ;
assign n18780 =  ( n18079 ) ? ( VREG_21_14 ) : ( n18779 ) ;
assign n18781 =  ( n18078 ) ? ( VREG_21_15 ) : ( n18780 ) ;
assign n18782 =  ( n18077 ) ? ( VREG_22_0 ) : ( n18781 ) ;
assign n18783 =  ( n18076 ) ? ( VREG_22_1 ) : ( n18782 ) ;
assign n18784 =  ( n18075 ) ? ( VREG_22_2 ) : ( n18783 ) ;
assign n18785 =  ( n18074 ) ? ( VREG_22_3 ) : ( n18784 ) ;
assign n18786 =  ( n18073 ) ? ( VREG_22_4 ) : ( n18785 ) ;
assign n18787 =  ( n18072 ) ? ( VREG_22_5 ) : ( n18786 ) ;
assign n18788 =  ( n18071 ) ? ( VREG_22_6 ) : ( n18787 ) ;
assign n18789 =  ( n18070 ) ? ( VREG_22_7 ) : ( n18788 ) ;
assign n18790 =  ( n18069 ) ? ( VREG_22_8 ) : ( n18789 ) ;
assign n18791 =  ( n18068 ) ? ( VREG_22_9 ) : ( n18790 ) ;
assign n18792 =  ( n18067 ) ? ( VREG_22_10 ) : ( n18791 ) ;
assign n18793 =  ( n18066 ) ? ( VREG_22_11 ) : ( n18792 ) ;
assign n18794 =  ( n18065 ) ? ( VREG_22_12 ) : ( n18793 ) ;
assign n18795 =  ( n18064 ) ? ( VREG_22_13 ) : ( n18794 ) ;
assign n18796 =  ( n18063 ) ? ( VREG_22_14 ) : ( n18795 ) ;
assign n18797 =  ( n18062 ) ? ( VREG_22_15 ) : ( n18796 ) ;
assign n18798 =  ( n18061 ) ? ( VREG_23_0 ) : ( n18797 ) ;
assign n18799 =  ( n18060 ) ? ( VREG_23_1 ) : ( n18798 ) ;
assign n18800 =  ( n18059 ) ? ( VREG_23_2 ) : ( n18799 ) ;
assign n18801 =  ( n18058 ) ? ( VREG_23_3 ) : ( n18800 ) ;
assign n18802 =  ( n18057 ) ? ( VREG_23_4 ) : ( n18801 ) ;
assign n18803 =  ( n18056 ) ? ( VREG_23_5 ) : ( n18802 ) ;
assign n18804 =  ( n18055 ) ? ( VREG_23_6 ) : ( n18803 ) ;
assign n18805 =  ( n18054 ) ? ( VREG_23_7 ) : ( n18804 ) ;
assign n18806 =  ( n18053 ) ? ( VREG_23_8 ) : ( n18805 ) ;
assign n18807 =  ( n18052 ) ? ( VREG_23_9 ) : ( n18806 ) ;
assign n18808 =  ( n18051 ) ? ( VREG_23_10 ) : ( n18807 ) ;
assign n18809 =  ( n18050 ) ? ( VREG_23_11 ) : ( n18808 ) ;
assign n18810 =  ( n18049 ) ? ( VREG_23_12 ) : ( n18809 ) ;
assign n18811 =  ( n18048 ) ? ( VREG_23_13 ) : ( n18810 ) ;
assign n18812 =  ( n18047 ) ? ( VREG_23_14 ) : ( n18811 ) ;
assign n18813 =  ( n18046 ) ? ( VREG_23_15 ) : ( n18812 ) ;
assign n18814 =  ( n18045 ) ? ( VREG_24_0 ) : ( n18813 ) ;
assign n18815 =  ( n18044 ) ? ( VREG_24_1 ) : ( n18814 ) ;
assign n18816 =  ( n18043 ) ? ( VREG_24_2 ) : ( n18815 ) ;
assign n18817 =  ( n18042 ) ? ( VREG_24_3 ) : ( n18816 ) ;
assign n18818 =  ( n18041 ) ? ( VREG_24_4 ) : ( n18817 ) ;
assign n18819 =  ( n18040 ) ? ( VREG_24_5 ) : ( n18818 ) ;
assign n18820 =  ( n18039 ) ? ( VREG_24_6 ) : ( n18819 ) ;
assign n18821 =  ( n18038 ) ? ( VREG_24_7 ) : ( n18820 ) ;
assign n18822 =  ( n18037 ) ? ( VREG_24_8 ) : ( n18821 ) ;
assign n18823 =  ( n18036 ) ? ( VREG_24_9 ) : ( n18822 ) ;
assign n18824 =  ( n18035 ) ? ( VREG_24_10 ) : ( n18823 ) ;
assign n18825 =  ( n18034 ) ? ( VREG_24_11 ) : ( n18824 ) ;
assign n18826 =  ( n18033 ) ? ( VREG_24_12 ) : ( n18825 ) ;
assign n18827 =  ( n18032 ) ? ( VREG_24_13 ) : ( n18826 ) ;
assign n18828 =  ( n18031 ) ? ( VREG_24_14 ) : ( n18827 ) ;
assign n18829 =  ( n18030 ) ? ( VREG_24_15 ) : ( n18828 ) ;
assign n18830 =  ( n18029 ) ? ( VREG_25_0 ) : ( n18829 ) ;
assign n18831 =  ( n18028 ) ? ( VREG_25_1 ) : ( n18830 ) ;
assign n18832 =  ( n18027 ) ? ( VREG_25_2 ) : ( n18831 ) ;
assign n18833 =  ( n18026 ) ? ( VREG_25_3 ) : ( n18832 ) ;
assign n18834 =  ( n18025 ) ? ( VREG_25_4 ) : ( n18833 ) ;
assign n18835 =  ( n18024 ) ? ( VREG_25_5 ) : ( n18834 ) ;
assign n18836 =  ( n18023 ) ? ( VREG_25_6 ) : ( n18835 ) ;
assign n18837 =  ( n18022 ) ? ( VREG_25_7 ) : ( n18836 ) ;
assign n18838 =  ( n18021 ) ? ( VREG_25_8 ) : ( n18837 ) ;
assign n18839 =  ( n18020 ) ? ( VREG_25_9 ) : ( n18838 ) ;
assign n18840 =  ( n18019 ) ? ( VREG_25_10 ) : ( n18839 ) ;
assign n18841 =  ( n18018 ) ? ( VREG_25_11 ) : ( n18840 ) ;
assign n18842 =  ( n18017 ) ? ( VREG_25_12 ) : ( n18841 ) ;
assign n18843 =  ( n18016 ) ? ( VREG_25_13 ) : ( n18842 ) ;
assign n18844 =  ( n18015 ) ? ( VREG_25_14 ) : ( n18843 ) ;
assign n18845 =  ( n18014 ) ? ( VREG_25_15 ) : ( n18844 ) ;
assign n18846 =  ( n18013 ) ? ( VREG_26_0 ) : ( n18845 ) ;
assign n18847 =  ( n18012 ) ? ( VREG_26_1 ) : ( n18846 ) ;
assign n18848 =  ( n18011 ) ? ( VREG_26_2 ) : ( n18847 ) ;
assign n18849 =  ( n18010 ) ? ( VREG_26_3 ) : ( n18848 ) ;
assign n18850 =  ( n18009 ) ? ( VREG_26_4 ) : ( n18849 ) ;
assign n18851 =  ( n18008 ) ? ( VREG_26_5 ) : ( n18850 ) ;
assign n18852 =  ( n18007 ) ? ( VREG_26_6 ) : ( n18851 ) ;
assign n18853 =  ( n18006 ) ? ( VREG_26_7 ) : ( n18852 ) ;
assign n18854 =  ( n18005 ) ? ( VREG_26_8 ) : ( n18853 ) ;
assign n18855 =  ( n18004 ) ? ( VREG_26_9 ) : ( n18854 ) ;
assign n18856 =  ( n18003 ) ? ( VREG_26_10 ) : ( n18855 ) ;
assign n18857 =  ( n18002 ) ? ( VREG_26_11 ) : ( n18856 ) ;
assign n18858 =  ( n18001 ) ? ( VREG_26_12 ) : ( n18857 ) ;
assign n18859 =  ( n18000 ) ? ( VREG_26_13 ) : ( n18858 ) ;
assign n18860 =  ( n17999 ) ? ( VREG_26_14 ) : ( n18859 ) ;
assign n18861 =  ( n17998 ) ? ( VREG_26_15 ) : ( n18860 ) ;
assign n18862 =  ( n17997 ) ? ( VREG_27_0 ) : ( n18861 ) ;
assign n18863 =  ( n17996 ) ? ( VREG_27_1 ) : ( n18862 ) ;
assign n18864 =  ( n17995 ) ? ( VREG_27_2 ) : ( n18863 ) ;
assign n18865 =  ( n17994 ) ? ( VREG_27_3 ) : ( n18864 ) ;
assign n18866 =  ( n17993 ) ? ( VREG_27_4 ) : ( n18865 ) ;
assign n18867 =  ( n17992 ) ? ( VREG_27_5 ) : ( n18866 ) ;
assign n18868 =  ( n17991 ) ? ( VREG_27_6 ) : ( n18867 ) ;
assign n18869 =  ( n17990 ) ? ( VREG_27_7 ) : ( n18868 ) ;
assign n18870 =  ( n17989 ) ? ( VREG_27_8 ) : ( n18869 ) ;
assign n18871 =  ( n17988 ) ? ( VREG_27_9 ) : ( n18870 ) ;
assign n18872 =  ( n17987 ) ? ( VREG_27_10 ) : ( n18871 ) ;
assign n18873 =  ( n17986 ) ? ( VREG_27_11 ) : ( n18872 ) ;
assign n18874 =  ( n17985 ) ? ( VREG_27_12 ) : ( n18873 ) ;
assign n18875 =  ( n17984 ) ? ( VREG_27_13 ) : ( n18874 ) ;
assign n18876 =  ( n17983 ) ? ( VREG_27_14 ) : ( n18875 ) ;
assign n18877 =  ( n17982 ) ? ( VREG_27_15 ) : ( n18876 ) ;
assign n18878 =  ( n17981 ) ? ( VREG_28_0 ) : ( n18877 ) ;
assign n18879 =  ( n17980 ) ? ( VREG_28_1 ) : ( n18878 ) ;
assign n18880 =  ( n17979 ) ? ( VREG_28_2 ) : ( n18879 ) ;
assign n18881 =  ( n17978 ) ? ( VREG_28_3 ) : ( n18880 ) ;
assign n18882 =  ( n17977 ) ? ( VREG_28_4 ) : ( n18881 ) ;
assign n18883 =  ( n17976 ) ? ( VREG_28_5 ) : ( n18882 ) ;
assign n18884 =  ( n17975 ) ? ( VREG_28_6 ) : ( n18883 ) ;
assign n18885 =  ( n17974 ) ? ( VREG_28_7 ) : ( n18884 ) ;
assign n18886 =  ( n17973 ) ? ( VREG_28_8 ) : ( n18885 ) ;
assign n18887 =  ( n17972 ) ? ( VREG_28_9 ) : ( n18886 ) ;
assign n18888 =  ( n17971 ) ? ( VREG_28_10 ) : ( n18887 ) ;
assign n18889 =  ( n17970 ) ? ( VREG_28_11 ) : ( n18888 ) ;
assign n18890 =  ( n17969 ) ? ( VREG_28_12 ) : ( n18889 ) ;
assign n18891 =  ( n17968 ) ? ( VREG_28_13 ) : ( n18890 ) ;
assign n18892 =  ( n17967 ) ? ( VREG_28_14 ) : ( n18891 ) ;
assign n18893 =  ( n17966 ) ? ( VREG_28_15 ) : ( n18892 ) ;
assign n18894 =  ( n17965 ) ? ( VREG_29_0 ) : ( n18893 ) ;
assign n18895 =  ( n17964 ) ? ( VREG_29_1 ) : ( n18894 ) ;
assign n18896 =  ( n17963 ) ? ( VREG_29_2 ) : ( n18895 ) ;
assign n18897 =  ( n17962 ) ? ( VREG_29_3 ) : ( n18896 ) ;
assign n18898 =  ( n17961 ) ? ( VREG_29_4 ) : ( n18897 ) ;
assign n18899 =  ( n17960 ) ? ( VREG_29_5 ) : ( n18898 ) ;
assign n18900 =  ( n17959 ) ? ( VREG_29_6 ) : ( n18899 ) ;
assign n18901 =  ( n17958 ) ? ( VREG_29_7 ) : ( n18900 ) ;
assign n18902 =  ( n17957 ) ? ( VREG_29_8 ) : ( n18901 ) ;
assign n18903 =  ( n17956 ) ? ( VREG_29_9 ) : ( n18902 ) ;
assign n18904 =  ( n17955 ) ? ( VREG_29_10 ) : ( n18903 ) ;
assign n18905 =  ( n17954 ) ? ( VREG_29_11 ) : ( n18904 ) ;
assign n18906 =  ( n17953 ) ? ( VREG_29_12 ) : ( n18905 ) ;
assign n18907 =  ( n17952 ) ? ( VREG_29_13 ) : ( n18906 ) ;
assign n18908 =  ( n17951 ) ? ( VREG_29_14 ) : ( n18907 ) ;
assign n18909 =  ( n17950 ) ? ( VREG_29_15 ) : ( n18908 ) ;
assign n18910 =  ( n17949 ) ? ( VREG_30_0 ) : ( n18909 ) ;
assign n18911 =  ( n17948 ) ? ( VREG_30_1 ) : ( n18910 ) ;
assign n18912 =  ( n17947 ) ? ( VREG_30_2 ) : ( n18911 ) ;
assign n18913 =  ( n17946 ) ? ( VREG_30_3 ) : ( n18912 ) ;
assign n18914 =  ( n17945 ) ? ( VREG_30_4 ) : ( n18913 ) ;
assign n18915 =  ( n17944 ) ? ( VREG_30_5 ) : ( n18914 ) ;
assign n18916 =  ( n17943 ) ? ( VREG_30_6 ) : ( n18915 ) ;
assign n18917 =  ( n17942 ) ? ( VREG_30_7 ) : ( n18916 ) ;
assign n18918 =  ( n17941 ) ? ( VREG_30_8 ) : ( n18917 ) ;
assign n18919 =  ( n17940 ) ? ( VREG_30_9 ) : ( n18918 ) ;
assign n18920 =  ( n17939 ) ? ( VREG_30_10 ) : ( n18919 ) ;
assign n18921 =  ( n17938 ) ? ( VREG_30_11 ) : ( n18920 ) ;
assign n18922 =  ( n17937 ) ? ( VREG_30_12 ) : ( n18921 ) ;
assign n18923 =  ( n17936 ) ? ( VREG_30_13 ) : ( n18922 ) ;
assign n18924 =  ( n17935 ) ? ( VREG_30_14 ) : ( n18923 ) ;
assign n18925 =  ( n17934 ) ? ( VREG_30_15 ) : ( n18924 ) ;
assign n18926 =  ( n17933 ) ? ( VREG_31_0 ) : ( n18925 ) ;
assign n18927 =  ( n17931 ) ? ( VREG_31_1 ) : ( n18926 ) ;
assign n18928 =  ( n17929 ) ? ( VREG_31_2 ) : ( n18927 ) ;
assign n18929 =  ( n17927 ) ? ( VREG_31_3 ) : ( n18928 ) ;
assign n18930 =  ( n17925 ) ? ( VREG_31_4 ) : ( n18929 ) ;
assign n18931 =  ( n17923 ) ? ( VREG_31_5 ) : ( n18930 ) ;
assign n18932 =  ( n17921 ) ? ( VREG_31_6 ) : ( n18931 ) ;
assign n18933 =  ( n17919 ) ? ( VREG_31_7 ) : ( n18932 ) ;
assign n18934 =  ( n17917 ) ? ( VREG_31_8 ) : ( n18933 ) ;
assign n18935 =  ( n17915 ) ? ( VREG_31_9 ) : ( n18934 ) ;
assign n18936 =  ( n17913 ) ? ( VREG_31_10 ) : ( n18935 ) ;
assign n18937 =  ( n17911 ) ? ( VREG_31_11 ) : ( n18936 ) ;
assign n18938 =  ( n17909 ) ? ( VREG_31_12 ) : ( n18937 ) ;
assign n18939 =  ( n17907 ) ? ( VREG_31_13 ) : ( n18938 ) ;
assign n18940 =  ( n17905 ) ? ( VREG_31_14 ) : ( n18939 ) ;
assign n18941 =  ( n17903 ) ? ( VREG_31_15 ) : ( n18940 ) ;
assign n18942 =  ( n18941 ) + ( n140 )  ;
assign n18943 =  ( n18941 ) - ( n140 )  ;
assign n18944 =  ( n18941 ) & ( n140 )  ;
assign n18945 =  ( n18941 ) | ( n140 )  ;
assign n18946 =  ( ( n18941 ) * ( n140 ))  ;
assign n18947 =  ( n148 ) ? ( n18946 ) : ( VREG_0_2 ) ;
assign n18948 =  ( n146 ) ? ( n18945 ) : ( n18947 ) ;
assign n18949 =  ( n144 ) ? ( n18944 ) : ( n18948 ) ;
assign n18950 =  ( n142 ) ? ( n18943 ) : ( n18949 ) ;
assign n18951 =  ( n10 ) ? ( n18942 ) : ( n18950 ) ;
assign n18952 =  ( n77 ) & ( n17902 )  ;
assign n18953 =  ( n77 ) & ( n17904 )  ;
assign n18954 =  ( n77 ) & ( n17906 )  ;
assign n18955 =  ( n77 ) & ( n17908 )  ;
assign n18956 =  ( n77 ) & ( n17910 )  ;
assign n18957 =  ( n77 ) & ( n17912 )  ;
assign n18958 =  ( n77 ) & ( n17914 )  ;
assign n18959 =  ( n77 ) & ( n17916 )  ;
assign n18960 =  ( n77 ) & ( n17918 )  ;
assign n18961 =  ( n77 ) & ( n17920 )  ;
assign n18962 =  ( n77 ) & ( n17922 )  ;
assign n18963 =  ( n77 ) & ( n17924 )  ;
assign n18964 =  ( n77 ) & ( n17926 )  ;
assign n18965 =  ( n77 ) & ( n17928 )  ;
assign n18966 =  ( n77 ) & ( n17930 )  ;
assign n18967 =  ( n77 ) & ( n17932 )  ;
assign n18968 =  ( n78 ) & ( n17902 )  ;
assign n18969 =  ( n78 ) & ( n17904 )  ;
assign n18970 =  ( n78 ) & ( n17906 )  ;
assign n18971 =  ( n78 ) & ( n17908 )  ;
assign n18972 =  ( n78 ) & ( n17910 )  ;
assign n18973 =  ( n78 ) & ( n17912 )  ;
assign n18974 =  ( n78 ) & ( n17914 )  ;
assign n18975 =  ( n78 ) & ( n17916 )  ;
assign n18976 =  ( n78 ) & ( n17918 )  ;
assign n18977 =  ( n78 ) & ( n17920 )  ;
assign n18978 =  ( n78 ) & ( n17922 )  ;
assign n18979 =  ( n78 ) & ( n17924 )  ;
assign n18980 =  ( n78 ) & ( n17926 )  ;
assign n18981 =  ( n78 ) & ( n17928 )  ;
assign n18982 =  ( n78 ) & ( n17930 )  ;
assign n18983 =  ( n78 ) & ( n17932 )  ;
assign n18984 =  ( n79 ) & ( n17902 )  ;
assign n18985 =  ( n79 ) & ( n17904 )  ;
assign n18986 =  ( n79 ) & ( n17906 )  ;
assign n18987 =  ( n79 ) & ( n17908 )  ;
assign n18988 =  ( n79 ) & ( n17910 )  ;
assign n18989 =  ( n79 ) & ( n17912 )  ;
assign n18990 =  ( n79 ) & ( n17914 )  ;
assign n18991 =  ( n79 ) & ( n17916 )  ;
assign n18992 =  ( n79 ) & ( n17918 )  ;
assign n18993 =  ( n79 ) & ( n17920 )  ;
assign n18994 =  ( n79 ) & ( n17922 )  ;
assign n18995 =  ( n79 ) & ( n17924 )  ;
assign n18996 =  ( n79 ) & ( n17926 )  ;
assign n18997 =  ( n79 ) & ( n17928 )  ;
assign n18998 =  ( n79 ) & ( n17930 )  ;
assign n18999 =  ( n79 ) & ( n17932 )  ;
assign n19000 =  ( n80 ) & ( n17902 )  ;
assign n19001 =  ( n80 ) & ( n17904 )  ;
assign n19002 =  ( n80 ) & ( n17906 )  ;
assign n19003 =  ( n80 ) & ( n17908 )  ;
assign n19004 =  ( n80 ) & ( n17910 )  ;
assign n19005 =  ( n80 ) & ( n17912 )  ;
assign n19006 =  ( n80 ) & ( n17914 )  ;
assign n19007 =  ( n80 ) & ( n17916 )  ;
assign n19008 =  ( n80 ) & ( n17918 )  ;
assign n19009 =  ( n80 ) & ( n17920 )  ;
assign n19010 =  ( n80 ) & ( n17922 )  ;
assign n19011 =  ( n80 ) & ( n17924 )  ;
assign n19012 =  ( n80 ) & ( n17926 )  ;
assign n19013 =  ( n80 ) & ( n17928 )  ;
assign n19014 =  ( n80 ) & ( n17930 )  ;
assign n19015 =  ( n80 ) & ( n17932 )  ;
assign n19016 =  ( n81 ) & ( n17902 )  ;
assign n19017 =  ( n81 ) & ( n17904 )  ;
assign n19018 =  ( n81 ) & ( n17906 )  ;
assign n19019 =  ( n81 ) & ( n17908 )  ;
assign n19020 =  ( n81 ) & ( n17910 )  ;
assign n19021 =  ( n81 ) & ( n17912 )  ;
assign n19022 =  ( n81 ) & ( n17914 )  ;
assign n19023 =  ( n81 ) & ( n17916 )  ;
assign n19024 =  ( n81 ) & ( n17918 )  ;
assign n19025 =  ( n81 ) & ( n17920 )  ;
assign n19026 =  ( n81 ) & ( n17922 )  ;
assign n19027 =  ( n81 ) & ( n17924 )  ;
assign n19028 =  ( n81 ) & ( n17926 )  ;
assign n19029 =  ( n81 ) & ( n17928 )  ;
assign n19030 =  ( n81 ) & ( n17930 )  ;
assign n19031 =  ( n81 ) & ( n17932 )  ;
assign n19032 =  ( n82 ) & ( n17902 )  ;
assign n19033 =  ( n82 ) & ( n17904 )  ;
assign n19034 =  ( n82 ) & ( n17906 )  ;
assign n19035 =  ( n82 ) & ( n17908 )  ;
assign n19036 =  ( n82 ) & ( n17910 )  ;
assign n19037 =  ( n82 ) & ( n17912 )  ;
assign n19038 =  ( n82 ) & ( n17914 )  ;
assign n19039 =  ( n82 ) & ( n17916 )  ;
assign n19040 =  ( n82 ) & ( n17918 )  ;
assign n19041 =  ( n82 ) & ( n17920 )  ;
assign n19042 =  ( n82 ) & ( n17922 )  ;
assign n19043 =  ( n82 ) & ( n17924 )  ;
assign n19044 =  ( n82 ) & ( n17926 )  ;
assign n19045 =  ( n82 ) & ( n17928 )  ;
assign n19046 =  ( n82 ) & ( n17930 )  ;
assign n19047 =  ( n82 ) & ( n17932 )  ;
assign n19048 =  ( n83 ) & ( n17902 )  ;
assign n19049 =  ( n83 ) & ( n17904 )  ;
assign n19050 =  ( n83 ) & ( n17906 )  ;
assign n19051 =  ( n83 ) & ( n17908 )  ;
assign n19052 =  ( n83 ) & ( n17910 )  ;
assign n19053 =  ( n83 ) & ( n17912 )  ;
assign n19054 =  ( n83 ) & ( n17914 )  ;
assign n19055 =  ( n83 ) & ( n17916 )  ;
assign n19056 =  ( n83 ) & ( n17918 )  ;
assign n19057 =  ( n83 ) & ( n17920 )  ;
assign n19058 =  ( n83 ) & ( n17922 )  ;
assign n19059 =  ( n83 ) & ( n17924 )  ;
assign n19060 =  ( n83 ) & ( n17926 )  ;
assign n19061 =  ( n83 ) & ( n17928 )  ;
assign n19062 =  ( n83 ) & ( n17930 )  ;
assign n19063 =  ( n83 ) & ( n17932 )  ;
assign n19064 =  ( n84 ) & ( n17902 )  ;
assign n19065 =  ( n84 ) & ( n17904 )  ;
assign n19066 =  ( n84 ) & ( n17906 )  ;
assign n19067 =  ( n84 ) & ( n17908 )  ;
assign n19068 =  ( n84 ) & ( n17910 )  ;
assign n19069 =  ( n84 ) & ( n17912 )  ;
assign n19070 =  ( n84 ) & ( n17914 )  ;
assign n19071 =  ( n84 ) & ( n17916 )  ;
assign n19072 =  ( n84 ) & ( n17918 )  ;
assign n19073 =  ( n84 ) & ( n17920 )  ;
assign n19074 =  ( n84 ) & ( n17922 )  ;
assign n19075 =  ( n84 ) & ( n17924 )  ;
assign n19076 =  ( n84 ) & ( n17926 )  ;
assign n19077 =  ( n84 ) & ( n17928 )  ;
assign n19078 =  ( n84 ) & ( n17930 )  ;
assign n19079 =  ( n84 ) & ( n17932 )  ;
assign n19080 =  ( n85 ) & ( n17902 )  ;
assign n19081 =  ( n85 ) & ( n17904 )  ;
assign n19082 =  ( n85 ) & ( n17906 )  ;
assign n19083 =  ( n85 ) & ( n17908 )  ;
assign n19084 =  ( n85 ) & ( n17910 )  ;
assign n19085 =  ( n85 ) & ( n17912 )  ;
assign n19086 =  ( n85 ) & ( n17914 )  ;
assign n19087 =  ( n85 ) & ( n17916 )  ;
assign n19088 =  ( n85 ) & ( n17918 )  ;
assign n19089 =  ( n85 ) & ( n17920 )  ;
assign n19090 =  ( n85 ) & ( n17922 )  ;
assign n19091 =  ( n85 ) & ( n17924 )  ;
assign n19092 =  ( n85 ) & ( n17926 )  ;
assign n19093 =  ( n85 ) & ( n17928 )  ;
assign n19094 =  ( n85 ) & ( n17930 )  ;
assign n19095 =  ( n85 ) & ( n17932 )  ;
assign n19096 =  ( n86 ) & ( n17902 )  ;
assign n19097 =  ( n86 ) & ( n17904 )  ;
assign n19098 =  ( n86 ) & ( n17906 )  ;
assign n19099 =  ( n86 ) & ( n17908 )  ;
assign n19100 =  ( n86 ) & ( n17910 )  ;
assign n19101 =  ( n86 ) & ( n17912 )  ;
assign n19102 =  ( n86 ) & ( n17914 )  ;
assign n19103 =  ( n86 ) & ( n17916 )  ;
assign n19104 =  ( n86 ) & ( n17918 )  ;
assign n19105 =  ( n86 ) & ( n17920 )  ;
assign n19106 =  ( n86 ) & ( n17922 )  ;
assign n19107 =  ( n86 ) & ( n17924 )  ;
assign n19108 =  ( n86 ) & ( n17926 )  ;
assign n19109 =  ( n86 ) & ( n17928 )  ;
assign n19110 =  ( n86 ) & ( n17930 )  ;
assign n19111 =  ( n86 ) & ( n17932 )  ;
assign n19112 =  ( n87 ) & ( n17902 )  ;
assign n19113 =  ( n87 ) & ( n17904 )  ;
assign n19114 =  ( n87 ) & ( n17906 )  ;
assign n19115 =  ( n87 ) & ( n17908 )  ;
assign n19116 =  ( n87 ) & ( n17910 )  ;
assign n19117 =  ( n87 ) & ( n17912 )  ;
assign n19118 =  ( n87 ) & ( n17914 )  ;
assign n19119 =  ( n87 ) & ( n17916 )  ;
assign n19120 =  ( n87 ) & ( n17918 )  ;
assign n19121 =  ( n87 ) & ( n17920 )  ;
assign n19122 =  ( n87 ) & ( n17922 )  ;
assign n19123 =  ( n87 ) & ( n17924 )  ;
assign n19124 =  ( n87 ) & ( n17926 )  ;
assign n19125 =  ( n87 ) & ( n17928 )  ;
assign n19126 =  ( n87 ) & ( n17930 )  ;
assign n19127 =  ( n87 ) & ( n17932 )  ;
assign n19128 =  ( n88 ) & ( n17902 )  ;
assign n19129 =  ( n88 ) & ( n17904 )  ;
assign n19130 =  ( n88 ) & ( n17906 )  ;
assign n19131 =  ( n88 ) & ( n17908 )  ;
assign n19132 =  ( n88 ) & ( n17910 )  ;
assign n19133 =  ( n88 ) & ( n17912 )  ;
assign n19134 =  ( n88 ) & ( n17914 )  ;
assign n19135 =  ( n88 ) & ( n17916 )  ;
assign n19136 =  ( n88 ) & ( n17918 )  ;
assign n19137 =  ( n88 ) & ( n17920 )  ;
assign n19138 =  ( n88 ) & ( n17922 )  ;
assign n19139 =  ( n88 ) & ( n17924 )  ;
assign n19140 =  ( n88 ) & ( n17926 )  ;
assign n19141 =  ( n88 ) & ( n17928 )  ;
assign n19142 =  ( n88 ) & ( n17930 )  ;
assign n19143 =  ( n88 ) & ( n17932 )  ;
assign n19144 =  ( n89 ) & ( n17902 )  ;
assign n19145 =  ( n89 ) & ( n17904 )  ;
assign n19146 =  ( n89 ) & ( n17906 )  ;
assign n19147 =  ( n89 ) & ( n17908 )  ;
assign n19148 =  ( n89 ) & ( n17910 )  ;
assign n19149 =  ( n89 ) & ( n17912 )  ;
assign n19150 =  ( n89 ) & ( n17914 )  ;
assign n19151 =  ( n89 ) & ( n17916 )  ;
assign n19152 =  ( n89 ) & ( n17918 )  ;
assign n19153 =  ( n89 ) & ( n17920 )  ;
assign n19154 =  ( n89 ) & ( n17922 )  ;
assign n19155 =  ( n89 ) & ( n17924 )  ;
assign n19156 =  ( n89 ) & ( n17926 )  ;
assign n19157 =  ( n89 ) & ( n17928 )  ;
assign n19158 =  ( n89 ) & ( n17930 )  ;
assign n19159 =  ( n89 ) & ( n17932 )  ;
assign n19160 =  ( n90 ) & ( n17902 )  ;
assign n19161 =  ( n90 ) & ( n17904 )  ;
assign n19162 =  ( n90 ) & ( n17906 )  ;
assign n19163 =  ( n90 ) & ( n17908 )  ;
assign n19164 =  ( n90 ) & ( n17910 )  ;
assign n19165 =  ( n90 ) & ( n17912 )  ;
assign n19166 =  ( n90 ) & ( n17914 )  ;
assign n19167 =  ( n90 ) & ( n17916 )  ;
assign n19168 =  ( n90 ) & ( n17918 )  ;
assign n19169 =  ( n90 ) & ( n17920 )  ;
assign n19170 =  ( n90 ) & ( n17922 )  ;
assign n19171 =  ( n90 ) & ( n17924 )  ;
assign n19172 =  ( n90 ) & ( n17926 )  ;
assign n19173 =  ( n90 ) & ( n17928 )  ;
assign n19174 =  ( n90 ) & ( n17930 )  ;
assign n19175 =  ( n90 ) & ( n17932 )  ;
assign n19176 =  ( n91 ) & ( n17902 )  ;
assign n19177 =  ( n91 ) & ( n17904 )  ;
assign n19178 =  ( n91 ) & ( n17906 )  ;
assign n19179 =  ( n91 ) & ( n17908 )  ;
assign n19180 =  ( n91 ) & ( n17910 )  ;
assign n19181 =  ( n91 ) & ( n17912 )  ;
assign n19182 =  ( n91 ) & ( n17914 )  ;
assign n19183 =  ( n91 ) & ( n17916 )  ;
assign n19184 =  ( n91 ) & ( n17918 )  ;
assign n19185 =  ( n91 ) & ( n17920 )  ;
assign n19186 =  ( n91 ) & ( n17922 )  ;
assign n19187 =  ( n91 ) & ( n17924 )  ;
assign n19188 =  ( n91 ) & ( n17926 )  ;
assign n19189 =  ( n91 ) & ( n17928 )  ;
assign n19190 =  ( n91 ) & ( n17930 )  ;
assign n19191 =  ( n91 ) & ( n17932 )  ;
assign n19192 =  ( n92 ) & ( n17902 )  ;
assign n19193 =  ( n92 ) & ( n17904 )  ;
assign n19194 =  ( n92 ) & ( n17906 )  ;
assign n19195 =  ( n92 ) & ( n17908 )  ;
assign n19196 =  ( n92 ) & ( n17910 )  ;
assign n19197 =  ( n92 ) & ( n17912 )  ;
assign n19198 =  ( n92 ) & ( n17914 )  ;
assign n19199 =  ( n92 ) & ( n17916 )  ;
assign n19200 =  ( n92 ) & ( n17918 )  ;
assign n19201 =  ( n92 ) & ( n17920 )  ;
assign n19202 =  ( n92 ) & ( n17922 )  ;
assign n19203 =  ( n92 ) & ( n17924 )  ;
assign n19204 =  ( n92 ) & ( n17926 )  ;
assign n19205 =  ( n92 ) & ( n17928 )  ;
assign n19206 =  ( n92 ) & ( n17930 )  ;
assign n19207 =  ( n92 ) & ( n17932 )  ;
assign n19208 =  ( n93 ) & ( n17902 )  ;
assign n19209 =  ( n93 ) & ( n17904 )  ;
assign n19210 =  ( n93 ) & ( n17906 )  ;
assign n19211 =  ( n93 ) & ( n17908 )  ;
assign n19212 =  ( n93 ) & ( n17910 )  ;
assign n19213 =  ( n93 ) & ( n17912 )  ;
assign n19214 =  ( n93 ) & ( n17914 )  ;
assign n19215 =  ( n93 ) & ( n17916 )  ;
assign n19216 =  ( n93 ) & ( n17918 )  ;
assign n19217 =  ( n93 ) & ( n17920 )  ;
assign n19218 =  ( n93 ) & ( n17922 )  ;
assign n19219 =  ( n93 ) & ( n17924 )  ;
assign n19220 =  ( n93 ) & ( n17926 )  ;
assign n19221 =  ( n93 ) & ( n17928 )  ;
assign n19222 =  ( n93 ) & ( n17930 )  ;
assign n19223 =  ( n93 ) & ( n17932 )  ;
assign n19224 =  ( n94 ) & ( n17902 )  ;
assign n19225 =  ( n94 ) & ( n17904 )  ;
assign n19226 =  ( n94 ) & ( n17906 )  ;
assign n19227 =  ( n94 ) & ( n17908 )  ;
assign n19228 =  ( n94 ) & ( n17910 )  ;
assign n19229 =  ( n94 ) & ( n17912 )  ;
assign n19230 =  ( n94 ) & ( n17914 )  ;
assign n19231 =  ( n94 ) & ( n17916 )  ;
assign n19232 =  ( n94 ) & ( n17918 )  ;
assign n19233 =  ( n94 ) & ( n17920 )  ;
assign n19234 =  ( n94 ) & ( n17922 )  ;
assign n19235 =  ( n94 ) & ( n17924 )  ;
assign n19236 =  ( n94 ) & ( n17926 )  ;
assign n19237 =  ( n94 ) & ( n17928 )  ;
assign n19238 =  ( n94 ) & ( n17930 )  ;
assign n19239 =  ( n94 ) & ( n17932 )  ;
assign n19240 =  ( n95 ) & ( n17902 )  ;
assign n19241 =  ( n95 ) & ( n17904 )  ;
assign n19242 =  ( n95 ) & ( n17906 )  ;
assign n19243 =  ( n95 ) & ( n17908 )  ;
assign n19244 =  ( n95 ) & ( n17910 )  ;
assign n19245 =  ( n95 ) & ( n17912 )  ;
assign n19246 =  ( n95 ) & ( n17914 )  ;
assign n19247 =  ( n95 ) & ( n17916 )  ;
assign n19248 =  ( n95 ) & ( n17918 )  ;
assign n19249 =  ( n95 ) & ( n17920 )  ;
assign n19250 =  ( n95 ) & ( n17922 )  ;
assign n19251 =  ( n95 ) & ( n17924 )  ;
assign n19252 =  ( n95 ) & ( n17926 )  ;
assign n19253 =  ( n95 ) & ( n17928 )  ;
assign n19254 =  ( n95 ) & ( n17930 )  ;
assign n19255 =  ( n95 ) & ( n17932 )  ;
assign n19256 =  ( n96 ) & ( n17902 )  ;
assign n19257 =  ( n96 ) & ( n17904 )  ;
assign n19258 =  ( n96 ) & ( n17906 )  ;
assign n19259 =  ( n96 ) & ( n17908 )  ;
assign n19260 =  ( n96 ) & ( n17910 )  ;
assign n19261 =  ( n96 ) & ( n17912 )  ;
assign n19262 =  ( n96 ) & ( n17914 )  ;
assign n19263 =  ( n96 ) & ( n17916 )  ;
assign n19264 =  ( n96 ) & ( n17918 )  ;
assign n19265 =  ( n96 ) & ( n17920 )  ;
assign n19266 =  ( n96 ) & ( n17922 )  ;
assign n19267 =  ( n96 ) & ( n17924 )  ;
assign n19268 =  ( n96 ) & ( n17926 )  ;
assign n19269 =  ( n96 ) & ( n17928 )  ;
assign n19270 =  ( n96 ) & ( n17930 )  ;
assign n19271 =  ( n96 ) & ( n17932 )  ;
assign n19272 =  ( n97 ) & ( n17902 )  ;
assign n19273 =  ( n97 ) & ( n17904 )  ;
assign n19274 =  ( n97 ) & ( n17906 )  ;
assign n19275 =  ( n97 ) & ( n17908 )  ;
assign n19276 =  ( n97 ) & ( n17910 )  ;
assign n19277 =  ( n97 ) & ( n17912 )  ;
assign n19278 =  ( n97 ) & ( n17914 )  ;
assign n19279 =  ( n97 ) & ( n17916 )  ;
assign n19280 =  ( n97 ) & ( n17918 )  ;
assign n19281 =  ( n97 ) & ( n17920 )  ;
assign n19282 =  ( n97 ) & ( n17922 )  ;
assign n19283 =  ( n97 ) & ( n17924 )  ;
assign n19284 =  ( n97 ) & ( n17926 )  ;
assign n19285 =  ( n97 ) & ( n17928 )  ;
assign n19286 =  ( n97 ) & ( n17930 )  ;
assign n19287 =  ( n97 ) & ( n17932 )  ;
assign n19288 =  ( n98 ) & ( n17902 )  ;
assign n19289 =  ( n98 ) & ( n17904 )  ;
assign n19290 =  ( n98 ) & ( n17906 )  ;
assign n19291 =  ( n98 ) & ( n17908 )  ;
assign n19292 =  ( n98 ) & ( n17910 )  ;
assign n19293 =  ( n98 ) & ( n17912 )  ;
assign n19294 =  ( n98 ) & ( n17914 )  ;
assign n19295 =  ( n98 ) & ( n17916 )  ;
assign n19296 =  ( n98 ) & ( n17918 )  ;
assign n19297 =  ( n98 ) & ( n17920 )  ;
assign n19298 =  ( n98 ) & ( n17922 )  ;
assign n19299 =  ( n98 ) & ( n17924 )  ;
assign n19300 =  ( n98 ) & ( n17926 )  ;
assign n19301 =  ( n98 ) & ( n17928 )  ;
assign n19302 =  ( n98 ) & ( n17930 )  ;
assign n19303 =  ( n98 ) & ( n17932 )  ;
assign n19304 =  ( n99 ) & ( n17902 )  ;
assign n19305 =  ( n99 ) & ( n17904 )  ;
assign n19306 =  ( n99 ) & ( n17906 )  ;
assign n19307 =  ( n99 ) & ( n17908 )  ;
assign n19308 =  ( n99 ) & ( n17910 )  ;
assign n19309 =  ( n99 ) & ( n17912 )  ;
assign n19310 =  ( n99 ) & ( n17914 )  ;
assign n19311 =  ( n99 ) & ( n17916 )  ;
assign n19312 =  ( n99 ) & ( n17918 )  ;
assign n19313 =  ( n99 ) & ( n17920 )  ;
assign n19314 =  ( n99 ) & ( n17922 )  ;
assign n19315 =  ( n99 ) & ( n17924 )  ;
assign n19316 =  ( n99 ) & ( n17926 )  ;
assign n19317 =  ( n99 ) & ( n17928 )  ;
assign n19318 =  ( n99 ) & ( n17930 )  ;
assign n19319 =  ( n99 ) & ( n17932 )  ;
assign n19320 =  ( n100 ) & ( n17902 )  ;
assign n19321 =  ( n100 ) & ( n17904 )  ;
assign n19322 =  ( n100 ) & ( n17906 )  ;
assign n19323 =  ( n100 ) & ( n17908 )  ;
assign n19324 =  ( n100 ) & ( n17910 )  ;
assign n19325 =  ( n100 ) & ( n17912 )  ;
assign n19326 =  ( n100 ) & ( n17914 )  ;
assign n19327 =  ( n100 ) & ( n17916 )  ;
assign n19328 =  ( n100 ) & ( n17918 )  ;
assign n19329 =  ( n100 ) & ( n17920 )  ;
assign n19330 =  ( n100 ) & ( n17922 )  ;
assign n19331 =  ( n100 ) & ( n17924 )  ;
assign n19332 =  ( n100 ) & ( n17926 )  ;
assign n19333 =  ( n100 ) & ( n17928 )  ;
assign n19334 =  ( n100 ) & ( n17930 )  ;
assign n19335 =  ( n100 ) & ( n17932 )  ;
assign n19336 =  ( n101 ) & ( n17902 )  ;
assign n19337 =  ( n101 ) & ( n17904 )  ;
assign n19338 =  ( n101 ) & ( n17906 )  ;
assign n19339 =  ( n101 ) & ( n17908 )  ;
assign n19340 =  ( n101 ) & ( n17910 )  ;
assign n19341 =  ( n101 ) & ( n17912 )  ;
assign n19342 =  ( n101 ) & ( n17914 )  ;
assign n19343 =  ( n101 ) & ( n17916 )  ;
assign n19344 =  ( n101 ) & ( n17918 )  ;
assign n19345 =  ( n101 ) & ( n17920 )  ;
assign n19346 =  ( n101 ) & ( n17922 )  ;
assign n19347 =  ( n101 ) & ( n17924 )  ;
assign n19348 =  ( n101 ) & ( n17926 )  ;
assign n19349 =  ( n101 ) & ( n17928 )  ;
assign n19350 =  ( n101 ) & ( n17930 )  ;
assign n19351 =  ( n101 ) & ( n17932 )  ;
assign n19352 =  ( n102 ) & ( n17902 )  ;
assign n19353 =  ( n102 ) & ( n17904 )  ;
assign n19354 =  ( n102 ) & ( n17906 )  ;
assign n19355 =  ( n102 ) & ( n17908 )  ;
assign n19356 =  ( n102 ) & ( n17910 )  ;
assign n19357 =  ( n102 ) & ( n17912 )  ;
assign n19358 =  ( n102 ) & ( n17914 )  ;
assign n19359 =  ( n102 ) & ( n17916 )  ;
assign n19360 =  ( n102 ) & ( n17918 )  ;
assign n19361 =  ( n102 ) & ( n17920 )  ;
assign n19362 =  ( n102 ) & ( n17922 )  ;
assign n19363 =  ( n102 ) & ( n17924 )  ;
assign n19364 =  ( n102 ) & ( n17926 )  ;
assign n19365 =  ( n102 ) & ( n17928 )  ;
assign n19366 =  ( n102 ) & ( n17930 )  ;
assign n19367 =  ( n102 ) & ( n17932 )  ;
assign n19368 =  ( n103 ) & ( n17902 )  ;
assign n19369 =  ( n103 ) & ( n17904 )  ;
assign n19370 =  ( n103 ) & ( n17906 )  ;
assign n19371 =  ( n103 ) & ( n17908 )  ;
assign n19372 =  ( n103 ) & ( n17910 )  ;
assign n19373 =  ( n103 ) & ( n17912 )  ;
assign n19374 =  ( n103 ) & ( n17914 )  ;
assign n19375 =  ( n103 ) & ( n17916 )  ;
assign n19376 =  ( n103 ) & ( n17918 )  ;
assign n19377 =  ( n103 ) & ( n17920 )  ;
assign n19378 =  ( n103 ) & ( n17922 )  ;
assign n19379 =  ( n103 ) & ( n17924 )  ;
assign n19380 =  ( n103 ) & ( n17926 )  ;
assign n19381 =  ( n103 ) & ( n17928 )  ;
assign n19382 =  ( n103 ) & ( n17930 )  ;
assign n19383 =  ( n103 ) & ( n17932 )  ;
assign n19384 =  ( n104 ) & ( n17902 )  ;
assign n19385 =  ( n104 ) & ( n17904 )  ;
assign n19386 =  ( n104 ) & ( n17906 )  ;
assign n19387 =  ( n104 ) & ( n17908 )  ;
assign n19388 =  ( n104 ) & ( n17910 )  ;
assign n19389 =  ( n104 ) & ( n17912 )  ;
assign n19390 =  ( n104 ) & ( n17914 )  ;
assign n19391 =  ( n104 ) & ( n17916 )  ;
assign n19392 =  ( n104 ) & ( n17918 )  ;
assign n19393 =  ( n104 ) & ( n17920 )  ;
assign n19394 =  ( n104 ) & ( n17922 )  ;
assign n19395 =  ( n104 ) & ( n17924 )  ;
assign n19396 =  ( n104 ) & ( n17926 )  ;
assign n19397 =  ( n104 ) & ( n17928 )  ;
assign n19398 =  ( n104 ) & ( n17930 )  ;
assign n19399 =  ( n104 ) & ( n17932 )  ;
assign n19400 =  ( n105 ) & ( n17902 )  ;
assign n19401 =  ( n105 ) & ( n17904 )  ;
assign n19402 =  ( n105 ) & ( n17906 )  ;
assign n19403 =  ( n105 ) & ( n17908 )  ;
assign n19404 =  ( n105 ) & ( n17910 )  ;
assign n19405 =  ( n105 ) & ( n17912 )  ;
assign n19406 =  ( n105 ) & ( n17914 )  ;
assign n19407 =  ( n105 ) & ( n17916 )  ;
assign n19408 =  ( n105 ) & ( n17918 )  ;
assign n19409 =  ( n105 ) & ( n17920 )  ;
assign n19410 =  ( n105 ) & ( n17922 )  ;
assign n19411 =  ( n105 ) & ( n17924 )  ;
assign n19412 =  ( n105 ) & ( n17926 )  ;
assign n19413 =  ( n105 ) & ( n17928 )  ;
assign n19414 =  ( n105 ) & ( n17930 )  ;
assign n19415 =  ( n105 ) & ( n17932 )  ;
assign n19416 =  ( n106 ) & ( n17902 )  ;
assign n19417 =  ( n106 ) & ( n17904 )  ;
assign n19418 =  ( n106 ) & ( n17906 )  ;
assign n19419 =  ( n106 ) & ( n17908 )  ;
assign n19420 =  ( n106 ) & ( n17910 )  ;
assign n19421 =  ( n106 ) & ( n17912 )  ;
assign n19422 =  ( n106 ) & ( n17914 )  ;
assign n19423 =  ( n106 ) & ( n17916 )  ;
assign n19424 =  ( n106 ) & ( n17918 )  ;
assign n19425 =  ( n106 ) & ( n17920 )  ;
assign n19426 =  ( n106 ) & ( n17922 )  ;
assign n19427 =  ( n106 ) & ( n17924 )  ;
assign n19428 =  ( n106 ) & ( n17926 )  ;
assign n19429 =  ( n106 ) & ( n17928 )  ;
assign n19430 =  ( n106 ) & ( n17930 )  ;
assign n19431 =  ( n106 ) & ( n17932 )  ;
assign n19432 =  ( n107 ) & ( n17902 )  ;
assign n19433 =  ( n107 ) & ( n17904 )  ;
assign n19434 =  ( n107 ) & ( n17906 )  ;
assign n19435 =  ( n107 ) & ( n17908 )  ;
assign n19436 =  ( n107 ) & ( n17910 )  ;
assign n19437 =  ( n107 ) & ( n17912 )  ;
assign n19438 =  ( n107 ) & ( n17914 )  ;
assign n19439 =  ( n107 ) & ( n17916 )  ;
assign n19440 =  ( n107 ) & ( n17918 )  ;
assign n19441 =  ( n107 ) & ( n17920 )  ;
assign n19442 =  ( n107 ) & ( n17922 )  ;
assign n19443 =  ( n107 ) & ( n17924 )  ;
assign n19444 =  ( n107 ) & ( n17926 )  ;
assign n19445 =  ( n107 ) & ( n17928 )  ;
assign n19446 =  ( n107 ) & ( n17930 )  ;
assign n19447 =  ( n107 ) & ( n17932 )  ;
assign n19448 =  ( n108 ) & ( n17902 )  ;
assign n19449 =  ( n108 ) & ( n17904 )  ;
assign n19450 =  ( n108 ) & ( n17906 )  ;
assign n19451 =  ( n108 ) & ( n17908 )  ;
assign n19452 =  ( n108 ) & ( n17910 )  ;
assign n19453 =  ( n108 ) & ( n17912 )  ;
assign n19454 =  ( n108 ) & ( n17914 )  ;
assign n19455 =  ( n108 ) & ( n17916 )  ;
assign n19456 =  ( n108 ) & ( n17918 )  ;
assign n19457 =  ( n108 ) & ( n17920 )  ;
assign n19458 =  ( n108 ) & ( n17922 )  ;
assign n19459 =  ( n108 ) & ( n17924 )  ;
assign n19460 =  ( n108 ) & ( n17926 )  ;
assign n19461 =  ( n108 ) & ( n17928 )  ;
assign n19462 =  ( n108 ) & ( n17930 )  ;
assign n19463 =  ( n108 ) & ( n17932 )  ;
assign n19464 =  ( n19463 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n19465 =  ( n19462 ) ? ( VREG_0_1 ) : ( n19464 ) ;
assign n19466 =  ( n19461 ) ? ( VREG_0_2 ) : ( n19465 ) ;
assign n19467 =  ( n19460 ) ? ( VREG_0_3 ) : ( n19466 ) ;
assign n19468 =  ( n19459 ) ? ( VREG_0_4 ) : ( n19467 ) ;
assign n19469 =  ( n19458 ) ? ( VREG_0_5 ) : ( n19468 ) ;
assign n19470 =  ( n19457 ) ? ( VREG_0_6 ) : ( n19469 ) ;
assign n19471 =  ( n19456 ) ? ( VREG_0_7 ) : ( n19470 ) ;
assign n19472 =  ( n19455 ) ? ( VREG_0_8 ) : ( n19471 ) ;
assign n19473 =  ( n19454 ) ? ( VREG_0_9 ) : ( n19472 ) ;
assign n19474 =  ( n19453 ) ? ( VREG_0_10 ) : ( n19473 ) ;
assign n19475 =  ( n19452 ) ? ( VREG_0_11 ) : ( n19474 ) ;
assign n19476 =  ( n19451 ) ? ( VREG_0_12 ) : ( n19475 ) ;
assign n19477 =  ( n19450 ) ? ( VREG_0_13 ) : ( n19476 ) ;
assign n19478 =  ( n19449 ) ? ( VREG_0_14 ) : ( n19477 ) ;
assign n19479 =  ( n19448 ) ? ( VREG_0_15 ) : ( n19478 ) ;
assign n19480 =  ( n19447 ) ? ( VREG_1_0 ) : ( n19479 ) ;
assign n19481 =  ( n19446 ) ? ( VREG_1_1 ) : ( n19480 ) ;
assign n19482 =  ( n19445 ) ? ( VREG_1_2 ) : ( n19481 ) ;
assign n19483 =  ( n19444 ) ? ( VREG_1_3 ) : ( n19482 ) ;
assign n19484 =  ( n19443 ) ? ( VREG_1_4 ) : ( n19483 ) ;
assign n19485 =  ( n19442 ) ? ( VREG_1_5 ) : ( n19484 ) ;
assign n19486 =  ( n19441 ) ? ( VREG_1_6 ) : ( n19485 ) ;
assign n19487 =  ( n19440 ) ? ( VREG_1_7 ) : ( n19486 ) ;
assign n19488 =  ( n19439 ) ? ( VREG_1_8 ) : ( n19487 ) ;
assign n19489 =  ( n19438 ) ? ( VREG_1_9 ) : ( n19488 ) ;
assign n19490 =  ( n19437 ) ? ( VREG_1_10 ) : ( n19489 ) ;
assign n19491 =  ( n19436 ) ? ( VREG_1_11 ) : ( n19490 ) ;
assign n19492 =  ( n19435 ) ? ( VREG_1_12 ) : ( n19491 ) ;
assign n19493 =  ( n19434 ) ? ( VREG_1_13 ) : ( n19492 ) ;
assign n19494 =  ( n19433 ) ? ( VREG_1_14 ) : ( n19493 ) ;
assign n19495 =  ( n19432 ) ? ( VREG_1_15 ) : ( n19494 ) ;
assign n19496 =  ( n19431 ) ? ( VREG_2_0 ) : ( n19495 ) ;
assign n19497 =  ( n19430 ) ? ( VREG_2_1 ) : ( n19496 ) ;
assign n19498 =  ( n19429 ) ? ( VREG_2_2 ) : ( n19497 ) ;
assign n19499 =  ( n19428 ) ? ( VREG_2_3 ) : ( n19498 ) ;
assign n19500 =  ( n19427 ) ? ( VREG_2_4 ) : ( n19499 ) ;
assign n19501 =  ( n19426 ) ? ( VREG_2_5 ) : ( n19500 ) ;
assign n19502 =  ( n19425 ) ? ( VREG_2_6 ) : ( n19501 ) ;
assign n19503 =  ( n19424 ) ? ( VREG_2_7 ) : ( n19502 ) ;
assign n19504 =  ( n19423 ) ? ( VREG_2_8 ) : ( n19503 ) ;
assign n19505 =  ( n19422 ) ? ( VREG_2_9 ) : ( n19504 ) ;
assign n19506 =  ( n19421 ) ? ( VREG_2_10 ) : ( n19505 ) ;
assign n19507 =  ( n19420 ) ? ( VREG_2_11 ) : ( n19506 ) ;
assign n19508 =  ( n19419 ) ? ( VREG_2_12 ) : ( n19507 ) ;
assign n19509 =  ( n19418 ) ? ( VREG_2_13 ) : ( n19508 ) ;
assign n19510 =  ( n19417 ) ? ( VREG_2_14 ) : ( n19509 ) ;
assign n19511 =  ( n19416 ) ? ( VREG_2_15 ) : ( n19510 ) ;
assign n19512 =  ( n19415 ) ? ( VREG_3_0 ) : ( n19511 ) ;
assign n19513 =  ( n19414 ) ? ( VREG_3_1 ) : ( n19512 ) ;
assign n19514 =  ( n19413 ) ? ( VREG_3_2 ) : ( n19513 ) ;
assign n19515 =  ( n19412 ) ? ( VREG_3_3 ) : ( n19514 ) ;
assign n19516 =  ( n19411 ) ? ( VREG_3_4 ) : ( n19515 ) ;
assign n19517 =  ( n19410 ) ? ( VREG_3_5 ) : ( n19516 ) ;
assign n19518 =  ( n19409 ) ? ( VREG_3_6 ) : ( n19517 ) ;
assign n19519 =  ( n19408 ) ? ( VREG_3_7 ) : ( n19518 ) ;
assign n19520 =  ( n19407 ) ? ( VREG_3_8 ) : ( n19519 ) ;
assign n19521 =  ( n19406 ) ? ( VREG_3_9 ) : ( n19520 ) ;
assign n19522 =  ( n19405 ) ? ( VREG_3_10 ) : ( n19521 ) ;
assign n19523 =  ( n19404 ) ? ( VREG_3_11 ) : ( n19522 ) ;
assign n19524 =  ( n19403 ) ? ( VREG_3_12 ) : ( n19523 ) ;
assign n19525 =  ( n19402 ) ? ( VREG_3_13 ) : ( n19524 ) ;
assign n19526 =  ( n19401 ) ? ( VREG_3_14 ) : ( n19525 ) ;
assign n19527 =  ( n19400 ) ? ( VREG_3_15 ) : ( n19526 ) ;
assign n19528 =  ( n19399 ) ? ( VREG_4_0 ) : ( n19527 ) ;
assign n19529 =  ( n19398 ) ? ( VREG_4_1 ) : ( n19528 ) ;
assign n19530 =  ( n19397 ) ? ( VREG_4_2 ) : ( n19529 ) ;
assign n19531 =  ( n19396 ) ? ( VREG_4_3 ) : ( n19530 ) ;
assign n19532 =  ( n19395 ) ? ( VREG_4_4 ) : ( n19531 ) ;
assign n19533 =  ( n19394 ) ? ( VREG_4_5 ) : ( n19532 ) ;
assign n19534 =  ( n19393 ) ? ( VREG_4_6 ) : ( n19533 ) ;
assign n19535 =  ( n19392 ) ? ( VREG_4_7 ) : ( n19534 ) ;
assign n19536 =  ( n19391 ) ? ( VREG_4_8 ) : ( n19535 ) ;
assign n19537 =  ( n19390 ) ? ( VREG_4_9 ) : ( n19536 ) ;
assign n19538 =  ( n19389 ) ? ( VREG_4_10 ) : ( n19537 ) ;
assign n19539 =  ( n19388 ) ? ( VREG_4_11 ) : ( n19538 ) ;
assign n19540 =  ( n19387 ) ? ( VREG_4_12 ) : ( n19539 ) ;
assign n19541 =  ( n19386 ) ? ( VREG_4_13 ) : ( n19540 ) ;
assign n19542 =  ( n19385 ) ? ( VREG_4_14 ) : ( n19541 ) ;
assign n19543 =  ( n19384 ) ? ( VREG_4_15 ) : ( n19542 ) ;
assign n19544 =  ( n19383 ) ? ( VREG_5_0 ) : ( n19543 ) ;
assign n19545 =  ( n19382 ) ? ( VREG_5_1 ) : ( n19544 ) ;
assign n19546 =  ( n19381 ) ? ( VREG_5_2 ) : ( n19545 ) ;
assign n19547 =  ( n19380 ) ? ( VREG_5_3 ) : ( n19546 ) ;
assign n19548 =  ( n19379 ) ? ( VREG_5_4 ) : ( n19547 ) ;
assign n19549 =  ( n19378 ) ? ( VREG_5_5 ) : ( n19548 ) ;
assign n19550 =  ( n19377 ) ? ( VREG_5_6 ) : ( n19549 ) ;
assign n19551 =  ( n19376 ) ? ( VREG_5_7 ) : ( n19550 ) ;
assign n19552 =  ( n19375 ) ? ( VREG_5_8 ) : ( n19551 ) ;
assign n19553 =  ( n19374 ) ? ( VREG_5_9 ) : ( n19552 ) ;
assign n19554 =  ( n19373 ) ? ( VREG_5_10 ) : ( n19553 ) ;
assign n19555 =  ( n19372 ) ? ( VREG_5_11 ) : ( n19554 ) ;
assign n19556 =  ( n19371 ) ? ( VREG_5_12 ) : ( n19555 ) ;
assign n19557 =  ( n19370 ) ? ( VREG_5_13 ) : ( n19556 ) ;
assign n19558 =  ( n19369 ) ? ( VREG_5_14 ) : ( n19557 ) ;
assign n19559 =  ( n19368 ) ? ( VREG_5_15 ) : ( n19558 ) ;
assign n19560 =  ( n19367 ) ? ( VREG_6_0 ) : ( n19559 ) ;
assign n19561 =  ( n19366 ) ? ( VREG_6_1 ) : ( n19560 ) ;
assign n19562 =  ( n19365 ) ? ( VREG_6_2 ) : ( n19561 ) ;
assign n19563 =  ( n19364 ) ? ( VREG_6_3 ) : ( n19562 ) ;
assign n19564 =  ( n19363 ) ? ( VREG_6_4 ) : ( n19563 ) ;
assign n19565 =  ( n19362 ) ? ( VREG_6_5 ) : ( n19564 ) ;
assign n19566 =  ( n19361 ) ? ( VREG_6_6 ) : ( n19565 ) ;
assign n19567 =  ( n19360 ) ? ( VREG_6_7 ) : ( n19566 ) ;
assign n19568 =  ( n19359 ) ? ( VREG_6_8 ) : ( n19567 ) ;
assign n19569 =  ( n19358 ) ? ( VREG_6_9 ) : ( n19568 ) ;
assign n19570 =  ( n19357 ) ? ( VREG_6_10 ) : ( n19569 ) ;
assign n19571 =  ( n19356 ) ? ( VREG_6_11 ) : ( n19570 ) ;
assign n19572 =  ( n19355 ) ? ( VREG_6_12 ) : ( n19571 ) ;
assign n19573 =  ( n19354 ) ? ( VREG_6_13 ) : ( n19572 ) ;
assign n19574 =  ( n19353 ) ? ( VREG_6_14 ) : ( n19573 ) ;
assign n19575 =  ( n19352 ) ? ( VREG_6_15 ) : ( n19574 ) ;
assign n19576 =  ( n19351 ) ? ( VREG_7_0 ) : ( n19575 ) ;
assign n19577 =  ( n19350 ) ? ( VREG_7_1 ) : ( n19576 ) ;
assign n19578 =  ( n19349 ) ? ( VREG_7_2 ) : ( n19577 ) ;
assign n19579 =  ( n19348 ) ? ( VREG_7_3 ) : ( n19578 ) ;
assign n19580 =  ( n19347 ) ? ( VREG_7_4 ) : ( n19579 ) ;
assign n19581 =  ( n19346 ) ? ( VREG_7_5 ) : ( n19580 ) ;
assign n19582 =  ( n19345 ) ? ( VREG_7_6 ) : ( n19581 ) ;
assign n19583 =  ( n19344 ) ? ( VREG_7_7 ) : ( n19582 ) ;
assign n19584 =  ( n19343 ) ? ( VREG_7_8 ) : ( n19583 ) ;
assign n19585 =  ( n19342 ) ? ( VREG_7_9 ) : ( n19584 ) ;
assign n19586 =  ( n19341 ) ? ( VREG_7_10 ) : ( n19585 ) ;
assign n19587 =  ( n19340 ) ? ( VREG_7_11 ) : ( n19586 ) ;
assign n19588 =  ( n19339 ) ? ( VREG_7_12 ) : ( n19587 ) ;
assign n19589 =  ( n19338 ) ? ( VREG_7_13 ) : ( n19588 ) ;
assign n19590 =  ( n19337 ) ? ( VREG_7_14 ) : ( n19589 ) ;
assign n19591 =  ( n19336 ) ? ( VREG_7_15 ) : ( n19590 ) ;
assign n19592 =  ( n19335 ) ? ( VREG_8_0 ) : ( n19591 ) ;
assign n19593 =  ( n19334 ) ? ( VREG_8_1 ) : ( n19592 ) ;
assign n19594 =  ( n19333 ) ? ( VREG_8_2 ) : ( n19593 ) ;
assign n19595 =  ( n19332 ) ? ( VREG_8_3 ) : ( n19594 ) ;
assign n19596 =  ( n19331 ) ? ( VREG_8_4 ) : ( n19595 ) ;
assign n19597 =  ( n19330 ) ? ( VREG_8_5 ) : ( n19596 ) ;
assign n19598 =  ( n19329 ) ? ( VREG_8_6 ) : ( n19597 ) ;
assign n19599 =  ( n19328 ) ? ( VREG_8_7 ) : ( n19598 ) ;
assign n19600 =  ( n19327 ) ? ( VREG_8_8 ) : ( n19599 ) ;
assign n19601 =  ( n19326 ) ? ( VREG_8_9 ) : ( n19600 ) ;
assign n19602 =  ( n19325 ) ? ( VREG_8_10 ) : ( n19601 ) ;
assign n19603 =  ( n19324 ) ? ( VREG_8_11 ) : ( n19602 ) ;
assign n19604 =  ( n19323 ) ? ( VREG_8_12 ) : ( n19603 ) ;
assign n19605 =  ( n19322 ) ? ( VREG_8_13 ) : ( n19604 ) ;
assign n19606 =  ( n19321 ) ? ( VREG_8_14 ) : ( n19605 ) ;
assign n19607 =  ( n19320 ) ? ( VREG_8_15 ) : ( n19606 ) ;
assign n19608 =  ( n19319 ) ? ( VREG_9_0 ) : ( n19607 ) ;
assign n19609 =  ( n19318 ) ? ( VREG_9_1 ) : ( n19608 ) ;
assign n19610 =  ( n19317 ) ? ( VREG_9_2 ) : ( n19609 ) ;
assign n19611 =  ( n19316 ) ? ( VREG_9_3 ) : ( n19610 ) ;
assign n19612 =  ( n19315 ) ? ( VREG_9_4 ) : ( n19611 ) ;
assign n19613 =  ( n19314 ) ? ( VREG_9_5 ) : ( n19612 ) ;
assign n19614 =  ( n19313 ) ? ( VREG_9_6 ) : ( n19613 ) ;
assign n19615 =  ( n19312 ) ? ( VREG_9_7 ) : ( n19614 ) ;
assign n19616 =  ( n19311 ) ? ( VREG_9_8 ) : ( n19615 ) ;
assign n19617 =  ( n19310 ) ? ( VREG_9_9 ) : ( n19616 ) ;
assign n19618 =  ( n19309 ) ? ( VREG_9_10 ) : ( n19617 ) ;
assign n19619 =  ( n19308 ) ? ( VREG_9_11 ) : ( n19618 ) ;
assign n19620 =  ( n19307 ) ? ( VREG_9_12 ) : ( n19619 ) ;
assign n19621 =  ( n19306 ) ? ( VREG_9_13 ) : ( n19620 ) ;
assign n19622 =  ( n19305 ) ? ( VREG_9_14 ) : ( n19621 ) ;
assign n19623 =  ( n19304 ) ? ( VREG_9_15 ) : ( n19622 ) ;
assign n19624 =  ( n19303 ) ? ( VREG_10_0 ) : ( n19623 ) ;
assign n19625 =  ( n19302 ) ? ( VREG_10_1 ) : ( n19624 ) ;
assign n19626 =  ( n19301 ) ? ( VREG_10_2 ) : ( n19625 ) ;
assign n19627 =  ( n19300 ) ? ( VREG_10_3 ) : ( n19626 ) ;
assign n19628 =  ( n19299 ) ? ( VREG_10_4 ) : ( n19627 ) ;
assign n19629 =  ( n19298 ) ? ( VREG_10_5 ) : ( n19628 ) ;
assign n19630 =  ( n19297 ) ? ( VREG_10_6 ) : ( n19629 ) ;
assign n19631 =  ( n19296 ) ? ( VREG_10_7 ) : ( n19630 ) ;
assign n19632 =  ( n19295 ) ? ( VREG_10_8 ) : ( n19631 ) ;
assign n19633 =  ( n19294 ) ? ( VREG_10_9 ) : ( n19632 ) ;
assign n19634 =  ( n19293 ) ? ( VREG_10_10 ) : ( n19633 ) ;
assign n19635 =  ( n19292 ) ? ( VREG_10_11 ) : ( n19634 ) ;
assign n19636 =  ( n19291 ) ? ( VREG_10_12 ) : ( n19635 ) ;
assign n19637 =  ( n19290 ) ? ( VREG_10_13 ) : ( n19636 ) ;
assign n19638 =  ( n19289 ) ? ( VREG_10_14 ) : ( n19637 ) ;
assign n19639 =  ( n19288 ) ? ( VREG_10_15 ) : ( n19638 ) ;
assign n19640 =  ( n19287 ) ? ( VREG_11_0 ) : ( n19639 ) ;
assign n19641 =  ( n19286 ) ? ( VREG_11_1 ) : ( n19640 ) ;
assign n19642 =  ( n19285 ) ? ( VREG_11_2 ) : ( n19641 ) ;
assign n19643 =  ( n19284 ) ? ( VREG_11_3 ) : ( n19642 ) ;
assign n19644 =  ( n19283 ) ? ( VREG_11_4 ) : ( n19643 ) ;
assign n19645 =  ( n19282 ) ? ( VREG_11_5 ) : ( n19644 ) ;
assign n19646 =  ( n19281 ) ? ( VREG_11_6 ) : ( n19645 ) ;
assign n19647 =  ( n19280 ) ? ( VREG_11_7 ) : ( n19646 ) ;
assign n19648 =  ( n19279 ) ? ( VREG_11_8 ) : ( n19647 ) ;
assign n19649 =  ( n19278 ) ? ( VREG_11_9 ) : ( n19648 ) ;
assign n19650 =  ( n19277 ) ? ( VREG_11_10 ) : ( n19649 ) ;
assign n19651 =  ( n19276 ) ? ( VREG_11_11 ) : ( n19650 ) ;
assign n19652 =  ( n19275 ) ? ( VREG_11_12 ) : ( n19651 ) ;
assign n19653 =  ( n19274 ) ? ( VREG_11_13 ) : ( n19652 ) ;
assign n19654 =  ( n19273 ) ? ( VREG_11_14 ) : ( n19653 ) ;
assign n19655 =  ( n19272 ) ? ( VREG_11_15 ) : ( n19654 ) ;
assign n19656 =  ( n19271 ) ? ( VREG_12_0 ) : ( n19655 ) ;
assign n19657 =  ( n19270 ) ? ( VREG_12_1 ) : ( n19656 ) ;
assign n19658 =  ( n19269 ) ? ( VREG_12_2 ) : ( n19657 ) ;
assign n19659 =  ( n19268 ) ? ( VREG_12_3 ) : ( n19658 ) ;
assign n19660 =  ( n19267 ) ? ( VREG_12_4 ) : ( n19659 ) ;
assign n19661 =  ( n19266 ) ? ( VREG_12_5 ) : ( n19660 ) ;
assign n19662 =  ( n19265 ) ? ( VREG_12_6 ) : ( n19661 ) ;
assign n19663 =  ( n19264 ) ? ( VREG_12_7 ) : ( n19662 ) ;
assign n19664 =  ( n19263 ) ? ( VREG_12_8 ) : ( n19663 ) ;
assign n19665 =  ( n19262 ) ? ( VREG_12_9 ) : ( n19664 ) ;
assign n19666 =  ( n19261 ) ? ( VREG_12_10 ) : ( n19665 ) ;
assign n19667 =  ( n19260 ) ? ( VREG_12_11 ) : ( n19666 ) ;
assign n19668 =  ( n19259 ) ? ( VREG_12_12 ) : ( n19667 ) ;
assign n19669 =  ( n19258 ) ? ( VREG_12_13 ) : ( n19668 ) ;
assign n19670 =  ( n19257 ) ? ( VREG_12_14 ) : ( n19669 ) ;
assign n19671 =  ( n19256 ) ? ( VREG_12_15 ) : ( n19670 ) ;
assign n19672 =  ( n19255 ) ? ( VREG_13_0 ) : ( n19671 ) ;
assign n19673 =  ( n19254 ) ? ( VREG_13_1 ) : ( n19672 ) ;
assign n19674 =  ( n19253 ) ? ( VREG_13_2 ) : ( n19673 ) ;
assign n19675 =  ( n19252 ) ? ( VREG_13_3 ) : ( n19674 ) ;
assign n19676 =  ( n19251 ) ? ( VREG_13_4 ) : ( n19675 ) ;
assign n19677 =  ( n19250 ) ? ( VREG_13_5 ) : ( n19676 ) ;
assign n19678 =  ( n19249 ) ? ( VREG_13_6 ) : ( n19677 ) ;
assign n19679 =  ( n19248 ) ? ( VREG_13_7 ) : ( n19678 ) ;
assign n19680 =  ( n19247 ) ? ( VREG_13_8 ) : ( n19679 ) ;
assign n19681 =  ( n19246 ) ? ( VREG_13_9 ) : ( n19680 ) ;
assign n19682 =  ( n19245 ) ? ( VREG_13_10 ) : ( n19681 ) ;
assign n19683 =  ( n19244 ) ? ( VREG_13_11 ) : ( n19682 ) ;
assign n19684 =  ( n19243 ) ? ( VREG_13_12 ) : ( n19683 ) ;
assign n19685 =  ( n19242 ) ? ( VREG_13_13 ) : ( n19684 ) ;
assign n19686 =  ( n19241 ) ? ( VREG_13_14 ) : ( n19685 ) ;
assign n19687 =  ( n19240 ) ? ( VREG_13_15 ) : ( n19686 ) ;
assign n19688 =  ( n19239 ) ? ( VREG_14_0 ) : ( n19687 ) ;
assign n19689 =  ( n19238 ) ? ( VREG_14_1 ) : ( n19688 ) ;
assign n19690 =  ( n19237 ) ? ( VREG_14_2 ) : ( n19689 ) ;
assign n19691 =  ( n19236 ) ? ( VREG_14_3 ) : ( n19690 ) ;
assign n19692 =  ( n19235 ) ? ( VREG_14_4 ) : ( n19691 ) ;
assign n19693 =  ( n19234 ) ? ( VREG_14_5 ) : ( n19692 ) ;
assign n19694 =  ( n19233 ) ? ( VREG_14_6 ) : ( n19693 ) ;
assign n19695 =  ( n19232 ) ? ( VREG_14_7 ) : ( n19694 ) ;
assign n19696 =  ( n19231 ) ? ( VREG_14_8 ) : ( n19695 ) ;
assign n19697 =  ( n19230 ) ? ( VREG_14_9 ) : ( n19696 ) ;
assign n19698 =  ( n19229 ) ? ( VREG_14_10 ) : ( n19697 ) ;
assign n19699 =  ( n19228 ) ? ( VREG_14_11 ) : ( n19698 ) ;
assign n19700 =  ( n19227 ) ? ( VREG_14_12 ) : ( n19699 ) ;
assign n19701 =  ( n19226 ) ? ( VREG_14_13 ) : ( n19700 ) ;
assign n19702 =  ( n19225 ) ? ( VREG_14_14 ) : ( n19701 ) ;
assign n19703 =  ( n19224 ) ? ( VREG_14_15 ) : ( n19702 ) ;
assign n19704 =  ( n19223 ) ? ( VREG_15_0 ) : ( n19703 ) ;
assign n19705 =  ( n19222 ) ? ( VREG_15_1 ) : ( n19704 ) ;
assign n19706 =  ( n19221 ) ? ( VREG_15_2 ) : ( n19705 ) ;
assign n19707 =  ( n19220 ) ? ( VREG_15_3 ) : ( n19706 ) ;
assign n19708 =  ( n19219 ) ? ( VREG_15_4 ) : ( n19707 ) ;
assign n19709 =  ( n19218 ) ? ( VREG_15_5 ) : ( n19708 ) ;
assign n19710 =  ( n19217 ) ? ( VREG_15_6 ) : ( n19709 ) ;
assign n19711 =  ( n19216 ) ? ( VREG_15_7 ) : ( n19710 ) ;
assign n19712 =  ( n19215 ) ? ( VREG_15_8 ) : ( n19711 ) ;
assign n19713 =  ( n19214 ) ? ( VREG_15_9 ) : ( n19712 ) ;
assign n19714 =  ( n19213 ) ? ( VREG_15_10 ) : ( n19713 ) ;
assign n19715 =  ( n19212 ) ? ( VREG_15_11 ) : ( n19714 ) ;
assign n19716 =  ( n19211 ) ? ( VREG_15_12 ) : ( n19715 ) ;
assign n19717 =  ( n19210 ) ? ( VREG_15_13 ) : ( n19716 ) ;
assign n19718 =  ( n19209 ) ? ( VREG_15_14 ) : ( n19717 ) ;
assign n19719 =  ( n19208 ) ? ( VREG_15_15 ) : ( n19718 ) ;
assign n19720 =  ( n19207 ) ? ( VREG_16_0 ) : ( n19719 ) ;
assign n19721 =  ( n19206 ) ? ( VREG_16_1 ) : ( n19720 ) ;
assign n19722 =  ( n19205 ) ? ( VREG_16_2 ) : ( n19721 ) ;
assign n19723 =  ( n19204 ) ? ( VREG_16_3 ) : ( n19722 ) ;
assign n19724 =  ( n19203 ) ? ( VREG_16_4 ) : ( n19723 ) ;
assign n19725 =  ( n19202 ) ? ( VREG_16_5 ) : ( n19724 ) ;
assign n19726 =  ( n19201 ) ? ( VREG_16_6 ) : ( n19725 ) ;
assign n19727 =  ( n19200 ) ? ( VREG_16_7 ) : ( n19726 ) ;
assign n19728 =  ( n19199 ) ? ( VREG_16_8 ) : ( n19727 ) ;
assign n19729 =  ( n19198 ) ? ( VREG_16_9 ) : ( n19728 ) ;
assign n19730 =  ( n19197 ) ? ( VREG_16_10 ) : ( n19729 ) ;
assign n19731 =  ( n19196 ) ? ( VREG_16_11 ) : ( n19730 ) ;
assign n19732 =  ( n19195 ) ? ( VREG_16_12 ) : ( n19731 ) ;
assign n19733 =  ( n19194 ) ? ( VREG_16_13 ) : ( n19732 ) ;
assign n19734 =  ( n19193 ) ? ( VREG_16_14 ) : ( n19733 ) ;
assign n19735 =  ( n19192 ) ? ( VREG_16_15 ) : ( n19734 ) ;
assign n19736 =  ( n19191 ) ? ( VREG_17_0 ) : ( n19735 ) ;
assign n19737 =  ( n19190 ) ? ( VREG_17_1 ) : ( n19736 ) ;
assign n19738 =  ( n19189 ) ? ( VREG_17_2 ) : ( n19737 ) ;
assign n19739 =  ( n19188 ) ? ( VREG_17_3 ) : ( n19738 ) ;
assign n19740 =  ( n19187 ) ? ( VREG_17_4 ) : ( n19739 ) ;
assign n19741 =  ( n19186 ) ? ( VREG_17_5 ) : ( n19740 ) ;
assign n19742 =  ( n19185 ) ? ( VREG_17_6 ) : ( n19741 ) ;
assign n19743 =  ( n19184 ) ? ( VREG_17_7 ) : ( n19742 ) ;
assign n19744 =  ( n19183 ) ? ( VREG_17_8 ) : ( n19743 ) ;
assign n19745 =  ( n19182 ) ? ( VREG_17_9 ) : ( n19744 ) ;
assign n19746 =  ( n19181 ) ? ( VREG_17_10 ) : ( n19745 ) ;
assign n19747 =  ( n19180 ) ? ( VREG_17_11 ) : ( n19746 ) ;
assign n19748 =  ( n19179 ) ? ( VREG_17_12 ) : ( n19747 ) ;
assign n19749 =  ( n19178 ) ? ( VREG_17_13 ) : ( n19748 ) ;
assign n19750 =  ( n19177 ) ? ( VREG_17_14 ) : ( n19749 ) ;
assign n19751 =  ( n19176 ) ? ( VREG_17_15 ) : ( n19750 ) ;
assign n19752 =  ( n19175 ) ? ( VREG_18_0 ) : ( n19751 ) ;
assign n19753 =  ( n19174 ) ? ( VREG_18_1 ) : ( n19752 ) ;
assign n19754 =  ( n19173 ) ? ( VREG_18_2 ) : ( n19753 ) ;
assign n19755 =  ( n19172 ) ? ( VREG_18_3 ) : ( n19754 ) ;
assign n19756 =  ( n19171 ) ? ( VREG_18_4 ) : ( n19755 ) ;
assign n19757 =  ( n19170 ) ? ( VREG_18_5 ) : ( n19756 ) ;
assign n19758 =  ( n19169 ) ? ( VREG_18_6 ) : ( n19757 ) ;
assign n19759 =  ( n19168 ) ? ( VREG_18_7 ) : ( n19758 ) ;
assign n19760 =  ( n19167 ) ? ( VREG_18_8 ) : ( n19759 ) ;
assign n19761 =  ( n19166 ) ? ( VREG_18_9 ) : ( n19760 ) ;
assign n19762 =  ( n19165 ) ? ( VREG_18_10 ) : ( n19761 ) ;
assign n19763 =  ( n19164 ) ? ( VREG_18_11 ) : ( n19762 ) ;
assign n19764 =  ( n19163 ) ? ( VREG_18_12 ) : ( n19763 ) ;
assign n19765 =  ( n19162 ) ? ( VREG_18_13 ) : ( n19764 ) ;
assign n19766 =  ( n19161 ) ? ( VREG_18_14 ) : ( n19765 ) ;
assign n19767 =  ( n19160 ) ? ( VREG_18_15 ) : ( n19766 ) ;
assign n19768 =  ( n19159 ) ? ( VREG_19_0 ) : ( n19767 ) ;
assign n19769 =  ( n19158 ) ? ( VREG_19_1 ) : ( n19768 ) ;
assign n19770 =  ( n19157 ) ? ( VREG_19_2 ) : ( n19769 ) ;
assign n19771 =  ( n19156 ) ? ( VREG_19_3 ) : ( n19770 ) ;
assign n19772 =  ( n19155 ) ? ( VREG_19_4 ) : ( n19771 ) ;
assign n19773 =  ( n19154 ) ? ( VREG_19_5 ) : ( n19772 ) ;
assign n19774 =  ( n19153 ) ? ( VREG_19_6 ) : ( n19773 ) ;
assign n19775 =  ( n19152 ) ? ( VREG_19_7 ) : ( n19774 ) ;
assign n19776 =  ( n19151 ) ? ( VREG_19_8 ) : ( n19775 ) ;
assign n19777 =  ( n19150 ) ? ( VREG_19_9 ) : ( n19776 ) ;
assign n19778 =  ( n19149 ) ? ( VREG_19_10 ) : ( n19777 ) ;
assign n19779 =  ( n19148 ) ? ( VREG_19_11 ) : ( n19778 ) ;
assign n19780 =  ( n19147 ) ? ( VREG_19_12 ) : ( n19779 ) ;
assign n19781 =  ( n19146 ) ? ( VREG_19_13 ) : ( n19780 ) ;
assign n19782 =  ( n19145 ) ? ( VREG_19_14 ) : ( n19781 ) ;
assign n19783 =  ( n19144 ) ? ( VREG_19_15 ) : ( n19782 ) ;
assign n19784 =  ( n19143 ) ? ( VREG_20_0 ) : ( n19783 ) ;
assign n19785 =  ( n19142 ) ? ( VREG_20_1 ) : ( n19784 ) ;
assign n19786 =  ( n19141 ) ? ( VREG_20_2 ) : ( n19785 ) ;
assign n19787 =  ( n19140 ) ? ( VREG_20_3 ) : ( n19786 ) ;
assign n19788 =  ( n19139 ) ? ( VREG_20_4 ) : ( n19787 ) ;
assign n19789 =  ( n19138 ) ? ( VREG_20_5 ) : ( n19788 ) ;
assign n19790 =  ( n19137 ) ? ( VREG_20_6 ) : ( n19789 ) ;
assign n19791 =  ( n19136 ) ? ( VREG_20_7 ) : ( n19790 ) ;
assign n19792 =  ( n19135 ) ? ( VREG_20_8 ) : ( n19791 ) ;
assign n19793 =  ( n19134 ) ? ( VREG_20_9 ) : ( n19792 ) ;
assign n19794 =  ( n19133 ) ? ( VREG_20_10 ) : ( n19793 ) ;
assign n19795 =  ( n19132 ) ? ( VREG_20_11 ) : ( n19794 ) ;
assign n19796 =  ( n19131 ) ? ( VREG_20_12 ) : ( n19795 ) ;
assign n19797 =  ( n19130 ) ? ( VREG_20_13 ) : ( n19796 ) ;
assign n19798 =  ( n19129 ) ? ( VREG_20_14 ) : ( n19797 ) ;
assign n19799 =  ( n19128 ) ? ( VREG_20_15 ) : ( n19798 ) ;
assign n19800 =  ( n19127 ) ? ( VREG_21_0 ) : ( n19799 ) ;
assign n19801 =  ( n19126 ) ? ( VREG_21_1 ) : ( n19800 ) ;
assign n19802 =  ( n19125 ) ? ( VREG_21_2 ) : ( n19801 ) ;
assign n19803 =  ( n19124 ) ? ( VREG_21_3 ) : ( n19802 ) ;
assign n19804 =  ( n19123 ) ? ( VREG_21_4 ) : ( n19803 ) ;
assign n19805 =  ( n19122 ) ? ( VREG_21_5 ) : ( n19804 ) ;
assign n19806 =  ( n19121 ) ? ( VREG_21_6 ) : ( n19805 ) ;
assign n19807 =  ( n19120 ) ? ( VREG_21_7 ) : ( n19806 ) ;
assign n19808 =  ( n19119 ) ? ( VREG_21_8 ) : ( n19807 ) ;
assign n19809 =  ( n19118 ) ? ( VREG_21_9 ) : ( n19808 ) ;
assign n19810 =  ( n19117 ) ? ( VREG_21_10 ) : ( n19809 ) ;
assign n19811 =  ( n19116 ) ? ( VREG_21_11 ) : ( n19810 ) ;
assign n19812 =  ( n19115 ) ? ( VREG_21_12 ) : ( n19811 ) ;
assign n19813 =  ( n19114 ) ? ( VREG_21_13 ) : ( n19812 ) ;
assign n19814 =  ( n19113 ) ? ( VREG_21_14 ) : ( n19813 ) ;
assign n19815 =  ( n19112 ) ? ( VREG_21_15 ) : ( n19814 ) ;
assign n19816 =  ( n19111 ) ? ( VREG_22_0 ) : ( n19815 ) ;
assign n19817 =  ( n19110 ) ? ( VREG_22_1 ) : ( n19816 ) ;
assign n19818 =  ( n19109 ) ? ( VREG_22_2 ) : ( n19817 ) ;
assign n19819 =  ( n19108 ) ? ( VREG_22_3 ) : ( n19818 ) ;
assign n19820 =  ( n19107 ) ? ( VREG_22_4 ) : ( n19819 ) ;
assign n19821 =  ( n19106 ) ? ( VREG_22_5 ) : ( n19820 ) ;
assign n19822 =  ( n19105 ) ? ( VREG_22_6 ) : ( n19821 ) ;
assign n19823 =  ( n19104 ) ? ( VREG_22_7 ) : ( n19822 ) ;
assign n19824 =  ( n19103 ) ? ( VREG_22_8 ) : ( n19823 ) ;
assign n19825 =  ( n19102 ) ? ( VREG_22_9 ) : ( n19824 ) ;
assign n19826 =  ( n19101 ) ? ( VREG_22_10 ) : ( n19825 ) ;
assign n19827 =  ( n19100 ) ? ( VREG_22_11 ) : ( n19826 ) ;
assign n19828 =  ( n19099 ) ? ( VREG_22_12 ) : ( n19827 ) ;
assign n19829 =  ( n19098 ) ? ( VREG_22_13 ) : ( n19828 ) ;
assign n19830 =  ( n19097 ) ? ( VREG_22_14 ) : ( n19829 ) ;
assign n19831 =  ( n19096 ) ? ( VREG_22_15 ) : ( n19830 ) ;
assign n19832 =  ( n19095 ) ? ( VREG_23_0 ) : ( n19831 ) ;
assign n19833 =  ( n19094 ) ? ( VREG_23_1 ) : ( n19832 ) ;
assign n19834 =  ( n19093 ) ? ( VREG_23_2 ) : ( n19833 ) ;
assign n19835 =  ( n19092 ) ? ( VREG_23_3 ) : ( n19834 ) ;
assign n19836 =  ( n19091 ) ? ( VREG_23_4 ) : ( n19835 ) ;
assign n19837 =  ( n19090 ) ? ( VREG_23_5 ) : ( n19836 ) ;
assign n19838 =  ( n19089 ) ? ( VREG_23_6 ) : ( n19837 ) ;
assign n19839 =  ( n19088 ) ? ( VREG_23_7 ) : ( n19838 ) ;
assign n19840 =  ( n19087 ) ? ( VREG_23_8 ) : ( n19839 ) ;
assign n19841 =  ( n19086 ) ? ( VREG_23_9 ) : ( n19840 ) ;
assign n19842 =  ( n19085 ) ? ( VREG_23_10 ) : ( n19841 ) ;
assign n19843 =  ( n19084 ) ? ( VREG_23_11 ) : ( n19842 ) ;
assign n19844 =  ( n19083 ) ? ( VREG_23_12 ) : ( n19843 ) ;
assign n19845 =  ( n19082 ) ? ( VREG_23_13 ) : ( n19844 ) ;
assign n19846 =  ( n19081 ) ? ( VREG_23_14 ) : ( n19845 ) ;
assign n19847 =  ( n19080 ) ? ( VREG_23_15 ) : ( n19846 ) ;
assign n19848 =  ( n19079 ) ? ( VREG_24_0 ) : ( n19847 ) ;
assign n19849 =  ( n19078 ) ? ( VREG_24_1 ) : ( n19848 ) ;
assign n19850 =  ( n19077 ) ? ( VREG_24_2 ) : ( n19849 ) ;
assign n19851 =  ( n19076 ) ? ( VREG_24_3 ) : ( n19850 ) ;
assign n19852 =  ( n19075 ) ? ( VREG_24_4 ) : ( n19851 ) ;
assign n19853 =  ( n19074 ) ? ( VREG_24_5 ) : ( n19852 ) ;
assign n19854 =  ( n19073 ) ? ( VREG_24_6 ) : ( n19853 ) ;
assign n19855 =  ( n19072 ) ? ( VREG_24_7 ) : ( n19854 ) ;
assign n19856 =  ( n19071 ) ? ( VREG_24_8 ) : ( n19855 ) ;
assign n19857 =  ( n19070 ) ? ( VREG_24_9 ) : ( n19856 ) ;
assign n19858 =  ( n19069 ) ? ( VREG_24_10 ) : ( n19857 ) ;
assign n19859 =  ( n19068 ) ? ( VREG_24_11 ) : ( n19858 ) ;
assign n19860 =  ( n19067 ) ? ( VREG_24_12 ) : ( n19859 ) ;
assign n19861 =  ( n19066 ) ? ( VREG_24_13 ) : ( n19860 ) ;
assign n19862 =  ( n19065 ) ? ( VREG_24_14 ) : ( n19861 ) ;
assign n19863 =  ( n19064 ) ? ( VREG_24_15 ) : ( n19862 ) ;
assign n19864 =  ( n19063 ) ? ( VREG_25_0 ) : ( n19863 ) ;
assign n19865 =  ( n19062 ) ? ( VREG_25_1 ) : ( n19864 ) ;
assign n19866 =  ( n19061 ) ? ( VREG_25_2 ) : ( n19865 ) ;
assign n19867 =  ( n19060 ) ? ( VREG_25_3 ) : ( n19866 ) ;
assign n19868 =  ( n19059 ) ? ( VREG_25_4 ) : ( n19867 ) ;
assign n19869 =  ( n19058 ) ? ( VREG_25_5 ) : ( n19868 ) ;
assign n19870 =  ( n19057 ) ? ( VREG_25_6 ) : ( n19869 ) ;
assign n19871 =  ( n19056 ) ? ( VREG_25_7 ) : ( n19870 ) ;
assign n19872 =  ( n19055 ) ? ( VREG_25_8 ) : ( n19871 ) ;
assign n19873 =  ( n19054 ) ? ( VREG_25_9 ) : ( n19872 ) ;
assign n19874 =  ( n19053 ) ? ( VREG_25_10 ) : ( n19873 ) ;
assign n19875 =  ( n19052 ) ? ( VREG_25_11 ) : ( n19874 ) ;
assign n19876 =  ( n19051 ) ? ( VREG_25_12 ) : ( n19875 ) ;
assign n19877 =  ( n19050 ) ? ( VREG_25_13 ) : ( n19876 ) ;
assign n19878 =  ( n19049 ) ? ( VREG_25_14 ) : ( n19877 ) ;
assign n19879 =  ( n19048 ) ? ( VREG_25_15 ) : ( n19878 ) ;
assign n19880 =  ( n19047 ) ? ( VREG_26_0 ) : ( n19879 ) ;
assign n19881 =  ( n19046 ) ? ( VREG_26_1 ) : ( n19880 ) ;
assign n19882 =  ( n19045 ) ? ( VREG_26_2 ) : ( n19881 ) ;
assign n19883 =  ( n19044 ) ? ( VREG_26_3 ) : ( n19882 ) ;
assign n19884 =  ( n19043 ) ? ( VREG_26_4 ) : ( n19883 ) ;
assign n19885 =  ( n19042 ) ? ( VREG_26_5 ) : ( n19884 ) ;
assign n19886 =  ( n19041 ) ? ( VREG_26_6 ) : ( n19885 ) ;
assign n19887 =  ( n19040 ) ? ( VREG_26_7 ) : ( n19886 ) ;
assign n19888 =  ( n19039 ) ? ( VREG_26_8 ) : ( n19887 ) ;
assign n19889 =  ( n19038 ) ? ( VREG_26_9 ) : ( n19888 ) ;
assign n19890 =  ( n19037 ) ? ( VREG_26_10 ) : ( n19889 ) ;
assign n19891 =  ( n19036 ) ? ( VREG_26_11 ) : ( n19890 ) ;
assign n19892 =  ( n19035 ) ? ( VREG_26_12 ) : ( n19891 ) ;
assign n19893 =  ( n19034 ) ? ( VREG_26_13 ) : ( n19892 ) ;
assign n19894 =  ( n19033 ) ? ( VREG_26_14 ) : ( n19893 ) ;
assign n19895 =  ( n19032 ) ? ( VREG_26_15 ) : ( n19894 ) ;
assign n19896 =  ( n19031 ) ? ( VREG_27_0 ) : ( n19895 ) ;
assign n19897 =  ( n19030 ) ? ( VREG_27_1 ) : ( n19896 ) ;
assign n19898 =  ( n19029 ) ? ( VREG_27_2 ) : ( n19897 ) ;
assign n19899 =  ( n19028 ) ? ( VREG_27_3 ) : ( n19898 ) ;
assign n19900 =  ( n19027 ) ? ( VREG_27_4 ) : ( n19899 ) ;
assign n19901 =  ( n19026 ) ? ( VREG_27_5 ) : ( n19900 ) ;
assign n19902 =  ( n19025 ) ? ( VREG_27_6 ) : ( n19901 ) ;
assign n19903 =  ( n19024 ) ? ( VREG_27_7 ) : ( n19902 ) ;
assign n19904 =  ( n19023 ) ? ( VREG_27_8 ) : ( n19903 ) ;
assign n19905 =  ( n19022 ) ? ( VREG_27_9 ) : ( n19904 ) ;
assign n19906 =  ( n19021 ) ? ( VREG_27_10 ) : ( n19905 ) ;
assign n19907 =  ( n19020 ) ? ( VREG_27_11 ) : ( n19906 ) ;
assign n19908 =  ( n19019 ) ? ( VREG_27_12 ) : ( n19907 ) ;
assign n19909 =  ( n19018 ) ? ( VREG_27_13 ) : ( n19908 ) ;
assign n19910 =  ( n19017 ) ? ( VREG_27_14 ) : ( n19909 ) ;
assign n19911 =  ( n19016 ) ? ( VREG_27_15 ) : ( n19910 ) ;
assign n19912 =  ( n19015 ) ? ( VREG_28_0 ) : ( n19911 ) ;
assign n19913 =  ( n19014 ) ? ( VREG_28_1 ) : ( n19912 ) ;
assign n19914 =  ( n19013 ) ? ( VREG_28_2 ) : ( n19913 ) ;
assign n19915 =  ( n19012 ) ? ( VREG_28_3 ) : ( n19914 ) ;
assign n19916 =  ( n19011 ) ? ( VREG_28_4 ) : ( n19915 ) ;
assign n19917 =  ( n19010 ) ? ( VREG_28_5 ) : ( n19916 ) ;
assign n19918 =  ( n19009 ) ? ( VREG_28_6 ) : ( n19917 ) ;
assign n19919 =  ( n19008 ) ? ( VREG_28_7 ) : ( n19918 ) ;
assign n19920 =  ( n19007 ) ? ( VREG_28_8 ) : ( n19919 ) ;
assign n19921 =  ( n19006 ) ? ( VREG_28_9 ) : ( n19920 ) ;
assign n19922 =  ( n19005 ) ? ( VREG_28_10 ) : ( n19921 ) ;
assign n19923 =  ( n19004 ) ? ( VREG_28_11 ) : ( n19922 ) ;
assign n19924 =  ( n19003 ) ? ( VREG_28_12 ) : ( n19923 ) ;
assign n19925 =  ( n19002 ) ? ( VREG_28_13 ) : ( n19924 ) ;
assign n19926 =  ( n19001 ) ? ( VREG_28_14 ) : ( n19925 ) ;
assign n19927 =  ( n19000 ) ? ( VREG_28_15 ) : ( n19926 ) ;
assign n19928 =  ( n18999 ) ? ( VREG_29_0 ) : ( n19927 ) ;
assign n19929 =  ( n18998 ) ? ( VREG_29_1 ) : ( n19928 ) ;
assign n19930 =  ( n18997 ) ? ( VREG_29_2 ) : ( n19929 ) ;
assign n19931 =  ( n18996 ) ? ( VREG_29_3 ) : ( n19930 ) ;
assign n19932 =  ( n18995 ) ? ( VREG_29_4 ) : ( n19931 ) ;
assign n19933 =  ( n18994 ) ? ( VREG_29_5 ) : ( n19932 ) ;
assign n19934 =  ( n18993 ) ? ( VREG_29_6 ) : ( n19933 ) ;
assign n19935 =  ( n18992 ) ? ( VREG_29_7 ) : ( n19934 ) ;
assign n19936 =  ( n18991 ) ? ( VREG_29_8 ) : ( n19935 ) ;
assign n19937 =  ( n18990 ) ? ( VREG_29_9 ) : ( n19936 ) ;
assign n19938 =  ( n18989 ) ? ( VREG_29_10 ) : ( n19937 ) ;
assign n19939 =  ( n18988 ) ? ( VREG_29_11 ) : ( n19938 ) ;
assign n19940 =  ( n18987 ) ? ( VREG_29_12 ) : ( n19939 ) ;
assign n19941 =  ( n18986 ) ? ( VREG_29_13 ) : ( n19940 ) ;
assign n19942 =  ( n18985 ) ? ( VREG_29_14 ) : ( n19941 ) ;
assign n19943 =  ( n18984 ) ? ( VREG_29_15 ) : ( n19942 ) ;
assign n19944 =  ( n18983 ) ? ( VREG_30_0 ) : ( n19943 ) ;
assign n19945 =  ( n18982 ) ? ( VREG_30_1 ) : ( n19944 ) ;
assign n19946 =  ( n18981 ) ? ( VREG_30_2 ) : ( n19945 ) ;
assign n19947 =  ( n18980 ) ? ( VREG_30_3 ) : ( n19946 ) ;
assign n19948 =  ( n18979 ) ? ( VREG_30_4 ) : ( n19947 ) ;
assign n19949 =  ( n18978 ) ? ( VREG_30_5 ) : ( n19948 ) ;
assign n19950 =  ( n18977 ) ? ( VREG_30_6 ) : ( n19949 ) ;
assign n19951 =  ( n18976 ) ? ( VREG_30_7 ) : ( n19950 ) ;
assign n19952 =  ( n18975 ) ? ( VREG_30_8 ) : ( n19951 ) ;
assign n19953 =  ( n18974 ) ? ( VREG_30_9 ) : ( n19952 ) ;
assign n19954 =  ( n18973 ) ? ( VREG_30_10 ) : ( n19953 ) ;
assign n19955 =  ( n18972 ) ? ( VREG_30_11 ) : ( n19954 ) ;
assign n19956 =  ( n18971 ) ? ( VREG_30_12 ) : ( n19955 ) ;
assign n19957 =  ( n18970 ) ? ( VREG_30_13 ) : ( n19956 ) ;
assign n19958 =  ( n18969 ) ? ( VREG_30_14 ) : ( n19957 ) ;
assign n19959 =  ( n18968 ) ? ( VREG_30_15 ) : ( n19958 ) ;
assign n19960 =  ( n18967 ) ? ( VREG_31_0 ) : ( n19959 ) ;
assign n19961 =  ( n18966 ) ? ( VREG_31_1 ) : ( n19960 ) ;
assign n19962 =  ( n18965 ) ? ( VREG_31_2 ) : ( n19961 ) ;
assign n19963 =  ( n18964 ) ? ( VREG_31_3 ) : ( n19962 ) ;
assign n19964 =  ( n18963 ) ? ( VREG_31_4 ) : ( n19963 ) ;
assign n19965 =  ( n18962 ) ? ( VREG_31_5 ) : ( n19964 ) ;
assign n19966 =  ( n18961 ) ? ( VREG_31_6 ) : ( n19965 ) ;
assign n19967 =  ( n18960 ) ? ( VREG_31_7 ) : ( n19966 ) ;
assign n19968 =  ( n18959 ) ? ( VREG_31_8 ) : ( n19967 ) ;
assign n19969 =  ( n18958 ) ? ( VREG_31_9 ) : ( n19968 ) ;
assign n19970 =  ( n18957 ) ? ( VREG_31_10 ) : ( n19969 ) ;
assign n19971 =  ( n18956 ) ? ( VREG_31_11 ) : ( n19970 ) ;
assign n19972 =  ( n18955 ) ? ( VREG_31_12 ) : ( n19971 ) ;
assign n19973 =  ( n18954 ) ? ( VREG_31_13 ) : ( n19972 ) ;
assign n19974 =  ( n18953 ) ? ( VREG_31_14 ) : ( n19973 ) ;
assign n19975 =  ( n18952 ) ? ( VREG_31_15 ) : ( n19974 ) ;
assign n19976 =  ( n18941 ) + ( n19975 )  ;
assign n19977 =  ( n18941 ) - ( n19975 )  ;
assign n19978 =  ( n18941 ) & ( n19975 )  ;
assign n19979 =  ( n18941 ) | ( n19975 )  ;
assign n19980 =  ( ( n18941 ) * ( n19975 ))  ;
assign n19981 =  ( n148 ) ? ( n19980 ) : ( VREG_0_2 ) ;
assign n19982 =  ( n146 ) ? ( n19979 ) : ( n19981 ) ;
assign n19983 =  ( n144 ) ? ( n19978 ) : ( n19982 ) ;
assign n19984 =  ( n142 ) ? ( n19977 ) : ( n19983 ) ;
assign n19985 =  ( n10 ) ? ( n19976 ) : ( n19984 ) ;
assign n19986 = n3030[2:2] ;
assign n19987 =  ( n19986 ) == ( 1'd0 )  ;
assign n19988 =  ( n19987 ) ? ( VREG_0_2 ) : ( n18951 ) ;
assign n19989 =  ( n19987 ) ? ( VREG_0_2 ) : ( n19985 ) ;
assign n19990 =  ( n3034 ) ? ( n19989 ) : ( VREG_0_2 ) ;
assign n19991 =  ( n2965 ) ? ( n19988 ) : ( n19990 ) ;
assign n19992 =  ( n1930 ) ? ( n19985 ) : ( n19991 ) ;
assign n19993 =  ( n879 ) ? ( n18951 ) : ( n19992 ) ;
assign n19994 =  ( n18941 ) + ( n164 )  ;
assign n19995 =  ( n18941 ) - ( n164 )  ;
assign n19996 =  ( n18941 ) & ( n164 )  ;
assign n19997 =  ( n18941 ) | ( n164 )  ;
assign n19998 =  ( ( n18941 ) * ( n164 ))  ;
assign n19999 =  ( n172 ) ? ( n19998 ) : ( VREG_0_2 ) ;
assign n20000 =  ( n170 ) ? ( n19997 ) : ( n19999 ) ;
assign n20001 =  ( n168 ) ? ( n19996 ) : ( n20000 ) ;
assign n20002 =  ( n166 ) ? ( n19995 ) : ( n20001 ) ;
assign n20003 =  ( n162 ) ? ( n19994 ) : ( n20002 ) ;
assign n20004 =  ( n18941 ) + ( n180 )  ;
assign n20005 =  ( n18941 ) - ( n180 )  ;
assign n20006 =  ( n18941 ) & ( n180 )  ;
assign n20007 =  ( n18941 ) | ( n180 )  ;
assign n20008 =  ( ( n18941 ) * ( n180 ))  ;
assign n20009 =  ( n172 ) ? ( n20008 ) : ( VREG_0_2 ) ;
assign n20010 =  ( n170 ) ? ( n20007 ) : ( n20009 ) ;
assign n20011 =  ( n168 ) ? ( n20006 ) : ( n20010 ) ;
assign n20012 =  ( n166 ) ? ( n20005 ) : ( n20011 ) ;
assign n20013 =  ( n162 ) ? ( n20004 ) : ( n20012 ) ;
assign n20014 =  ( n19987 ) ? ( VREG_0_2 ) : ( n20013 ) ;
assign n20015 =  ( n3051 ) ? ( n20014 ) : ( VREG_0_2 ) ;
assign n20016 =  ( n3040 ) ? ( n20003 ) : ( n20015 ) ;
assign n20017 =  ( n192 ) ? ( VREG_0_2 ) : ( VREG_0_2 ) ;
assign n20018 =  ( n157 ) ? ( n20016 ) : ( n20017 ) ;
assign n20019 =  ( n6 ) ? ( n19993 ) : ( n20018 ) ;
assign n20020 =  ( n4 ) ? ( n20019 ) : ( VREG_0_2 ) ;
assign n20021 =  ( 32'd3 ) == ( 32'd15 )  ;
assign n20022 =  ( n12 ) & ( n20021 )  ;
assign n20023 =  ( 32'd3 ) == ( 32'd14 )  ;
assign n20024 =  ( n12 ) & ( n20023 )  ;
assign n20025 =  ( 32'd3 ) == ( 32'd13 )  ;
assign n20026 =  ( n12 ) & ( n20025 )  ;
assign n20027 =  ( 32'd3 ) == ( 32'd12 )  ;
assign n20028 =  ( n12 ) & ( n20027 )  ;
assign n20029 =  ( 32'd3 ) == ( 32'd11 )  ;
assign n20030 =  ( n12 ) & ( n20029 )  ;
assign n20031 =  ( 32'd3 ) == ( 32'd10 )  ;
assign n20032 =  ( n12 ) & ( n20031 )  ;
assign n20033 =  ( 32'd3 ) == ( 32'd9 )  ;
assign n20034 =  ( n12 ) & ( n20033 )  ;
assign n20035 =  ( 32'd3 ) == ( 32'd8 )  ;
assign n20036 =  ( n12 ) & ( n20035 )  ;
assign n20037 =  ( 32'd3 ) == ( 32'd7 )  ;
assign n20038 =  ( n12 ) & ( n20037 )  ;
assign n20039 =  ( 32'd3 ) == ( 32'd6 )  ;
assign n20040 =  ( n12 ) & ( n20039 )  ;
assign n20041 =  ( 32'd3 ) == ( 32'd5 )  ;
assign n20042 =  ( n12 ) & ( n20041 )  ;
assign n20043 =  ( 32'd3 ) == ( 32'd4 )  ;
assign n20044 =  ( n12 ) & ( n20043 )  ;
assign n20045 =  ( 32'd3 ) == ( 32'd3 )  ;
assign n20046 =  ( n12 ) & ( n20045 )  ;
assign n20047 =  ( 32'd3 ) == ( 32'd2 )  ;
assign n20048 =  ( n12 ) & ( n20047 )  ;
assign n20049 =  ( 32'd3 ) == ( 32'd1 )  ;
assign n20050 =  ( n12 ) & ( n20049 )  ;
assign n20051 =  ( 32'd3 ) == ( 32'd0 )  ;
assign n20052 =  ( n12 ) & ( n20051 )  ;
assign n20053 =  ( n13 ) & ( n20021 )  ;
assign n20054 =  ( n13 ) & ( n20023 )  ;
assign n20055 =  ( n13 ) & ( n20025 )  ;
assign n20056 =  ( n13 ) & ( n20027 )  ;
assign n20057 =  ( n13 ) & ( n20029 )  ;
assign n20058 =  ( n13 ) & ( n20031 )  ;
assign n20059 =  ( n13 ) & ( n20033 )  ;
assign n20060 =  ( n13 ) & ( n20035 )  ;
assign n20061 =  ( n13 ) & ( n20037 )  ;
assign n20062 =  ( n13 ) & ( n20039 )  ;
assign n20063 =  ( n13 ) & ( n20041 )  ;
assign n20064 =  ( n13 ) & ( n20043 )  ;
assign n20065 =  ( n13 ) & ( n20045 )  ;
assign n20066 =  ( n13 ) & ( n20047 )  ;
assign n20067 =  ( n13 ) & ( n20049 )  ;
assign n20068 =  ( n13 ) & ( n20051 )  ;
assign n20069 =  ( n14 ) & ( n20021 )  ;
assign n20070 =  ( n14 ) & ( n20023 )  ;
assign n20071 =  ( n14 ) & ( n20025 )  ;
assign n20072 =  ( n14 ) & ( n20027 )  ;
assign n20073 =  ( n14 ) & ( n20029 )  ;
assign n20074 =  ( n14 ) & ( n20031 )  ;
assign n20075 =  ( n14 ) & ( n20033 )  ;
assign n20076 =  ( n14 ) & ( n20035 )  ;
assign n20077 =  ( n14 ) & ( n20037 )  ;
assign n20078 =  ( n14 ) & ( n20039 )  ;
assign n20079 =  ( n14 ) & ( n20041 )  ;
assign n20080 =  ( n14 ) & ( n20043 )  ;
assign n20081 =  ( n14 ) & ( n20045 )  ;
assign n20082 =  ( n14 ) & ( n20047 )  ;
assign n20083 =  ( n14 ) & ( n20049 )  ;
assign n20084 =  ( n14 ) & ( n20051 )  ;
assign n20085 =  ( n15 ) & ( n20021 )  ;
assign n20086 =  ( n15 ) & ( n20023 )  ;
assign n20087 =  ( n15 ) & ( n20025 )  ;
assign n20088 =  ( n15 ) & ( n20027 )  ;
assign n20089 =  ( n15 ) & ( n20029 )  ;
assign n20090 =  ( n15 ) & ( n20031 )  ;
assign n20091 =  ( n15 ) & ( n20033 )  ;
assign n20092 =  ( n15 ) & ( n20035 )  ;
assign n20093 =  ( n15 ) & ( n20037 )  ;
assign n20094 =  ( n15 ) & ( n20039 )  ;
assign n20095 =  ( n15 ) & ( n20041 )  ;
assign n20096 =  ( n15 ) & ( n20043 )  ;
assign n20097 =  ( n15 ) & ( n20045 )  ;
assign n20098 =  ( n15 ) & ( n20047 )  ;
assign n20099 =  ( n15 ) & ( n20049 )  ;
assign n20100 =  ( n15 ) & ( n20051 )  ;
assign n20101 =  ( n16 ) & ( n20021 )  ;
assign n20102 =  ( n16 ) & ( n20023 )  ;
assign n20103 =  ( n16 ) & ( n20025 )  ;
assign n20104 =  ( n16 ) & ( n20027 )  ;
assign n20105 =  ( n16 ) & ( n20029 )  ;
assign n20106 =  ( n16 ) & ( n20031 )  ;
assign n20107 =  ( n16 ) & ( n20033 )  ;
assign n20108 =  ( n16 ) & ( n20035 )  ;
assign n20109 =  ( n16 ) & ( n20037 )  ;
assign n20110 =  ( n16 ) & ( n20039 )  ;
assign n20111 =  ( n16 ) & ( n20041 )  ;
assign n20112 =  ( n16 ) & ( n20043 )  ;
assign n20113 =  ( n16 ) & ( n20045 )  ;
assign n20114 =  ( n16 ) & ( n20047 )  ;
assign n20115 =  ( n16 ) & ( n20049 )  ;
assign n20116 =  ( n16 ) & ( n20051 )  ;
assign n20117 =  ( n17 ) & ( n20021 )  ;
assign n20118 =  ( n17 ) & ( n20023 )  ;
assign n20119 =  ( n17 ) & ( n20025 )  ;
assign n20120 =  ( n17 ) & ( n20027 )  ;
assign n20121 =  ( n17 ) & ( n20029 )  ;
assign n20122 =  ( n17 ) & ( n20031 )  ;
assign n20123 =  ( n17 ) & ( n20033 )  ;
assign n20124 =  ( n17 ) & ( n20035 )  ;
assign n20125 =  ( n17 ) & ( n20037 )  ;
assign n20126 =  ( n17 ) & ( n20039 )  ;
assign n20127 =  ( n17 ) & ( n20041 )  ;
assign n20128 =  ( n17 ) & ( n20043 )  ;
assign n20129 =  ( n17 ) & ( n20045 )  ;
assign n20130 =  ( n17 ) & ( n20047 )  ;
assign n20131 =  ( n17 ) & ( n20049 )  ;
assign n20132 =  ( n17 ) & ( n20051 )  ;
assign n20133 =  ( n18 ) & ( n20021 )  ;
assign n20134 =  ( n18 ) & ( n20023 )  ;
assign n20135 =  ( n18 ) & ( n20025 )  ;
assign n20136 =  ( n18 ) & ( n20027 )  ;
assign n20137 =  ( n18 ) & ( n20029 )  ;
assign n20138 =  ( n18 ) & ( n20031 )  ;
assign n20139 =  ( n18 ) & ( n20033 )  ;
assign n20140 =  ( n18 ) & ( n20035 )  ;
assign n20141 =  ( n18 ) & ( n20037 )  ;
assign n20142 =  ( n18 ) & ( n20039 )  ;
assign n20143 =  ( n18 ) & ( n20041 )  ;
assign n20144 =  ( n18 ) & ( n20043 )  ;
assign n20145 =  ( n18 ) & ( n20045 )  ;
assign n20146 =  ( n18 ) & ( n20047 )  ;
assign n20147 =  ( n18 ) & ( n20049 )  ;
assign n20148 =  ( n18 ) & ( n20051 )  ;
assign n20149 =  ( n19 ) & ( n20021 )  ;
assign n20150 =  ( n19 ) & ( n20023 )  ;
assign n20151 =  ( n19 ) & ( n20025 )  ;
assign n20152 =  ( n19 ) & ( n20027 )  ;
assign n20153 =  ( n19 ) & ( n20029 )  ;
assign n20154 =  ( n19 ) & ( n20031 )  ;
assign n20155 =  ( n19 ) & ( n20033 )  ;
assign n20156 =  ( n19 ) & ( n20035 )  ;
assign n20157 =  ( n19 ) & ( n20037 )  ;
assign n20158 =  ( n19 ) & ( n20039 )  ;
assign n20159 =  ( n19 ) & ( n20041 )  ;
assign n20160 =  ( n19 ) & ( n20043 )  ;
assign n20161 =  ( n19 ) & ( n20045 )  ;
assign n20162 =  ( n19 ) & ( n20047 )  ;
assign n20163 =  ( n19 ) & ( n20049 )  ;
assign n20164 =  ( n19 ) & ( n20051 )  ;
assign n20165 =  ( n20 ) & ( n20021 )  ;
assign n20166 =  ( n20 ) & ( n20023 )  ;
assign n20167 =  ( n20 ) & ( n20025 )  ;
assign n20168 =  ( n20 ) & ( n20027 )  ;
assign n20169 =  ( n20 ) & ( n20029 )  ;
assign n20170 =  ( n20 ) & ( n20031 )  ;
assign n20171 =  ( n20 ) & ( n20033 )  ;
assign n20172 =  ( n20 ) & ( n20035 )  ;
assign n20173 =  ( n20 ) & ( n20037 )  ;
assign n20174 =  ( n20 ) & ( n20039 )  ;
assign n20175 =  ( n20 ) & ( n20041 )  ;
assign n20176 =  ( n20 ) & ( n20043 )  ;
assign n20177 =  ( n20 ) & ( n20045 )  ;
assign n20178 =  ( n20 ) & ( n20047 )  ;
assign n20179 =  ( n20 ) & ( n20049 )  ;
assign n20180 =  ( n20 ) & ( n20051 )  ;
assign n20181 =  ( n21 ) & ( n20021 )  ;
assign n20182 =  ( n21 ) & ( n20023 )  ;
assign n20183 =  ( n21 ) & ( n20025 )  ;
assign n20184 =  ( n21 ) & ( n20027 )  ;
assign n20185 =  ( n21 ) & ( n20029 )  ;
assign n20186 =  ( n21 ) & ( n20031 )  ;
assign n20187 =  ( n21 ) & ( n20033 )  ;
assign n20188 =  ( n21 ) & ( n20035 )  ;
assign n20189 =  ( n21 ) & ( n20037 )  ;
assign n20190 =  ( n21 ) & ( n20039 )  ;
assign n20191 =  ( n21 ) & ( n20041 )  ;
assign n20192 =  ( n21 ) & ( n20043 )  ;
assign n20193 =  ( n21 ) & ( n20045 )  ;
assign n20194 =  ( n21 ) & ( n20047 )  ;
assign n20195 =  ( n21 ) & ( n20049 )  ;
assign n20196 =  ( n21 ) & ( n20051 )  ;
assign n20197 =  ( n22 ) & ( n20021 )  ;
assign n20198 =  ( n22 ) & ( n20023 )  ;
assign n20199 =  ( n22 ) & ( n20025 )  ;
assign n20200 =  ( n22 ) & ( n20027 )  ;
assign n20201 =  ( n22 ) & ( n20029 )  ;
assign n20202 =  ( n22 ) & ( n20031 )  ;
assign n20203 =  ( n22 ) & ( n20033 )  ;
assign n20204 =  ( n22 ) & ( n20035 )  ;
assign n20205 =  ( n22 ) & ( n20037 )  ;
assign n20206 =  ( n22 ) & ( n20039 )  ;
assign n20207 =  ( n22 ) & ( n20041 )  ;
assign n20208 =  ( n22 ) & ( n20043 )  ;
assign n20209 =  ( n22 ) & ( n20045 )  ;
assign n20210 =  ( n22 ) & ( n20047 )  ;
assign n20211 =  ( n22 ) & ( n20049 )  ;
assign n20212 =  ( n22 ) & ( n20051 )  ;
assign n20213 =  ( n23 ) & ( n20021 )  ;
assign n20214 =  ( n23 ) & ( n20023 )  ;
assign n20215 =  ( n23 ) & ( n20025 )  ;
assign n20216 =  ( n23 ) & ( n20027 )  ;
assign n20217 =  ( n23 ) & ( n20029 )  ;
assign n20218 =  ( n23 ) & ( n20031 )  ;
assign n20219 =  ( n23 ) & ( n20033 )  ;
assign n20220 =  ( n23 ) & ( n20035 )  ;
assign n20221 =  ( n23 ) & ( n20037 )  ;
assign n20222 =  ( n23 ) & ( n20039 )  ;
assign n20223 =  ( n23 ) & ( n20041 )  ;
assign n20224 =  ( n23 ) & ( n20043 )  ;
assign n20225 =  ( n23 ) & ( n20045 )  ;
assign n20226 =  ( n23 ) & ( n20047 )  ;
assign n20227 =  ( n23 ) & ( n20049 )  ;
assign n20228 =  ( n23 ) & ( n20051 )  ;
assign n20229 =  ( n24 ) & ( n20021 )  ;
assign n20230 =  ( n24 ) & ( n20023 )  ;
assign n20231 =  ( n24 ) & ( n20025 )  ;
assign n20232 =  ( n24 ) & ( n20027 )  ;
assign n20233 =  ( n24 ) & ( n20029 )  ;
assign n20234 =  ( n24 ) & ( n20031 )  ;
assign n20235 =  ( n24 ) & ( n20033 )  ;
assign n20236 =  ( n24 ) & ( n20035 )  ;
assign n20237 =  ( n24 ) & ( n20037 )  ;
assign n20238 =  ( n24 ) & ( n20039 )  ;
assign n20239 =  ( n24 ) & ( n20041 )  ;
assign n20240 =  ( n24 ) & ( n20043 )  ;
assign n20241 =  ( n24 ) & ( n20045 )  ;
assign n20242 =  ( n24 ) & ( n20047 )  ;
assign n20243 =  ( n24 ) & ( n20049 )  ;
assign n20244 =  ( n24 ) & ( n20051 )  ;
assign n20245 =  ( n25 ) & ( n20021 )  ;
assign n20246 =  ( n25 ) & ( n20023 )  ;
assign n20247 =  ( n25 ) & ( n20025 )  ;
assign n20248 =  ( n25 ) & ( n20027 )  ;
assign n20249 =  ( n25 ) & ( n20029 )  ;
assign n20250 =  ( n25 ) & ( n20031 )  ;
assign n20251 =  ( n25 ) & ( n20033 )  ;
assign n20252 =  ( n25 ) & ( n20035 )  ;
assign n20253 =  ( n25 ) & ( n20037 )  ;
assign n20254 =  ( n25 ) & ( n20039 )  ;
assign n20255 =  ( n25 ) & ( n20041 )  ;
assign n20256 =  ( n25 ) & ( n20043 )  ;
assign n20257 =  ( n25 ) & ( n20045 )  ;
assign n20258 =  ( n25 ) & ( n20047 )  ;
assign n20259 =  ( n25 ) & ( n20049 )  ;
assign n20260 =  ( n25 ) & ( n20051 )  ;
assign n20261 =  ( n26 ) & ( n20021 )  ;
assign n20262 =  ( n26 ) & ( n20023 )  ;
assign n20263 =  ( n26 ) & ( n20025 )  ;
assign n20264 =  ( n26 ) & ( n20027 )  ;
assign n20265 =  ( n26 ) & ( n20029 )  ;
assign n20266 =  ( n26 ) & ( n20031 )  ;
assign n20267 =  ( n26 ) & ( n20033 )  ;
assign n20268 =  ( n26 ) & ( n20035 )  ;
assign n20269 =  ( n26 ) & ( n20037 )  ;
assign n20270 =  ( n26 ) & ( n20039 )  ;
assign n20271 =  ( n26 ) & ( n20041 )  ;
assign n20272 =  ( n26 ) & ( n20043 )  ;
assign n20273 =  ( n26 ) & ( n20045 )  ;
assign n20274 =  ( n26 ) & ( n20047 )  ;
assign n20275 =  ( n26 ) & ( n20049 )  ;
assign n20276 =  ( n26 ) & ( n20051 )  ;
assign n20277 =  ( n27 ) & ( n20021 )  ;
assign n20278 =  ( n27 ) & ( n20023 )  ;
assign n20279 =  ( n27 ) & ( n20025 )  ;
assign n20280 =  ( n27 ) & ( n20027 )  ;
assign n20281 =  ( n27 ) & ( n20029 )  ;
assign n20282 =  ( n27 ) & ( n20031 )  ;
assign n20283 =  ( n27 ) & ( n20033 )  ;
assign n20284 =  ( n27 ) & ( n20035 )  ;
assign n20285 =  ( n27 ) & ( n20037 )  ;
assign n20286 =  ( n27 ) & ( n20039 )  ;
assign n20287 =  ( n27 ) & ( n20041 )  ;
assign n20288 =  ( n27 ) & ( n20043 )  ;
assign n20289 =  ( n27 ) & ( n20045 )  ;
assign n20290 =  ( n27 ) & ( n20047 )  ;
assign n20291 =  ( n27 ) & ( n20049 )  ;
assign n20292 =  ( n27 ) & ( n20051 )  ;
assign n20293 =  ( n28 ) & ( n20021 )  ;
assign n20294 =  ( n28 ) & ( n20023 )  ;
assign n20295 =  ( n28 ) & ( n20025 )  ;
assign n20296 =  ( n28 ) & ( n20027 )  ;
assign n20297 =  ( n28 ) & ( n20029 )  ;
assign n20298 =  ( n28 ) & ( n20031 )  ;
assign n20299 =  ( n28 ) & ( n20033 )  ;
assign n20300 =  ( n28 ) & ( n20035 )  ;
assign n20301 =  ( n28 ) & ( n20037 )  ;
assign n20302 =  ( n28 ) & ( n20039 )  ;
assign n20303 =  ( n28 ) & ( n20041 )  ;
assign n20304 =  ( n28 ) & ( n20043 )  ;
assign n20305 =  ( n28 ) & ( n20045 )  ;
assign n20306 =  ( n28 ) & ( n20047 )  ;
assign n20307 =  ( n28 ) & ( n20049 )  ;
assign n20308 =  ( n28 ) & ( n20051 )  ;
assign n20309 =  ( n29 ) & ( n20021 )  ;
assign n20310 =  ( n29 ) & ( n20023 )  ;
assign n20311 =  ( n29 ) & ( n20025 )  ;
assign n20312 =  ( n29 ) & ( n20027 )  ;
assign n20313 =  ( n29 ) & ( n20029 )  ;
assign n20314 =  ( n29 ) & ( n20031 )  ;
assign n20315 =  ( n29 ) & ( n20033 )  ;
assign n20316 =  ( n29 ) & ( n20035 )  ;
assign n20317 =  ( n29 ) & ( n20037 )  ;
assign n20318 =  ( n29 ) & ( n20039 )  ;
assign n20319 =  ( n29 ) & ( n20041 )  ;
assign n20320 =  ( n29 ) & ( n20043 )  ;
assign n20321 =  ( n29 ) & ( n20045 )  ;
assign n20322 =  ( n29 ) & ( n20047 )  ;
assign n20323 =  ( n29 ) & ( n20049 )  ;
assign n20324 =  ( n29 ) & ( n20051 )  ;
assign n20325 =  ( n30 ) & ( n20021 )  ;
assign n20326 =  ( n30 ) & ( n20023 )  ;
assign n20327 =  ( n30 ) & ( n20025 )  ;
assign n20328 =  ( n30 ) & ( n20027 )  ;
assign n20329 =  ( n30 ) & ( n20029 )  ;
assign n20330 =  ( n30 ) & ( n20031 )  ;
assign n20331 =  ( n30 ) & ( n20033 )  ;
assign n20332 =  ( n30 ) & ( n20035 )  ;
assign n20333 =  ( n30 ) & ( n20037 )  ;
assign n20334 =  ( n30 ) & ( n20039 )  ;
assign n20335 =  ( n30 ) & ( n20041 )  ;
assign n20336 =  ( n30 ) & ( n20043 )  ;
assign n20337 =  ( n30 ) & ( n20045 )  ;
assign n20338 =  ( n30 ) & ( n20047 )  ;
assign n20339 =  ( n30 ) & ( n20049 )  ;
assign n20340 =  ( n30 ) & ( n20051 )  ;
assign n20341 =  ( n31 ) & ( n20021 )  ;
assign n20342 =  ( n31 ) & ( n20023 )  ;
assign n20343 =  ( n31 ) & ( n20025 )  ;
assign n20344 =  ( n31 ) & ( n20027 )  ;
assign n20345 =  ( n31 ) & ( n20029 )  ;
assign n20346 =  ( n31 ) & ( n20031 )  ;
assign n20347 =  ( n31 ) & ( n20033 )  ;
assign n20348 =  ( n31 ) & ( n20035 )  ;
assign n20349 =  ( n31 ) & ( n20037 )  ;
assign n20350 =  ( n31 ) & ( n20039 )  ;
assign n20351 =  ( n31 ) & ( n20041 )  ;
assign n20352 =  ( n31 ) & ( n20043 )  ;
assign n20353 =  ( n31 ) & ( n20045 )  ;
assign n20354 =  ( n31 ) & ( n20047 )  ;
assign n20355 =  ( n31 ) & ( n20049 )  ;
assign n20356 =  ( n31 ) & ( n20051 )  ;
assign n20357 =  ( n32 ) & ( n20021 )  ;
assign n20358 =  ( n32 ) & ( n20023 )  ;
assign n20359 =  ( n32 ) & ( n20025 )  ;
assign n20360 =  ( n32 ) & ( n20027 )  ;
assign n20361 =  ( n32 ) & ( n20029 )  ;
assign n20362 =  ( n32 ) & ( n20031 )  ;
assign n20363 =  ( n32 ) & ( n20033 )  ;
assign n20364 =  ( n32 ) & ( n20035 )  ;
assign n20365 =  ( n32 ) & ( n20037 )  ;
assign n20366 =  ( n32 ) & ( n20039 )  ;
assign n20367 =  ( n32 ) & ( n20041 )  ;
assign n20368 =  ( n32 ) & ( n20043 )  ;
assign n20369 =  ( n32 ) & ( n20045 )  ;
assign n20370 =  ( n32 ) & ( n20047 )  ;
assign n20371 =  ( n32 ) & ( n20049 )  ;
assign n20372 =  ( n32 ) & ( n20051 )  ;
assign n20373 =  ( n33 ) & ( n20021 )  ;
assign n20374 =  ( n33 ) & ( n20023 )  ;
assign n20375 =  ( n33 ) & ( n20025 )  ;
assign n20376 =  ( n33 ) & ( n20027 )  ;
assign n20377 =  ( n33 ) & ( n20029 )  ;
assign n20378 =  ( n33 ) & ( n20031 )  ;
assign n20379 =  ( n33 ) & ( n20033 )  ;
assign n20380 =  ( n33 ) & ( n20035 )  ;
assign n20381 =  ( n33 ) & ( n20037 )  ;
assign n20382 =  ( n33 ) & ( n20039 )  ;
assign n20383 =  ( n33 ) & ( n20041 )  ;
assign n20384 =  ( n33 ) & ( n20043 )  ;
assign n20385 =  ( n33 ) & ( n20045 )  ;
assign n20386 =  ( n33 ) & ( n20047 )  ;
assign n20387 =  ( n33 ) & ( n20049 )  ;
assign n20388 =  ( n33 ) & ( n20051 )  ;
assign n20389 =  ( n34 ) & ( n20021 )  ;
assign n20390 =  ( n34 ) & ( n20023 )  ;
assign n20391 =  ( n34 ) & ( n20025 )  ;
assign n20392 =  ( n34 ) & ( n20027 )  ;
assign n20393 =  ( n34 ) & ( n20029 )  ;
assign n20394 =  ( n34 ) & ( n20031 )  ;
assign n20395 =  ( n34 ) & ( n20033 )  ;
assign n20396 =  ( n34 ) & ( n20035 )  ;
assign n20397 =  ( n34 ) & ( n20037 )  ;
assign n20398 =  ( n34 ) & ( n20039 )  ;
assign n20399 =  ( n34 ) & ( n20041 )  ;
assign n20400 =  ( n34 ) & ( n20043 )  ;
assign n20401 =  ( n34 ) & ( n20045 )  ;
assign n20402 =  ( n34 ) & ( n20047 )  ;
assign n20403 =  ( n34 ) & ( n20049 )  ;
assign n20404 =  ( n34 ) & ( n20051 )  ;
assign n20405 =  ( n35 ) & ( n20021 )  ;
assign n20406 =  ( n35 ) & ( n20023 )  ;
assign n20407 =  ( n35 ) & ( n20025 )  ;
assign n20408 =  ( n35 ) & ( n20027 )  ;
assign n20409 =  ( n35 ) & ( n20029 )  ;
assign n20410 =  ( n35 ) & ( n20031 )  ;
assign n20411 =  ( n35 ) & ( n20033 )  ;
assign n20412 =  ( n35 ) & ( n20035 )  ;
assign n20413 =  ( n35 ) & ( n20037 )  ;
assign n20414 =  ( n35 ) & ( n20039 )  ;
assign n20415 =  ( n35 ) & ( n20041 )  ;
assign n20416 =  ( n35 ) & ( n20043 )  ;
assign n20417 =  ( n35 ) & ( n20045 )  ;
assign n20418 =  ( n35 ) & ( n20047 )  ;
assign n20419 =  ( n35 ) & ( n20049 )  ;
assign n20420 =  ( n35 ) & ( n20051 )  ;
assign n20421 =  ( n36 ) & ( n20021 )  ;
assign n20422 =  ( n36 ) & ( n20023 )  ;
assign n20423 =  ( n36 ) & ( n20025 )  ;
assign n20424 =  ( n36 ) & ( n20027 )  ;
assign n20425 =  ( n36 ) & ( n20029 )  ;
assign n20426 =  ( n36 ) & ( n20031 )  ;
assign n20427 =  ( n36 ) & ( n20033 )  ;
assign n20428 =  ( n36 ) & ( n20035 )  ;
assign n20429 =  ( n36 ) & ( n20037 )  ;
assign n20430 =  ( n36 ) & ( n20039 )  ;
assign n20431 =  ( n36 ) & ( n20041 )  ;
assign n20432 =  ( n36 ) & ( n20043 )  ;
assign n20433 =  ( n36 ) & ( n20045 )  ;
assign n20434 =  ( n36 ) & ( n20047 )  ;
assign n20435 =  ( n36 ) & ( n20049 )  ;
assign n20436 =  ( n36 ) & ( n20051 )  ;
assign n20437 =  ( n37 ) & ( n20021 )  ;
assign n20438 =  ( n37 ) & ( n20023 )  ;
assign n20439 =  ( n37 ) & ( n20025 )  ;
assign n20440 =  ( n37 ) & ( n20027 )  ;
assign n20441 =  ( n37 ) & ( n20029 )  ;
assign n20442 =  ( n37 ) & ( n20031 )  ;
assign n20443 =  ( n37 ) & ( n20033 )  ;
assign n20444 =  ( n37 ) & ( n20035 )  ;
assign n20445 =  ( n37 ) & ( n20037 )  ;
assign n20446 =  ( n37 ) & ( n20039 )  ;
assign n20447 =  ( n37 ) & ( n20041 )  ;
assign n20448 =  ( n37 ) & ( n20043 )  ;
assign n20449 =  ( n37 ) & ( n20045 )  ;
assign n20450 =  ( n37 ) & ( n20047 )  ;
assign n20451 =  ( n37 ) & ( n20049 )  ;
assign n20452 =  ( n37 ) & ( n20051 )  ;
assign n20453 =  ( n38 ) & ( n20021 )  ;
assign n20454 =  ( n38 ) & ( n20023 )  ;
assign n20455 =  ( n38 ) & ( n20025 )  ;
assign n20456 =  ( n38 ) & ( n20027 )  ;
assign n20457 =  ( n38 ) & ( n20029 )  ;
assign n20458 =  ( n38 ) & ( n20031 )  ;
assign n20459 =  ( n38 ) & ( n20033 )  ;
assign n20460 =  ( n38 ) & ( n20035 )  ;
assign n20461 =  ( n38 ) & ( n20037 )  ;
assign n20462 =  ( n38 ) & ( n20039 )  ;
assign n20463 =  ( n38 ) & ( n20041 )  ;
assign n20464 =  ( n38 ) & ( n20043 )  ;
assign n20465 =  ( n38 ) & ( n20045 )  ;
assign n20466 =  ( n38 ) & ( n20047 )  ;
assign n20467 =  ( n38 ) & ( n20049 )  ;
assign n20468 =  ( n38 ) & ( n20051 )  ;
assign n20469 =  ( n39 ) & ( n20021 )  ;
assign n20470 =  ( n39 ) & ( n20023 )  ;
assign n20471 =  ( n39 ) & ( n20025 )  ;
assign n20472 =  ( n39 ) & ( n20027 )  ;
assign n20473 =  ( n39 ) & ( n20029 )  ;
assign n20474 =  ( n39 ) & ( n20031 )  ;
assign n20475 =  ( n39 ) & ( n20033 )  ;
assign n20476 =  ( n39 ) & ( n20035 )  ;
assign n20477 =  ( n39 ) & ( n20037 )  ;
assign n20478 =  ( n39 ) & ( n20039 )  ;
assign n20479 =  ( n39 ) & ( n20041 )  ;
assign n20480 =  ( n39 ) & ( n20043 )  ;
assign n20481 =  ( n39 ) & ( n20045 )  ;
assign n20482 =  ( n39 ) & ( n20047 )  ;
assign n20483 =  ( n39 ) & ( n20049 )  ;
assign n20484 =  ( n39 ) & ( n20051 )  ;
assign n20485 =  ( n40 ) & ( n20021 )  ;
assign n20486 =  ( n40 ) & ( n20023 )  ;
assign n20487 =  ( n40 ) & ( n20025 )  ;
assign n20488 =  ( n40 ) & ( n20027 )  ;
assign n20489 =  ( n40 ) & ( n20029 )  ;
assign n20490 =  ( n40 ) & ( n20031 )  ;
assign n20491 =  ( n40 ) & ( n20033 )  ;
assign n20492 =  ( n40 ) & ( n20035 )  ;
assign n20493 =  ( n40 ) & ( n20037 )  ;
assign n20494 =  ( n40 ) & ( n20039 )  ;
assign n20495 =  ( n40 ) & ( n20041 )  ;
assign n20496 =  ( n40 ) & ( n20043 )  ;
assign n20497 =  ( n40 ) & ( n20045 )  ;
assign n20498 =  ( n40 ) & ( n20047 )  ;
assign n20499 =  ( n40 ) & ( n20049 )  ;
assign n20500 =  ( n40 ) & ( n20051 )  ;
assign n20501 =  ( n41 ) & ( n20021 )  ;
assign n20502 =  ( n41 ) & ( n20023 )  ;
assign n20503 =  ( n41 ) & ( n20025 )  ;
assign n20504 =  ( n41 ) & ( n20027 )  ;
assign n20505 =  ( n41 ) & ( n20029 )  ;
assign n20506 =  ( n41 ) & ( n20031 )  ;
assign n20507 =  ( n41 ) & ( n20033 )  ;
assign n20508 =  ( n41 ) & ( n20035 )  ;
assign n20509 =  ( n41 ) & ( n20037 )  ;
assign n20510 =  ( n41 ) & ( n20039 )  ;
assign n20511 =  ( n41 ) & ( n20041 )  ;
assign n20512 =  ( n41 ) & ( n20043 )  ;
assign n20513 =  ( n41 ) & ( n20045 )  ;
assign n20514 =  ( n41 ) & ( n20047 )  ;
assign n20515 =  ( n41 ) & ( n20049 )  ;
assign n20516 =  ( n41 ) & ( n20051 )  ;
assign n20517 =  ( n42 ) & ( n20021 )  ;
assign n20518 =  ( n42 ) & ( n20023 )  ;
assign n20519 =  ( n42 ) & ( n20025 )  ;
assign n20520 =  ( n42 ) & ( n20027 )  ;
assign n20521 =  ( n42 ) & ( n20029 )  ;
assign n20522 =  ( n42 ) & ( n20031 )  ;
assign n20523 =  ( n42 ) & ( n20033 )  ;
assign n20524 =  ( n42 ) & ( n20035 )  ;
assign n20525 =  ( n42 ) & ( n20037 )  ;
assign n20526 =  ( n42 ) & ( n20039 )  ;
assign n20527 =  ( n42 ) & ( n20041 )  ;
assign n20528 =  ( n42 ) & ( n20043 )  ;
assign n20529 =  ( n42 ) & ( n20045 )  ;
assign n20530 =  ( n42 ) & ( n20047 )  ;
assign n20531 =  ( n42 ) & ( n20049 )  ;
assign n20532 =  ( n42 ) & ( n20051 )  ;
assign n20533 =  ( n43 ) & ( n20021 )  ;
assign n20534 =  ( n43 ) & ( n20023 )  ;
assign n20535 =  ( n43 ) & ( n20025 )  ;
assign n20536 =  ( n43 ) & ( n20027 )  ;
assign n20537 =  ( n43 ) & ( n20029 )  ;
assign n20538 =  ( n43 ) & ( n20031 )  ;
assign n20539 =  ( n43 ) & ( n20033 )  ;
assign n20540 =  ( n43 ) & ( n20035 )  ;
assign n20541 =  ( n43 ) & ( n20037 )  ;
assign n20542 =  ( n43 ) & ( n20039 )  ;
assign n20543 =  ( n43 ) & ( n20041 )  ;
assign n20544 =  ( n43 ) & ( n20043 )  ;
assign n20545 =  ( n43 ) & ( n20045 )  ;
assign n20546 =  ( n43 ) & ( n20047 )  ;
assign n20547 =  ( n43 ) & ( n20049 )  ;
assign n20548 =  ( n43 ) & ( n20051 )  ;
assign n20549 =  ( n20548 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n20550 =  ( n20547 ) ? ( VREG_0_1 ) : ( n20549 ) ;
assign n20551 =  ( n20546 ) ? ( VREG_0_2 ) : ( n20550 ) ;
assign n20552 =  ( n20545 ) ? ( VREG_0_3 ) : ( n20551 ) ;
assign n20553 =  ( n20544 ) ? ( VREG_0_4 ) : ( n20552 ) ;
assign n20554 =  ( n20543 ) ? ( VREG_0_5 ) : ( n20553 ) ;
assign n20555 =  ( n20542 ) ? ( VREG_0_6 ) : ( n20554 ) ;
assign n20556 =  ( n20541 ) ? ( VREG_0_7 ) : ( n20555 ) ;
assign n20557 =  ( n20540 ) ? ( VREG_0_8 ) : ( n20556 ) ;
assign n20558 =  ( n20539 ) ? ( VREG_0_9 ) : ( n20557 ) ;
assign n20559 =  ( n20538 ) ? ( VREG_0_10 ) : ( n20558 ) ;
assign n20560 =  ( n20537 ) ? ( VREG_0_11 ) : ( n20559 ) ;
assign n20561 =  ( n20536 ) ? ( VREG_0_12 ) : ( n20560 ) ;
assign n20562 =  ( n20535 ) ? ( VREG_0_13 ) : ( n20561 ) ;
assign n20563 =  ( n20534 ) ? ( VREG_0_14 ) : ( n20562 ) ;
assign n20564 =  ( n20533 ) ? ( VREG_0_15 ) : ( n20563 ) ;
assign n20565 =  ( n20532 ) ? ( VREG_1_0 ) : ( n20564 ) ;
assign n20566 =  ( n20531 ) ? ( VREG_1_1 ) : ( n20565 ) ;
assign n20567 =  ( n20530 ) ? ( VREG_1_2 ) : ( n20566 ) ;
assign n20568 =  ( n20529 ) ? ( VREG_1_3 ) : ( n20567 ) ;
assign n20569 =  ( n20528 ) ? ( VREG_1_4 ) : ( n20568 ) ;
assign n20570 =  ( n20527 ) ? ( VREG_1_5 ) : ( n20569 ) ;
assign n20571 =  ( n20526 ) ? ( VREG_1_6 ) : ( n20570 ) ;
assign n20572 =  ( n20525 ) ? ( VREG_1_7 ) : ( n20571 ) ;
assign n20573 =  ( n20524 ) ? ( VREG_1_8 ) : ( n20572 ) ;
assign n20574 =  ( n20523 ) ? ( VREG_1_9 ) : ( n20573 ) ;
assign n20575 =  ( n20522 ) ? ( VREG_1_10 ) : ( n20574 ) ;
assign n20576 =  ( n20521 ) ? ( VREG_1_11 ) : ( n20575 ) ;
assign n20577 =  ( n20520 ) ? ( VREG_1_12 ) : ( n20576 ) ;
assign n20578 =  ( n20519 ) ? ( VREG_1_13 ) : ( n20577 ) ;
assign n20579 =  ( n20518 ) ? ( VREG_1_14 ) : ( n20578 ) ;
assign n20580 =  ( n20517 ) ? ( VREG_1_15 ) : ( n20579 ) ;
assign n20581 =  ( n20516 ) ? ( VREG_2_0 ) : ( n20580 ) ;
assign n20582 =  ( n20515 ) ? ( VREG_2_1 ) : ( n20581 ) ;
assign n20583 =  ( n20514 ) ? ( VREG_2_2 ) : ( n20582 ) ;
assign n20584 =  ( n20513 ) ? ( VREG_2_3 ) : ( n20583 ) ;
assign n20585 =  ( n20512 ) ? ( VREG_2_4 ) : ( n20584 ) ;
assign n20586 =  ( n20511 ) ? ( VREG_2_5 ) : ( n20585 ) ;
assign n20587 =  ( n20510 ) ? ( VREG_2_6 ) : ( n20586 ) ;
assign n20588 =  ( n20509 ) ? ( VREG_2_7 ) : ( n20587 ) ;
assign n20589 =  ( n20508 ) ? ( VREG_2_8 ) : ( n20588 ) ;
assign n20590 =  ( n20507 ) ? ( VREG_2_9 ) : ( n20589 ) ;
assign n20591 =  ( n20506 ) ? ( VREG_2_10 ) : ( n20590 ) ;
assign n20592 =  ( n20505 ) ? ( VREG_2_11 ) : ( n20591 ) ;
assign n20593 =  ( n20504 ) ? ( VREG_2_12 ) : ( n20592 ) ;
assign n20594 =  ( n20503 ) ? ( VREG_2_13 ) : ( n20593 ) ;
assign n20595 =  ( n20502 ) ? ( VREG_2_14 ) : ( n20594 ) ;
assign n20596 =  ( n20501 ) ? ( VREG_2_15 ) : ( n20595 ) ;
assign n20597 =  ( n20500 ) ? ( VREG_3_0 ) : ( n20596 ) ;
assign n20598 =  ( n20499 ) ? ( VREG_3_1 ) : ( n20597 ) ;
assign n20599 =  ( n20498 ) ? ( VREG_3_2 ) : ( n20598 ) ;
assign n20600 =  ( n20497 ) ? ( VREG_3_3 ) : ( n20599 ) ;
assign n20601 =  ( n20496 ) ? ( VREG_3_4 ) : ( n20600 ) ;
assign n20602 =  ( n20495 ) ? ( VREG_3_5 ) : ( n20601 ) ;
assign n20603 =  ( n20494 ) ? ( VREG_3_6 ) : ( n20602 ) ;
assign n20604 =  ( n20493 ) ? ( VREG_3_7 ) : ( n20603 ) ;
assign n20605 =  ( n20492 ) ? ( VREG_3_8 ) : ( n20604 ) ;
assign n20606 =  ( n20491 ) ? ( VREG_3_9 ) : ( n20605 ) ;
assign n20607 =  ( n20490 ) ? ( VREG_3_10 ) : ( n20606 ) ;
assign n20608 =  ( n20489 ) ? ( VREG_3_11 ) : ( n20607 ) ;
assign n20609 =  ( n20488 ) ? ( VREG_3_12 ) : ( n20608 ) ;
assign n20610 =  ( n20487 ) ? ( VREG_3_13 ) : ( n20609 ) ;
assign n20611 =  ( n20486 ) ? ( VREG_3_14 ) : ( n20610 ) ;
assign n20612 =  ( n20485 ) ? ( VREG_3_15 ) : ( n20611 ) ;
assign n20613 =  ( n20484 ) ? ( VREG_4_0 ) : ( n20612 ) ;
assign n20614 =  ( n20483 ) ? ( VREG_4_1 ) : ( n20613 ) ;
assign n20615 =  ( n20482 ) ? ( VREG_4_2 ) : ( n20614 ) ;
assign n20616 =  ( n20481 ) ? ( VREG_4_3 ) : ( n20615 ) ;
assign n20617 =  ( n20480 ) ? ( VREG_4_4 ) : ( n20616 ) ;
assign n20618 =  ( n20479 ) ? ( VREG_4_5 ) : ( n20617 ) ;
assign n20619 =  ( n20478 ) ? ( VREG_4_6 ) : ( n20618 ) ;
assign n20620 =  ( n20477 ) ? ( VREG_4_7 ) : ( n20619 ) ;
assign n20621 =  ( n20476 ) ? ( VREG_4_8 ) : ( n20620 ) ;
assign n20622 =  ( n20475 ) ? ( VREG_4_9 ) : ( n20621 ) ;
assign n20623 =  ( n20474 ) ? ( VREG_4_10 ) : ( n20622 ) ;
assign n20624 =  ( n20473 ) ? ( VREG_4_11 ) : ( n20623 ) ;
assign n20625 =  ( n20472 ) ? ( VREG_4_12 ) : ( n20624 ) ;
assign n20626 =  ( n20471 ) ? ( VREG_4_13 ) : ( n20625 ) ;
assign n20627 =  ( n20470 ) ? ( VREG_4_14 ) : ( n20626 ) ;
assign n20628 =  ( n20469 ) ? ( VREG_4_15 ) : ( n20627 ) ;
assign n20629 =  ( n20468 ) ? ( VREG_5_0 ) : ( n20628 ) ;
assign n20630 =  ( n20467 ) ? ( VREG_5_1 ) : ( n20629 ) ;
assign n20631 =  ( n20466 ) ? ( VREG_5_2 ) : ( n20630 ) ;
assign n20632 =  ( n20465 ) ? ( VREG_5_3 ) : ( n20631 ) ;
assign n20633 =  ( n20464 ) ? ( VREG_5_4 ) : ( n20632 ) ;
assign n20634 =  ( n20463 ) ? ( VREG_5_5 ) : ( n20633 ) ;
assign n20635 =  ( n20462 ) ? ( VREG_5_6 ) : ( n20634 ) ;
assign n20636 =  ( n20461 ) ? ( VREG_5_7 ) : ( n20635 ) ;
assign n20637 =  ( n20460 ) ? ( VREG_5_8 ) : ( n20636 ) ;
assign n20638 =  ( n20459 ) ? ( VREG_5_9 ) : ( n20637 ) ;
assign n20639 =  ( n20458 ) ? ( VREG_5_10 ) : ( n20638 ) ;
assign n20640 =  ( n20457 ) ? ( VREG_5_11 ) : ( n20639 ) ;
assign n20641 =  ( n20456 ) ? ( VREG_5_12 ) : ( n20640 ) ;
assign n20642 =  ( n20455 ) ? ( VREG_5_13 ) : ( n20641 ) ;
assign n20643 =  ( n20454 ) ? ( VREG_5_14 ) : ( n20642 ) ;
assign n20644 =  ( n20453 ) ? ( VREG_5_15 ) : ( n20643 ) ;
assign n20645 =  ( n20452 ) ? ( VREG_6_0 ) : ( n20644 ) ;
assign n20646 =  ( n20451 ) ? ( VREG_6_1 ) : ( n20645 ) ;
assign n20647 =  ( n20450 ) ? ( VREG_6_2 ) : ( n20646 ) ;
assign n20648 =  ( n20449 ) ? ( VREG_6_3 ) : ( n20647 ) ;
assign n20649 =  ( n20448 ) ? ( VREG_6_4 ) : ( n20648 ) ;
assign n20650 =  ( n20447 ) ? ( VREG_6_5 ) : ( n20649 ) ;
assign n20651 =  ( n20446 ) ? ( VREG_6_6 ) : ( n20650 ) ;
assign n20652 =  ( n20445 ) ? ( VREG_6_7 ) : ( n20651 ) ;
assign n20653 =  ( n20444 ) ? ( VREG_6_8 ) : ( n20652 ) ;
assign n20654 =  ( n20443 ) ? ( VREG_6_9 ) : ( n20653 ) ;
assign n20655 =  ( n20442 ) ? ( VREG_6_10 ) : ( n20654 ) ;
assign n20656 =  ( n20441 ) ? ( VREG_6_11 ) : ( n20655 ) ;
assign n20657 =  ( n20440 ) ? ( VREG_6_12 ) : ( n20656 ) ;
assign n20658 =  ( n20439 ) ? ( VREG_6_13 ) : ( n20657 ) ;
assign n20659 =  ( n20438 ) ? ( VREG_6_14 ) : ( n20658 ) ;
assign n20660 =  ( n20437 ) ? ( VREG_6_15 ) : ( n20659 ) ;
assign n20661 =  ( n20436 ) ? ( VREG_7_0 ) : ( n20660 ) ;
assign n20662 =  ( n20435 ) ? ( VREG_7_1 ) : ( n20661 ) ;
assign n20663 =  ( n20434 ) ? ( VREG_7_2 ) : ( n20662 ) ;
assign n20664 =  ( n20433 ) ? ( VREG_7_3 ) : ( n20663 ) ;
assign n20665 =  ( n20432 ) ? ( VREG_7_4 ) : ( n20664 ) ;
assign n20666 =  ( n20431 ) ? ( VREG_7_5 ) : ( n20665 ) ;
assign n20667 =  ( n20430 ) ? ( VREG_7_6 ) : ( n20666 ) ;
assign n20668 =  ( n20429 ) ? ( VREG_7_7 ) : ( n20667 ) ;
assign n20669 =  ( n20428 ) ? ( VREG_7_8 ) : ( n20668 ) ;
assign n20670 =  ( n20427 ) ? ( VREG_7_9 ) : ( n20669 ) ;
assign n20671 =  ( n20426 ) ? ( VREG_7_10 ) : ( n20670 ) ;
assign n20672 =  ( n20425 ) ? ( VREG_7_11 ) : ( n20671 ) ;
assign n20673 =  ( n20424 ) ? ( VREG_7_12 ) : ( n20672 ) ;
assign n20674 =  ( n20423 ) ? ( VREG_7_13 ) : ( n20673 ) ;
assign n20675 =  ( n20422 ) ? ( VREG_7_14 ) : ( n20674 ) ;
assign n20676 =  ( n20421 ) ? ( VREG_7_15 ) : ( n20675 ) ;
assign n20677 =  ( n20420 ) ? ( VREG_8_0 ) : ( n20676 ) ;
assign n20678 =  ( n20419 ) ? ( VREG_8_1 ) : ( n20677 ) ;
assign n20679 =  ( n20418 ) ? ( VREG_8_2 ) : ( n20678 ) ;
assign n20680 =  ( n20417 ) ? ( VREG_8_3 ) : ( n20679 ) ;
assign n20681 =  ( n20416 ) ? ( VREG_8_4 ) : ( n20680 ) ;
assign n20682 =  ( n20415 ) ? ( VREG_8_5 ) : ( n20681 ) ;
assign n20683 =  ( n20414 ) ? ( VREG_8_6 ) : ( n20682 ) ;
assign n20684 =  ( n20413 ) ? ( VREG_8_7 ) : ( n20683 ) ;
assign n20685 =  ( n20412 ) ? ( VREG_8_8 ) : ( n20684 ) ;
assign n20686 =  ( n20411 ) ? ( VREG_8_9 ) : ( n20685 ) ;
assign n20687 =  ( n20410 ) ? ( VREG_8_10 ) : ( n20686 ) ;
assign n20688 =  ( n20409 ) ? ( VREG_8_11 ) : ( n20687 ) ;
assign n20689 =  ( n20408 ) ? ( VREG_8_12 ) : ( n20688 ) ;
assign n20690 =  ( n20407 ) ? ( VREG_8_13 ) : ( n20689 ) ;
assign n20691 =  ( n20406 ) ? ( VREG_8_14 ) : ( n20690 ) ;
assign n20692 =  ( n20405 ) ? ( VREG_8_15 ) : ( n20691 ) ;
assign n20693 =  ( n20404 ) ? ( VREG_9_0 ) : ( n20692 ) ;
assign n20694 =  ( n20403 ) ? ( VREG_9_1 ) : ( n20693 ) ;
assign n20695 =  ( n20402 ) ? ( VREG_9_2 ) : ( n20694 ) ;
assign n20696 =  ( n20401 ) ? ( VREG_9_3 ) : ( n20695 ) ;
assign n20697 =  ( n20400 ) ? ( VREG_9_4 ) : ( n20696 ) ;
assign n20698 =  ( n20399 ) ? ( VREG_9_5 ) : ( n20697 ) ;
assign n20699 =  ( n20398 ) ? ( VREG_9_6 ) : ( n20698 ) ;
assign n20700 =  ( n20397 ) ? ( VREG_9_7 ) : ( n20699 ) ;
assign n20701 =  ( n20396 ) ? ( VREG_9_8 ) : ( n20700 ) ;
assign n20702 =  ( n20395 ) ? ( VREG_9_9 ) : ( n20701 ) ;
assign n20703 =  ( n20394 ) ? ( VREG_9_10 ) : ( n20702 ) ;
assign n20704 =  ( n20393 ) ? ( VREG_9_11 ) : ( n20703 ) ;
assign n20705 =  ( n20392 ) ? ( VREG_9_12 ) : ( n20704 ) ;
assign n20706 =  ( n20391 ) ? ( VREG_9_13 ) : ( n20705 ) ;
assign n20707 =  ( n20390 ) ? ( VREG_9_14 ) : ( n20706 ) ;
assign n20708 =  ( n20389 ) ? ( VREG_9_15 ) : ( n20707 ) ;
assign n20709 =  ( n20388 ) ? ( VREG_10_0 ) : ( n20708 ) ;
assign n20710 =  ( n20387 ) ? ( VREG_10_1 ) : ( n20709 ) ;
assign n20711 =  ( n20386 ) ? ( VREG_10_2 ) : ( n20710 ) ;
assign n20712 =  ( n20385 ) ? ( VREG_10_3 ) : ( n20711 ) ;
assign n20713 =  ( n20384 ) ? ( VREG_10_4 ) : ( n20712 ) ;
assign n20714 =  ( n20383 ) ? ( VREG_10_5 ) : ( n20713 ) ;
assign n20715 =  ( n20382 ) ? ( VREG_10_6 ) : ( n20714 ) ;
assign n20716 =  ( n20381 ) ? ( VREG_10_7 ) : ( n20715 ) ;
assign n20717 =  ( n20380 ) ? ( VREG_10_8 ) : ( n20716 ) ;
assign n20718 =  ( n20379 ) ? ( VREG_10_9 ) : ( n20717 ) ;
assign n20719 =  ( n20378 ) ? ( VREG_10_10 ) : ( n20718 ) ;
assign n20720 =  ( n20377 ) ? ( VREG_10_11 ) : ( n20719 ) ;
assign n20721 =  ( n20376 ) ? ( VREG_10_12 ) : ( n20720 ) ;
assign n20722 =  ( n20375 ) ? ( VREG_10_13 ) : ( n20721 ) ;
assign n20723 =  ( n20374 ) ? ( VREG_10_14 ) : ( n20722 ) ;
assign n20724 =  ( n20373 ) ? ( VREG_10_15 ) : ( n20723 ) ;
assign n20725 =  ( n20372 ) ? ( VREG_11_0 ) : ( n20724 ) ;
assign n20726 =  ( n20371 ) ? ( VREG_11_1 ) : ( n20725 ) ;
assign n20727 =  ( n20370 ) ? ( VREG_11_2 ) : ( n20726 ) ;
assign n20728 =  ( n20369 ) ? ( VREG_11_3 ) : ( n20727 ) ;
assign n20729 =  ( n20368 ) ? ( VREG_11_4 ) : ( n20728 ) ;
assign n20730 =  ( n20367 ) ? ( VREG_11_5 ) : ( n20729 ) ;
assign n20731 =  ( n20366 ) ? ( VREG_11_6 ) : ( n20730 ) ;
assign n20732 =  ( n20365 ) ? ( VREG_11_7 ) : ( n20731 ) ;
assign n20733 =  ( n20364 ) ? ( VREG_11_8 ) : ( n20732 ) ;
assign n20734 =  ( n20363 ) ? ( VREG_11_9 ) : ( n20733 ) ;
assign n20735 =  ( n20362 ) ? ( VREG_11_10 ) : ( n20734 ) ;
assign n20736 =  ( n20361 ) ? ( VREG_11_11 ) : ( n20735 ) ;
assign n20737 =  ( n20360 ) ? ( VREG_11_12 ) : ( n20736 ) ;
assign n20738 =  ( n20359 ) ? ( VREG_11_13 ) : ( n20737 ) ;
assign n20739 =  ( n20358 ) ? ( VREG_11_14 ) : ( n20738 ) ;
assign n20740 =  ( n20357 ) ? ( VREG_11_15 ) : ( n20739 ) ;
assign n20741 =  ( n20356 ) ? ( VREG_12_0 ) : ( n20740 ) ;
assign n20742 =  ( n20355 ) ? ( VREG_12_1 ) : ( n20741 ) ;
assign n20743 =  ( n20354 ) ? ( VREG_12_2 ) : ( n20742 ) ;
assign n20744 =  ( n20353 ) ? ( VREG_12_3 ) : ( n20743 ) ;
assign n20745 =  ( n20352 ) ? ( VREG_12_4 ) : ( n20744 ) ;
assign n20746 =  ( n20351 ) ? ( VREG_12_5 ) : ( n20745 ) ;
assign n20747 =  ( n20350 ) ? ( VREG_12_6 ) : ( n20746 ) ;
assign n20748 =  ( n20349 ) ? ( VREG_12_7 ) : ( n20747 ) ;
assign n20749 =  ( n20348 ) ? ( VREG_12_8 ) : ( n20748 ) ;
assign n20750 =  ( n20347 ) ? ( VREG_12_9 ) : ( n20749 ) ;
assign n20751 =  ( n20346 ) ? ( VREG_12_10 ) : ( n20750 ) ;
assign n20752 =  ( n20345 ) ? ( VREG_12_11 ) : ( n20751 ) ;
assign n20753 =  ( n20344 ) ? ( VREG_12_12 ) : ( n20752 ) ;
assign n20754 =  ( n20343 ) ? ( VREG_12_13 ) : ( n20753 ) ;
assign n20755 =  ( n20342 ) ? ( VREG_12_14 ) : ( n20754 ) ;
assign n20756 =  ( n20341 ) ? ( VREG_12_15 ) : ( n20755 ) ;
assign n20757 =  ( n20340 ) ? ( VREG_13_0 ) : ( n20756 ) ;
assign n20758 =  ( n20339 ) ? ( VREG_13_1 ) : ( n20757 ) ;
assign n20759 =  ( n20338 ) ? ( VREG_13_2 ) : ( n20758 ) ;
assign n20760 =  ( n20337 ) ? ( VREG_13_3 ) : ( n20759 ) ;
assign n20761 =  ( n20336 ) ? ( VREG_13_4 ) : ( n20760 ) ;
assign n20762 =  ( n20335 ) ? ( VREG_13_5 ) : ( n20761 ) ;
assign n20763 =  ( n20334 ) ? ( VREG_13_6 ) : ( n20762 ) ;
assign n20764 =  ( n20333 ) ? ( VREG_13_7 ) : ( n20763 ) ;
assign n20765 =  ( n20332 ) ? ( VREG_13_8 ) : ( n20764 ) ;
assign n20766 =  ( n20331 ) ? ( VREG_13_9 ) : ( n20765 ) ;
assign n20767 =  ( n20330 ) ? ( VREG_13_10 ) : ( n20766 ) ;
assign n20768 =  ( n20329 ) ? ( VREG_13_11 ) : ( n20767 ) ;
assign n20769 =  ( n20328 ) ? ( VREG_13_12 ) : ( n20768 ) ;
assign n20770 =  ( n20327 ) ? ( VREG_13_13 ) : ( n20769 ) ;
assign n20771 =  ( n20326 ) ? ( VREG_13_14 ) : ( n20770 ) ;
assign n20772 =  ( n20325 ) ? ( VREG_13_15 ) : ( n20771 ) ;
assign n20773 =  ( n20324 ) ? ( VREG_14_0 ) : ( n20772 ) ;
assign n20774 =  ( n20323 ) ? ( VREG_14_1 ) : ( n20773 ) ;
assign n20775 =  ( n20322 ) ? ( VREG_14_2 ) : ( n20774 ) ;
assign n20776 =  ( n20321 ) ? ( VREG_14_3 ) : ( n20775 ) ;
assign n20777 =  ( n20320 ) ? ( VREG_14_4 ) : ( n20776 ) ;
assign n20778 =  ( n20319 ) ? ( VREG_14_5 ) : ( n20777 ) ;
assign n20779 =  ( n20318 ) ? ( VREG_14_6 ) : ( n20778 ) ;
assign n20780 =  ( n20317 ) ? ( VREG_14_7 ) : ( n20779 ) ;
assign n20781 =  ( n20316 ) ? ( VREG_14_8 ) : ( n20780 ) ;
assign n20782 =  ( n20315 ) ? ( VREG_14_9 ) : ( n20781 ) ;
assign n20783 =  ( n20314 ) ? ( VREG_14_10 ) : ( n20782 ) ;
assign n20784 =  ( n20313 ) ? ( VREG_14_11 ) : ( n20783 ) ;
assign n20785 =  ( n20312 ) ? ( VREG_14_12 ) : ( n20784 ) ;
assign n20786 =  ( n20311 ) ? ( VREG_14_13 ) : ( n20785 ) ;
assign n20787 =  ( n20310 ) ? ( VREG_14_14 ) : ( n20786 ) ;
assign n20788 =  ( n20309 ) ? ( VREG_14_15 ) : ( n20787 ) ;
assign n20789 =  ( n20308 ) ? ( VREG_15_0 ) : ( n20788 ) ;
assign n20790 =  ( n20307 ) ? ( VREG_15_1 ) : ( n20789 ) ;
assign n20791 =  ( n20306 ) ? ( VREG_15_2 ) : ( n20790 ) ;
assign n20792 =  ( n20305 ) ? ( VREG_15_3 ) : ( n20791 ) ;
assign n20793 =  ( n20304 ) ? ( VREG_15_4 ) : ( n20792 ) ;
assign n20794 =  ( n20303 ) ? ( VREG_15_5 ) : ( n20793 ) ;
assign n20795 =  ( n20302 ) ? ( VREG_15_6 ) : ( n20794 ) ;
assign n20796 =  ( n20301 ) ? ( VREG_15_7 ) : ( n20795 ) ;
assign n20797 =  ( n20300 ) ? ( VREG_15_8 ) : ( n20796 ) ;
assign n20798 =  ( n20299 ) ? ( VREG_15_9 ) : ( n20797 ) ;
assign n20799 =  ( n20298 ) ? ( VREG_15_10 ) : ( n20798 ) ;
assign n20800 =  ( n20297 ) ? ( VREG_15_11 ) : ( n20799 ) ;
assign n20801 =  ( n20296 ) ? ( VREG_15_12 ) : ( n20800 ) ;
assign n20802 =  ( n20295 ) ? ( VREG_15_13 ) : ( n20801 ) ;
assign n20803 =  ( n20294 ) ? ( VREG_15_14 ) : ( n20802 ) ;
assign n20804 =  ( n20293 ) ? ( VREG_15_15 ) : ( n20803 ) ;
assign n20805 =  ( n20292 ) ? ( VREG_16_0 ) : ( n20804 ) ;
assign n20806 =  ( n20291 ) ? ( VREG_16_1 ) : ( n20805 ) ;
assign n20807 =  ( n20290 ) ? ( VREG_16_2 ) : ( n20806 ) ;
assign n20808 =  ( n20289 ) ? ( VREG_16_3 ) : ( n20807 ) ;
assign n20809 =  ( n20288 ) ? ( VREG_16_4 ) : ( n20808 ) ;
assign n20810 =  ( n20287 ) ? ( VREG_16_5 ) : ( n20809 ) ;
assign n20811 =  ( n20286 ) ? ( VREG_16_6 ) : ( n20810 ) ;
assign n20812 =  ( n20285 ) ? ( VREG_16_7 ) : ( n20811 ) ;
assign n20813 =  ( n20284 ) ? ( VREG_16_8 ) : ( n20812 ) ;
assign n20814 =  ( n20283 ) ? ( VREG_16_9 ) : ( n20813 ) ;
assign n20815 =  ( n20282 ) ? ( VREG_16_10 ) : ( n20814 ) ;
assign n20816 =  ( n20281 ) ? ( VREG_16_11 ) : ( n20815 ) ;
assign n20817 =  ( n20280 ) ? ( VREG_16_12 ) : ( n20816 ) ;
assign n20818 =  ( n20279 ) ? ( VREG_16_13 ) : ( n20817 ) ;
assign n20819 =  ( n20278 ) ? ( VREG_16_14 ) : ( n20818 ) ;
assign n20820 =  ( n20277 ) ? ( VREG_16_15 ) : ( n20819 ) ;
assign n20821 =  ( n20276 ) ? ( VREG_17_0 ) : ( n20820 ) ;
assign n20822 =  ( n20275 ) ? ( VREG_17_1 ) : ( n20821 ) ;
assign n20823 =  ( n20274 ) ? ( VREG_17_2 ) : ( n20822 ) ;
assign n20824 =  ( n20273 ) ? ( VREG_17_3 ) : ( n20823 ) ;
assign n20825 =  ( n20272 ) ? ( VREG_17_4 ) : ( n20824 ) ;
assign n20826 =  ( n20271 ) ? ( VREG_17_5 ) : ( n20825 ) ;
assign n20827 =  ( n20270 ) ? ( VREG_17_6 ) : ( n20826 ) ;
assign n20828 =  ( n20269 ) ? ( VREG_17_7 ) : ( n20827 ) ;
assign n20829 =  ( n20268 ) ? ( VREG_17_8 ) : ( n20828 ) ;
assign n20830 =  ( n20267 ) ? ( VREG_17_9 ) : ( n20829 ) ;
assign n20831 =  ( n20266 ) ? ( VREG_17_10 ) : ( n20830 ) ;
assign n20832 =  ( n20265 ) ? ( VREG_17_11 ) : ( n20831 ) ;
assign n20833 =  ( n20264 ) ? ( VREG_17_12 ) : ( n20832 ) ;
assign n20834 =  ( n20263 ) ? ( VREG_17_13 ) : ( n20833 ) ;
assign n20835 =  ( n20262 ) ? ( VREG_17_14 ) : ( n20834 ) ;
assign n20836 =  ( n20261 ) ? ( VREG_17_15 ) : ( n20835 ) ;
assign n20837 =  ( n20260 ) ? ( VREG_18_0 ) : ( n20836 ) ;
assign n20838 =  ( n20259 ) ? ( VREG_18_1 ) : ( n20837 ) ;
assign n20839 =  ( n20258 ) ? ( VREG_18_2 ) : ( n20838 ) ;
assign n20840 =  ( n20257 ) ? ( VREG_18_3 ) : ( n20839 ) ;
assign n20841 =  ( n20256 ) ? ( VREG_18_4 ) : ( n20840 ) ;
assign n20842 =  ( n20255 ) ? ( VREG_18_5 ) : ( n20841 ) ;
assign n20843 =  ( n20254 ) ? ( VREG_18_6 ) : ( n20842 ) ;
assign n20844 =  ( n20253 ) ? ( VREG_18_7 ) : ( n20843 ) ;
assign n20845 =  ( n20252 ) ? ( VREG_18_8 ) : ( n20844 ) ;
assign n20846 =  ( n20251 ) ? ( VREG_18_9 ) : ( n20845 ) ;
assign n20847 =  ( n20250 ) ? ( VREG_18_10 ) : ( n20846 ) ;
assign n20848 =  ( n20249 ) ? ( VREG_18_11 ) : ( n20847 ) ;
assign n20849 =  ( n20248 ) ? ( VREG_18_12 ) : ( n20848 ) ;
assign n20850 =  ( n20247 ) ? ( VREG_18_13 ) : ( n20849 ) ;
assign n20851 =  ( n20246 ) ? ( VREG_18_14 ) : ( n20850 ) ;
assign n20852 =  ( n20245 ) ? ( VREG_18_15 ) : ( n20851 ) ;
assign n20853 =  ( n20244 ) ? ( VREG_19_0 ) : ( n20852 ) ;
assign n20854 =  ( n20243 ) ? ( VREG_19_1 ) : ( n20853 ) ;
assign n20855 =  ( n20242 ) ? ( VREG_19_2 ) : ( n20854 ) ;
assign n20856 =  ( n20241 ) ? ( VREG_19_3 ) : ( n20855 ) ;
assign n20857 =  ( n20240 ) ? ( VREG_19_4 ) : ( n20856 ) ;
assign n20858 =  ( n20239 ) ? ( VREG_19_5 ) : ( n20857 ) ;
assign n20859 =  ( n20238 ) ? ( VREG_19_6 ) : ( n20858 ) ;
assign n20860 =  ( n20237 ) ? ( VREG_19_7 ) : ( n20859 ) ;
assign n20861 =  ( n20236 ) ? ( VREG_19_8 ) : ( n20860 ) ;
assign n20862 =  ( n20235 ) ? ( VREG_19_9 ) : ( n20861 ) ;
assign n20863 =  ( n20234 ) ? ( VREG_19_10 ) : ( n20862 ) ;
assign n20864 =  ( n20233 ) ? ( VREG_19_11 ) : ( n20863 ) ;
assign n20865 =  ( n20232 ) ? ( VREG_19_12 ) : ( n20864 ) ;
assign n20866 =  ( n20231 ) ? ( VREG_19_13 ) : ( n20865 ) ;
assign n20867 =  ( n20230 ) ? ( VREG_19_14 ) : ( n20866 ) ;
assign n20868 =  ( n20229 ) ? ( VREG_19_15 ) : ( n20867 ) ;
assign n20869 =  ( n20228 ) ? ( VREG_20_0 ) : ( n20868 ) ;
assign n20870 =  ( n20227 ) ? ( VREG_20_1 ) : ( n20869 ) ;
assign n20871 =  ( n20226 ) ? ( VREG_20_2 ) : ( n20870 ) ;
assign n20872 =  ( n20225 ) ? ( VREG_20_3 ) : ( n20871 ) ;
assign n20873 =  ( n20224 ) ? ( VREG_20_4 ) : ( n20872 ) ;
assign n20874 =  ( n20223 ) ? ( VREG_20_5 ) : ( n20873 ) ;
assign n20875 =  ( n20222 ) ? ( VREG_20_6 ) : ( n20874 ) ;
assign n20876 =  ( n20221 ) ? ( VREG_20_7 ) : ( n20875 ) ;
assign n20877 =  ( n20220 ) ? ( VREG_20_8 ) : ( n20876 ) ;
assign n20878 =  ( n20219 ) ? ( VREG_20_9 ) : ( n20877 ) ;
assign n20879 =  ( n20218 ) ? ( VREG_20_10 ) : ( n20878 ) ;
assign n20880 =  ( n20217 ) ? ( VREG_20_11 ) : ( n20879 ) ;
assign n20881 =  ( n20216 ) ? ( VREG_20_12 ) : ( n20880 ) ;
assign n20882 =  ( n20215 ) ? ( VREG_20_13 ) : ( n20881 ) ;
assign n20883 =  ( n20214 ) ? ( VREG_20_14 ) : ( n20882 ) ;
assign n20884 =  ( n20213 ) ? ( VREG_20_15 ) : ( n20883 ) ;
assign n20885 =  ( n20212 ) ? ( VREG_21_0 ) : ( n20884 ) ;
assign n20886 =  ( n20211 ) ? ( VREG_21_1 ) : ( n20885 ) ;
assign n20887 =  ( n20210 ) ? ( VREG_21_2 ) : ( n20886 ) ;
assign n20888 =  ( n20209 ) ? ( VREG_21_3 ) : ( n20887 ) ;
assign n20889 =  ( n20208 ) ? ( VREG_21_4 ) : ( n20888 ) ;
assign n20890 =  ( n20207 ) ? ( VREG_21_5 ) : ( n20889 ) ;
assign n20891 =  ( n20206 ) ? ( VREG_21_6 ) : ( n20890 ) ;
assign n20892 =  ( n20205 ) ? ( VREG_21_7 ) : ( n20891 ) ;
assign n20893 =  ( n20204 ) ? ( VREG_21_8 ) : ( n20892 ) ;
assign n20894 =  ( n20203 ) ? ( VREG_21_9 ) : ( n20893 ) ;
assign n20895 =  ( n20202 ) ? ( VREG_21_10 ) : ( n20894 ) ;
assign n20896 =  ( n20201 ) ? ( VREG_21_11 ) : ( n20895 ) ;
assign n20897 =  ( n20200 ) ? ( VREG_21_12 ) : ( n20896 ) ;
assign n20898 =  ( n20199 ) ? ( VREG_21_13 ) : ( n20897 ) ;
assign n20899 =  ( n20198 ) ? ( VREG_21_14 ) : ( n20898 ) ;
assign n20900 =  ( n20197 ) ? ( VREG_21_15 ) : ( n20899 ) ;
assign n20901 =  ( n20196 ) ? ( VREG_22_0 ) : ( n20900 ) ;
assign n20902 =  ( n20195 ) ? ( VREG_22_1 ) : ( n20901 ) ;
assign n20903 =  ( n20194 ) ? ( VREG_22_2 ) : ( n20902 ) ;
assign n20904 =  ( n20193 ) ? ( VREG_22_3 ) : ( n20903 ) ;
assign n20905 =  ( n20192 ) ? ( VREG_22_4 ) : ( n20904 ) ;
assign n20906 =  ( n20191 ) ? ( VREG_22_5 ) : ( n20905 ) ;
assign n20907 =  ( n20190 ) ? ( VREG_22_6 ) : ( n20906 ) ;
assign n20908 =  ( n20189 ) ? ( VREG_22_7 ) : ( n20907 ) ;
assign n20909 =  ( n20188 ) ? ( VREG_22_8 ) : ( n20908 ) ;
assign n20910 =  ( n20187 ) ? ( VREG_22_9 ) : ( n20909 ) ;
assign n20911 =  ( n20186 ) ? ( VREG_22_10 ) : ( n20910 ) ;
assign n20912 =  ( n20185 ) ? ( VREG_22_11 ) : ( n20911 ) ;
assign n20913 =  ( n20184 ) ? ( VREG_22_12 ) : ( n20912 ) ;
assign n20914 =  ( n20183 ) ? ( VREG_22_13 ) : ( n20913 ) ;
assign n20915 =  ( n20182 ) ? ( VREG_22_14 ) : ( n20914 ) ;
assign n20916 =  ( n20181 ) ? ( VREG_22_15 ) : ( n20915 ) ;
assign n20917 =  ( n20180 ) ? ( VREG_23_0 ) : ( n20916 ) ;
assign n20918 =  ( n20179 ) ? ( VREG_23_1 ) : ( n20917 ) ;
assign n20919 =  ( n20178 ) ? ( VREG_23_2 ) : ( n20918 ) ;
assign n20920 =  ( n20177 ) ? ( VREG_23_3 ) : ( n20919 ) ;
assign n20921 =  ( n20176 ) ? ( VREG_23_4 ) : ( n20920 ) ;
assign n20922 =  ( n20175 ) ? ( VREG_23_5 ) : ( n20921 ) ;
assign n20923 =  ( n20174 ) ? ( VREG_23_6 ) : ( n20922 ) ;
assign n20924 =  ( n20173 ) ? ( VREG_23_7 ) : ( n20923 ) ;
assign n20925 =  ( n20172 ) ? ( VREG_23_8 ) : ( n20924 ) ;
assign n20926 =  ( n20171 ) ? ( VREG_23_9 ) : ( n20925 ) ;
assign n20927 =  ( n20170 ) ? ( VREG_23_10 ) : ( n20926 ) ;
assign n20928 =  ( n20169 ) ? ( VREG_23_11 ) : ( n20927 ) ;
assign n20929 =  ( n20168 ) ? ( VREG_23_12 ) : ( n20928 ) ;
assign n20930 =  ( n20167 ) ? ( VREG_23_13 ) : ( n20929 ) ;
assign n20931 =  ( n20166 ) ? ( VREG_23_14 ) : ( n20930 ) ;
assign n20932 =  ( n20165 ) ? ( VREG_23_15 ) : ( n20931 ) ;
assign n20933 =  ( n20164 ) ? ( VREG_24_0 ) : ( n20932 ) ;
assign n20934 =  ( n20163 ) ? ( VREG_24_1 ) : ( n20933 ) ;
assign n20935 =  ( n20162 ) ? ( VREG_24_2 ) : ( n20934 ) ;
assign n20936 =  ( n20161 ) ? ( VREG_24_3 ) : ( n20935 ) ;
assign n20937 =  ( n20160 ) ? ( VREG_24_4 ) : ( n20936 ) ;
assign n20938 =  ( n20159 ) ? ( VREG_24_5 ) : ( n20937 ) ;
assign n20939 =  ( n20158 ) ? ( VREG_24_6 ) : ( n20938 ) ;
assign n20940 =  ( n20157 ) ? ( VREG_24_7 ) : ( n20939 ) ;
assign n20941 =  ( n20156 ) ? ( VREG_24_8 ) : ( n20940 ) ;
assign n20942 =  ( n20155 ) ? ( VREG_24_9 ) : ( n20941 ) ;
assign n20943 =  ( n20154 ) ? ( VREG_24_10 ) : ( n20942 ) ;
assign n20944 =  ( n20153 ) ? ( VREG_24_11 ) : ( n20943 ) ;
assign n20945 =  ( n20152 ) ? ( VREG_24_12 ) : ( n20944 ) ;
assign n20946 =  ( n20151 ) ? ( VREG_24_13 ) : ( n20945 ) ;
assign n20947 =  ( n20150 ) ? ( VREG_24_14 ) : ( n20946 ) ;
assign n20948 =  ( n20149 ) ? ( VREG_24_15 ) : ( n20947 ) ;
assign n20949 =  ( n20148 ) ? ( VREG_25_0 ) : ( n20948 ) ;
assign n20950 =  ( n20147 ) ? ( VREG_25_1 ) : ( n20949 ) ;
assign n20951 =  ( n20146 ) ? ( VREG_25_2 ) : ( n20950 ) ;
assign n20952 =  ( n20145 ) ? ( VREG_25_3 ) : ( n20951 ) ;
assign n20953 =  ( n20144 ) ? ( VREG_25_4 ) : ( n20952 ) ;
assign n20954 =  ( n20143 ) ? ( VREG_25_5 ) : ( n20953 ) ;
assign n20955 =  ( n20142 ) ? ( VREG_25_6 ) : ( n20954 ) ;
assign n20956 =  ( n20141 ) ? ( VREG_25_7 ) : ( n20955 ) ;
assign n20957 =  ( n20140 ) ? ( VREG_25_8 ) : ( n20956 ) ;
assign n20958 =  ( n20139 ) ? ( VREG_25_9 ) : ( n20957 ) ;
assign n20959 =  ( n20138 ) ? ( VREG_25_10 ) : ( n20958 ) ;
assign n20960 =  ( n20137 ) ? ( VREG_25_11 ) : ( n20959 ) ;
assign n20961 =  ( n20136 ) ? ( VREG_25_12 ) : ( n20960 ) ;
assign n20962 =  ( n20135 ) ? ( VREG_25_13 ) : ( n20961 ) ;
assign n20963 =  ( n20134 ) ? ( VREG_25_14 ) : ( n20962 ) ;
assign n20964 =  ( n20133 ) ? ( VREG_25_15 ) : ( n20963 ) ;
assign n20965 =  ( n20132 ) ? ( VREG_26_0 ) : ( n20964 ) ;
assign n20966 =  ( n20131 ) ? ( VREG_26_1 ) : ( n20965 ) ;
assign n20967 =  ( n20130 ) ? ( VREG_26_2 ) : ( n20966 ) ;
assign n20968 =  ( n20129 ) ? ( VREG_26_3 ) : ( n20967 ) ;
assign n20969 =  ( n20128 ) ? ( VREG_26_4 ) : ( n20968 ) ;
assign n20970 =  ( n20127 ) ? ( VREG_26_5 ) : ( n20969 ) ;
assign n20971 =  ( n20126 ) ? ( VREG_26_6 ) : ( n20970 ) ;
assign n20972 =  ( n20125 ) ? ( VREG_26_7 ) : ( n20971 ) ;
assign n20973 =  ( n20124 ) ? ( VREG_26_8 ) : ( n20972 ) ;
assign n20974 =  ( n20123 ) ? ( VREG_26_9 ) : ( n20973 ) ;
assign n20975 =  ( n20122 ) ? ( VREG_26_10 ) : ( n20974 ) ;
assign n20976 =  ( n20121 ) ? ( VREG_26_11 ) : ( n20975 ) ;
assign n20977 =  ( n20120 ) ? ( VREG_26_12 ) : ( n20976 ) ;
assign n20978 =  ( n20119 ) ? ( VREG_26_13 ) : ( n20977 ) ;
assign n20979 =  ( n20118 ) ? ( VREG_26_14 ) : ( n20978 ) ;
assign n20980 =  ( n20117 ) ? ( VREG_26_15 ) : ( n20979 ) ;
assign n20981 =  ( n20116 ) ? ( VREG_27_0 ) : ( n20980 ) ;
assign n20982 =  ( n20115 ) ? ( VREG_27_1 ) : ( n20981 ) ;
assign n20983 =  ( n20114 ) ? ( VREG_27_2 ) : ( n20982 ) ;
assign n20984 =  ( n20113 ) ? ( VREG_27_3 ) : ( n20983 ) ;
assign n20985 =  ( n20112 ) ? ( VREG_27_4 ) : ( n20984 ) ;
assign n20986 =  ( n20111 ) ? ( VREG_27_5 ) : ( n20985 ) ;
assign n20987 =  ( n20110 ) ? ( VREG_27_6 ) : ( n20986 ) ;
assign n20988 =  ( n20109 ) ? ( VREG_27_7 ) : ( n20987 ) ;
assign n20989 =  ( n20108 ) ? ( VREG_27_8 ) : ( n20988 ) ;
assign n20990 =  ( n20107 ) ? ( VREG_27_9 ) : ( n20989 ) ;
assign n20991 =  ( n20106 ) ? ( VREG_27_10 ) : ( n20990 ) ;
assign n20992 =  ( n20105 ) ? ( VREG_27_11 ) : ( n20991 ) ;
assign n20993 =  ( n20104 ) ? ( VREG_27_12 ) : ( n20992 ) ;
assign n20994 =  ( n20103 ) ? ( VREG_27_13 ) : ( n20993 ) ;
assign n20995 =  ( n20102 ) ? ( VREG_27_14 ) : ( n20994 ) ;
assign n20996 =  ( n20101 ) ? ( VREG_27_15 ) : ( n20995 ) ;
assign n20997 =  ( n20100 ) ? ( VREG_28_0 ) : ( n20996 ) ;
assign n20998 =  ( n20099 ) ? ( VREG_28_1 ) : ( n20997 ) ;
assign n20999 =  ( n20098 ) ? ( VREG_28_2 ) : ( n20998 ) ;
assign n21000 =  ( n20097 ) ? ( VREG_28_3 ) : ( n20999 ) ;
assign n21001 =  ( n20096 ) ? ( VREG_28_4 ) : ( n21000 ) ;
assign n21002 =  ( n20095 ) ? ( VREG_28_5 ) : ( n21001 ) ;
assign n21003 =  ( n20094 ) ? ( VREG_28_6 ) : ( n21002 ) ;
assign n21004 =  ( n20093 ) ? ( VREG_28_7 ) : ( n21003 ) ;
assign n21005 =  ( n20092 ) ? ( VREG_28_8 ) : ( n21004 ) ;
assign n21006 =  ( n20091 ) ? ( VREG_28_9 ) : ( n21005 ) ;
assign n21007 =  ( n20090 ) ? ( VREG_28_10 ) : ( n21006 ) ;
assign n21008 =  ( n20089 ) ? ( VREG_28_11 ) : ( n21007 ) ;
assign n21009 =  ( n20088 ) ? ( VREG_28_12 ) : ( n21008 ) ;
assign n21010 =  ( n20087 ) ? ( VREG_28_13 ) : ( n21009 ) ;
assign n21011 =  ( n20086 ) ? ( VREG_28_14 ) : ( n21010 ) ;
assign n21012 =  ( n20085 ) ? ( VREG_28_15 ) : ( n21011 ) ;
assign n21013 =  ( n20084 ) ? ( VREG_29_0 ) : ( n21012 ) ;
assign n21014 =  ( n20083 ) ? ( VREG_29_1 ) : ( n21013 ) ;
assign n21015 =  ( n20082 ) ? ( VREG_29_2 ) : ( n21014 ) ;
assign n21016 =  ( n20081 ) ? ( VREG_29_3 ) : ( n21015 ) ;
assign n21017 =  ( n20080 ) ? ( VREG_29_4 ) : ( n21016 ) ;
assign n21018 =  ( n20079 ) ? ( VREG_29_5 ) : ( n21017 ) ;
assign n21019 =  ( n20078 ) ? ( VREG_29_6 ) : ( n21018 ) ;
assign n21020 =  ( n20077 ) ? ( VREG_29_7 ) : ( n21019 ) ;
assign n21021 =  ( n20076 ) ? ( VREG_29_8 ) : ( n21020 ) ;
assign n21022 =  ( n20075 ) ? ( VREG_29_9 ) : ( n21021 ) ;
assign n21023 =  ( n20074 ) ? ( VREG_29_10 ) : ( n21022 ) ;
assign n21024 =  ( n20073 ) ? ( VREG_29_11 ) : ( n21023 ) ;
assign n21025 =  ( n20072 ) ? ( VREG_29_12 ) : ( n21024 ) ;
assign n21026 =  ( n20071 ) ? ( VREG_29_13 ) : ( n21025 ) ;
assign n21027 =  ( n20070 ) ? ( VREG_29_14 ) : ( n21026 ) ;
assign n21028 =  ( n20069 ) ? ( VREG_29_15 ) : ( n21027 ) ;
assign n21029 =  ( n20068 ) ? ( VREG_30_0 ) : ( n21028 ) ;
assign n21030 =  ( n20067 ) ? ( VREG_30_1 ) : ( n21029 ) ;
assign n21031 =  ( n20066 ) ? ( VREG_30_2 ) : ( n21030 ) ;
assign n21032 =  ( n20065 ) ? ( VREG_30_3 ) : ( n21031 ) ;
assign n21033 =  ( n20064 ) ? ( VREG_30_4 ) : ( n21032 ) ;
assign n21034 =  ( n20063 ) ? ( VREG_30_5 ) : ( n21033 ) ;
assign n21035 =  ( n20062 ) ? ( VREG_30_6 ) : ( n21034 ) ;
assign n21036 =  ( n20061 ) ? ( VREG_30_7 ) : ( n21035 ) ;
assign n21037 =  ( n20060 ) ? ( VREG_30_8 ) : ( n21036 ) ;
assign n21038 =  ( n20059 ) ? ( VREG_30_9 ) : ( n21037 ) ;
assign n21039 =  ( n20058 ) ? ( VREG_30_10 ) : ( n21038 ) ;
assign n21040 =  ( n20057 ) ? ( VREG_30_11 ) : ( n21039 ) ;
assign n21041 =  ( n20056 ) ? ( VREG_30_12 ) : ( n21040 ) ;
assign n21042 =  ( n20055 ) ? ( VREG_30_13 ) : ( n21041 ) ;
assign n21043 =  ( n20054 ) ? ( VREG_30_14 ) : ( n21042 ) ;
assign n21044 =  ( n20053 ) ? ( VREG_30_15 ) : ( n21043 ) ;
assign n21045 =  ( n20052 ) ? ( VREG_31_0 ) : ( n21044 ) ;
assign n21046 =  ( n20050 ) ? ( VREG_31_1 ) : ( n21045 ) ;
assign n21047 =  ( n20048 ) ? ( VREG_31_2 ) : ( n21046 ) ;
assign n21048 =  ( n20046 ) ? ( VREG_31_3 ) : ( n21047 ) ;
assign n21049 =  ( n20044 ) ? ( VREG_31_4 ) : ( n21048 ) ;
assign n21050 =  ( n20042 ) ? ( VREG_31_5 ) : ( n21049 ) ;
assign n21051 =  ( n20040 ) ? ( VREG_31_6 ) : ( n21050 ) ;
assign n21052 =  ( n20038 ) ? ( VREG_31_7 ) : ( n21051 ) ;
assign n21053 =  ( n20036 ) ? ( VREG_31_8 ) : ( n21052 ) ;
assign n21054 =  ( n20034 ) ? ( VREG_31_9 ) : ( n21053 ) ;
assign n21055 =  ( n20032 ) ? ( VREG_31_10 ) : ( n21054 ) ;
assign n21056 =  ( n20030 ) ? ( VREG_31_11 ) : ( n21055 ) ;
assign n21057 =  ( n20028 ) ? ( VREG_31_12 ) : ( n21056 ) ;
assign n21058 =  ( n20026 ) ? ( VREG_31_13 ) : ( n21057 ) ;
assign n21059 =  ( n20024 ) ? ( VREG_31_14 ) : ( n21058 ) ;
assign n21060 =  ( n20022 ) ? ( VREG_31_15 ) : ( n21059 ) ;
assign n21061 =  ( n21060 ) + ( n140 )  ;
assign n21062 =  ( n21060 ) - ( n140 )  ;
assign n21063 =  ( n21060 ) & ( n140 )  ;
assign n21064 =  ( n21060 ) | ( n140 )  ;
assign n21065 =  ( ( n21060 ) * ( n140 ))  ;
assign n21066 =  ( n148 ) ? ( n21065 ) : ( VREG_0_3 ) ;
assign n21067 =  ( n146 ) ? ( n21064 ) : ( n21066 ) ;
assign n21068 =  ( n144 ) ? ( n21063 ) : ( n21067 ) ;
assign n21069 =  ( n142 ) ? ( n21062 ) : ( n21068 ) ;
assign n21070 =  ( n10 ) ? ( n21061 ) : ( n21069 ) ;
assign n21071 =  ( n77 ) & ( n20021 )  ;
assign n21072 =  ( n77 ) & ( n20023 )  ;
assign n21073 =  ( n77 ) & ( n20025 )  ;
assign n21074 =  ( n77 ) & ( n20027 )  ;
assign n21075 =  ( n77 ) & ( n20029 )  ;
assign n21076 =  ( n77 ) & ( n20031 )  ;
assign n21077 =  ( n77 ) & ( n20033 )  ;
assign n21078 =  ( n77 ) & ( n20035 )  ;
assign n21079 =  ( n77 ) & ( n20037 )  ;
assign n21080 =  ( n77 ) & ( n20039 )  ;
assign n21081 =  ( n77 ) & ( n20041 )  ;
assign n21082 =  ( n77 ) & ( n20043 )  ;
assign n21083 =  ( n77 ) & ( n20045 )  ;
assign n21084 =  ( n77 ) & ( n20047 )  ;
assign n21085 =  ( n77 ) & ( n20049 )  ;
assign n21086 =  ( n77 ) & ( n20051 )  ;
assign n21087 =  ( n78 ) & ( n20021 )  ;
assign n21088 =  ( n78 ) & ( n20023 )  ;
assign n21089 =  ( n78 ) & ( n20025 )  ;
assign n21090 =  ( n78 ) & ( n20027 )  ;
assign n21091 =  ( n78 ) & ( n20029 )  ;
assign n21092 =  ( n78 ) & ( n20031 )  ;
assign n21093 =  ( n78 ) & ( n20033 )  ;
assign n21094 =  ( n78 ) & ( n20035 )  ;
assign n21095 =  ( n78 ) & ( n20037 )  ;
assign n21096 =  ( n78 ) & ( n20039 )  ;
assign n21097 =  ( n78 ) & ( n20041 )  ;
assign n21098 =  ( n78 ) & ( n20043 )  ;
assign n21099 =  ( n78 ) & ( n20045 )  ;
assign n21100 =  ( n78 ) & ( n20047 )  ;
assign n21101 =  ( n78 ) & ( n20049 )  ;
assign n21102 =  ( n78 ) & ( n20051 )  ;
assign n21103 =  ( n79 ) & ( n20021 )  ;
assign n21104 =  ( n79 ) & ( n20023 )  ;
assign n21105 =  ( n79 ) & ( n20025 )  ;
assign n21106 =  ( n79 ) & ( n20027 )  ;
assign n21107 =  ( n79 ) & ( n20029 )  ;
assign n21108 =  ( n79 ) & ( n20031 )  ;
assign n21109 =  ( n79 ) & ( n20033 )  ;
assign n21110 =  ( n79 ) & ( n20035 )  ;
assign n21111 =  ( n79 ) & ( n20037 )  ;
assign n21112 =  ( n79 ) & ( n20039 )  ;
assign n21113 =  ( n79 ) & ( n20041 )  ;
assign n21114 =  ( n79 ) & ( n20043 )  ;
assign n21115 =  ( n79 ) & ( n20045 )  ;
assign n21116 =  ( n79 ) & ( n20047 )  ;
assign n21117 =  ( n79 ) & ( n20049 )  ;
assign n21118 =  ( n79 ) & ( n20051 )  ;
assign n21119 =  ( n80 ) & ( n20021 )  ;
assign n21120 =  ( n80 ) & ( n20023 )  ;
assign n21121 =  ( n80 ) & ( n20025 )  ;
assign n21122 =  ( n80 ) & ( n20027 )  ;
assign n21123 =  ( n80 ) & ( n20029 )  ;
assign n21124 =  ( n80 ) & ( n20031 )  ;
assign n21125 =  ( n80 ) & ( n20033 )  ;
assign n21126 =  ( n80 ) & ( n20035 )  ;
assign n21127 =  ( n80 ) & ( n20037 )  ;
assign n21128 =  ( n80 ) & ( n20039 )  ;
assign n21129 =  ( n80 ) & ( n20041 )  ;
assign n21130 =  ( n80 ) & ( n20043 )  ;
assign n21131 =  ( n80 ) & ( n20045 )  ;
assign n21132 =  ( n80 ) & ( n20047 )  ;
assign n21133 =  ( n80 ) & ( n20049 )  ;
assign n21134 =  ( n80 ) & ( n20051 )  ;
assign n21135 =  ( n81 ) & ( n20021 )  ;
assign n21136 =  ( n81 ) & ( n20023 )  ;
assign n21137 =  ( n81 ) & ( n20025 )  ;
assign n21138 =  ( n81 ) & ( n20027 )  ;
assign n21139 =  ( n81 ) & ( n20029 )  ;
assign n21140 =  ( n81 ) & ( n20031 )  ;
assign n21141 =  ( n81 ) & ( n20033 )  ;
assign n21142 =  ( n81 ) & ( n20035 )  ;
assign n21143 =  ( n81 ) & ( n20037 )  ;
assign n21144 =  ( n81 ) & ( n20039 )  ;
assign n21145 =  ( n81 ) & ( n20041 )  ;
assign n21146 =  ( n81 ) & ( n20043 )  ;
assign n21147 =  ( n81 ) & ( n20045 )  ;
assign n21148 =  ( n81 ) & ( n20047 )  ;
assign n21149 =  ( n81 ) & ( n20049 )  ;
assign n21150 =  ( n81 ) & ( n20051 )  ;
assign n21151 =  ( n82 ) & ( n20021 )  ;
assign n21152 =  ( n82 ) & ( n20023 )  ;
assign n21153 =  ( n82 ) & ( n20025 )  ;
assign n21154 =  ( n82 ) & ( n20027 )  ;
assign n21155 =  ( n82 ) & ( n20029 )  ;
assign n21156 =  ( n82 ) & ( n20031 )  ;
assign n21157 =  ( n82 ) & ( n20033 )  ;
assign n21158 =  ( n82 ) & ( n20035 )  ;
assign n21159 =  ( n82 ) & ( n20037 )  ;
assign n21160 =  ( n82 ) & ( n20039 )  ;
assign n21161 =  ( n82 ) & ( n20041 )  ;
assign n21162 =  ( n82 ) & ( n20043 )  ;
assign n21163 =  ( n82 ) & ( n20045 )  ;
assign n21164 =  ( n82 ) & ( n20047 )  ;
assign n21165 =  ( n82 ) & ( n20049 )  ;
assign n21166 =  ( n82 ) & ( n20051 )  ;
assign n21167 =  ( n83 ) & ( n20021 )  ;
assign n21168 =  ( n83 ) & ( n20023 )  ;
assign n21169 =  ( n83 ) & ( n20025 )  ;
assign n21170 =  ( n83 ) & ( n20027 )  ;
assign n21171 =  ( n83 ) & ( n20029 )  ;
assign n21172 =  ( n83 ) & ( n20031 )  ;
assign n21173 =  ( n83 ) & ( n20033 )  ;
assign n21174 =  ( n83 ) & ( n20035 )  ;
assign n21175 =  ( n83 ) & ( n20037 )  ;
assign n21176 =  ( n83 ) & ( n20039 )  ;
assign n21177 =  ( n83 ) & ( n20041 )  ;
assign n21178 =  ( n83 ) & ( n20043 )  ;
assign n21179 =  ( n83 ) & ( n20045 )  ;
assign n21180 =  ( n83 ) & ( n20047 )  ;
assign n21181 =  ( n83 ) & ( n20049 )  ;
assign n21182 =  ( n83 ) & ( n20051 )  ;
assign n21183 =  ( n84 ) & ( n20021 )  ;
assign n21184 =  ( n84 ) & ( n20023 )  ;
assign n21185 =  ( n84 ) & ( n20025 )  ;
assign n21186 =  ( n84 ) & ( n20027 )  ;
assign n21187 =  ( n84 ) & ( n20029 )  ;
assign n21188 =  ( n84 ) & ( n20031 )  ;
assign n21189 =  ( n84 ) & ( n20033 )  ;
assign n21190 =  ( n84 ) & ( n20035 )  ;
assign n21191 =  ( n84 ) & ( n20037 )  ;
assign n21192 =  ( n84 ) & ( n20039 )  ;
assign n21193 =  ( n84 ) & ( n20041 )  ;
assign n21194 =  ( n84 ) & ( n20043 )  ;
assign n21195 =  ( n84 ) & ( n20045 )  ;
assign n21196 =  ( n84 ) & ( n20047 )  ;
assign n21197 =  ( n84 ) & ( n20049 )  ;
assign n21198 =  ( n84 ) & ( n20051 )  ;
assign n21199 =  ( n85 ) & ( n20021 )  ;
assign n21200 =  ( n85 ) & ( n20023 )  ;
assign n21201 =  ( n85 ) & ( n20025 )  ;
assign n21202 =  ( n85 ) & ( n20027 )  ;
assign n21203 =  ( n85 ) & ( n20029 )  ;
assign n21204 =  ( n85 ) & ( n20031 )  ;
assign n21205 =  ( n85 ) & ( n20033 )  ;
assign n21206 =  ( n85 ) & ( n20035 )  ;
assign n21207 =  ( n85 ) & ( n20037 )  ;
assign n21208 =  ( n85 ) & ( n20039 )  ;
assign n21209 =  ( n85 ) & ( n20041 )  ;
assign n21210 =  ( n85 ) & ( n20043 )  ;
assign n21211 =  ( n85 ) & ( n20045 )  ;
assign n21212 =  ( n85 ) & ( n20047 )  ;
assign n21213 =  ( n85 ) & ( n20049 )  ;
assign n21214 =  ( n85 ) & ( n20051 )  ;
assign n21215 =  ( n86 ) & ( n20021 )  ;
assign n21216 =  ( n86 ) & ( n20023 )  ;
assign n21217 =  ( n86 ) & ( n20025 )  ;
assign n21218 =  ( n86 ) & ( n20027 )  ;
assign n21219 =  ( n86 ) & ( n20029 )  ;
assign n21220 =  ( n86 ) & ( n20031 )  ;
assign n21221 =  ( n86 ) & ( n20033 )  ;
assign n21222 =  ( n86 ) & ( n20035 )  ;
assign n21223 =  ( n86 ) & ( n20037 )  ;
assign n21224 =  ( n86 ) & ( n20039 )  ;
assign n21225 =  ( n86 ) & ( n20041 )  ;
assign n21226 =  ( n86 ) & ( n20043 )  ;
assign n21227 =  ( n86 ) & ( n20045 )  ;
assign n21228 =  ( n86 ) & ( n20047 )  ;
assign n21229 =  ( n86 ) & ( n20049 )  ;
assign n21230 =  ( n86 ) & ( n20051 )  ;
assign n21231 =  ( n87 ) & ( n20021 )  ;
assign n21232 =  ( n87 ) & ( n20023 )  ;
assign n21233 =  ( n87 ) & ( n20025 )  ;
assign n21234 =  ( n87 ) & ( n20027 )  ;
assign n21235 =  ( n87 ) & ( n20029 )  ;
assign n21236 =  ( n87 ) & ( n20031 )  ;
assign n21237 =  ( n87 ) & ( n20033 )  ;
assign n21238 =  ( n87 ) & ( n20035 )  ;
assign n21239 =  ( n87 ) & ( n20037 )  ;
assign n21240 =  ( n87 ) & ( n20039 )  ;
assign n21241 =  ( n87 ) & ( n20041 )  ;
assign n21242 =  ( n87 ) & ( n20043 )  ;
assign n21243 =  ( n87 ) & ( n20045 )  ;
assign n21244 =  ( n87 ) & ( n20047 )  ;
assign n21245 =  ( n87 ) & ( n20049 )  ;
assign n21246 =  ( n87 ) & ( n20051 )  ;
assign n21247 =  ( n88 ) & ( n20021 )  ;
assign n21248 =  ( n88 ) & ( n20023 )  ;
assign n21249 =  ( n88 ) & ( n20025 )  ;
assign n21250 =  ( n88 ) & ( n20027 )  ;
assign n21251 =  ( n88 ) & ( n20029 )  ;
assign n21252 =  ( n88 ) & ( n20031 )  ;
assign n21253 =  ( n88 ) & ( n20033 )  ;
assign n21254 =  ( n88 ) & ( n20035 )  ;
assign n21255 =  ( n88 ) & ( n20037 )  ;
assign n21256 =  ( n88 ) & ( n20039 )  ;
assign n21257 =  ( n88 ) & ( n20041 )  ;
assign n21258 =  ( n88 ) & ( n20043 )  ;
assign n21259 =  ( n88 ) & ( n20045 )  ;
assign n21260 =  ( n88 ) & ( n20047 )  ;
assign n21261 =  ( n88 ) & ( n20049 )  ;
assign n21262 =  ( n88 ) & ( n20051 )  ;
assign n21263 =  ( n89 ) & ( n20021 )  ;
assign n21264 =  ( n89 ) & ( n20023 )  ;
assign n21265 =  ( n89 ) & ( n20025 )  ;
assign n21266 =  ( n89 ) & ( n20027 )  ;
assign n21267 =  ( n89 ) & ( n20029 )  ;
assign n21268 =  ( n89 ) & ( n20031 )  ;
assign n21269 =  ( n89 ) & ( n20033 )  ;
assign n21270 =  ( n89 ) & ( n20035 )  ;
assign n21271 =  ( n89 ) & ( n20037 )  ;
assign n21272 =  ( n89 ) & ( n20039 )  ;
assign n21273 =  ( n89 ) & ( n20041 )  ;
assign n21274 =  ( n89 ) & ( n20043 )  ;
assign n21275 =  ( n89 ) & ( n20045 )  ;
assign n21276 =  ( n89 ) & ( n20047 )  ;
assign n21277 =  ( n89 ) & ( n20049 )  ;
assign n21278 =  ( n89 ) & ( n20051 )  ;
assign n21279 =  ( n90 ) & ( n20021 )  ;
assign n21280 =  ( n90 ) & ( n20023 )  ;
assign n21281 =  ( n90 ) & ( n20025 )  ;
assign n21282 =  ( n90 ) & ( n20027 )  ;
assign n21283 =  ( n90 ) & ( n20029 )  ;
assign n21284 =  ( n90 ) & ( n20031 )  ;
assign n21285 =  ( n90 ) & ( n20033 )  ;
assign n21286 =  ( n90 ) & ( n20035 )  ;
assign n21287 =  ( n90 ) & ( n20037 )  ;
assign n21288 =  ( n90 ) & ( n20039 )  ;
assign n21289 =  ( n90 ) & ( n20041 )  ;
assign n21290 =  ( n90 ) & ( n20043 )  ;
assign n21291 =  ( n90 ) & ( n20045 )  ;
assign n21292 =  ( n90 ) & ( n20047 )  ;
assign n21293 =  ( n90 ) & ( n20049 )  ;
assign n21294 =  ( n90 ) & ( n20051 )  ;
assign n21295 =  ( n91 ) & ( n20021 )  ;
assign n21296 =  ( n91 ) & ( n20023 )  ;
assign n21297 =  ( n91 ) & ( n20025 )  ;
assign n21298 =  ( n91 ) & ( n20027 )  ;
assign n21299 =  ( n91 ) & ( n20029 )  ;
assign n21300 =  ( n91 ) & ( n20031 )  ;
assign n21301 =  ( n91 ) & ( n20033 )  ;
assign n21302 =  ( n91 ) & ( n20035 )  ;
assign n21303 =  ( n91 ) & ( n20037 )  ;
assign n21304 =  ( n91 ) & ( n20039 )  ;
assign n21305 =  ( n91 ) & ( n20041 )  ;
assign n21306 =  ( n91 ) & ( n20043 )  ;
assign n21307 =  ( n91 ) & ( n20045 )  ;
assign n21308 =  ( n91 ) & ( n20047 )  ;
assign n21309 =  ( n91 ) & ( n20049 )  ;
assign n21310 =  ( n91 ) & ( n20051 )  ;
assign n21311 =  ( n92 ) & ( n20021 )  ;
assign n21312 =  ( n92 ) & ( n20023 )  ;
assign n21313 =  ( n92 ) & ( n20025 )  ;
assign n21314 =  ( n92 ) & ( n20027 )  ;
assign n21315 =  ( n92 ) & ( n20029 )  ;
assign n21316 =  ( n92 ) & ( n20031 )  ;
assign n21317 =  ( n92 ) & ( n20033 )  ;
assign n21318 =  ( n92 ) & ( n20035 )  ;
assign n21319 =  ( n92 ) & ( n20037 )  ;
assign n21320 =  ( n92 ) & ( n20039 )  ;
assign n21321 =  ( n92 ) & ( n20041 )  ;
assign n21322 =  ( n92 ) & ( n20043 )  ;
assign n21323 =  ( n92 ) & ( n20045 )  ;
assign n21324 =  ( n92 ) & ( n20047 )  ;
assign n21325 =  ( n92 ) & ( n20049 )  ;
assign n21326 =  ( n92 ) & ( n20051 )  ;
assign n21327 =  ( n93 ) & ( n20021 )  ;
assign n21328 =  ( n93 ) & ( n20023 )  ;
assign n21329 =  ( n93 ) & ( n20025 )  ;
assign n21330 =  ( n93 ) & ( n20027 )  ;
assign n21331 =  ( n93 ) & ( n20029 )  ;
assign n21332 =  ( n93 ) & ( n20031 )  ;
assign n21333 =  ( n93 ) & ( n20033 )  ;
assign n21334 =  ( n93 ) & ( n20035 )  ;
assign n21335 =  ( n93 ) & ( n20037 )  ;
assign n21336 =  ( n93 ) & ( n20039 )  ;
assign n21337 =  ( n93 ) & ( n20041 )  ;
assign n21338 =  ( n93 ) & ( n20043 )  ;
assign n21339 =  ( n93 ) & ( n20045 )  ;
assign n21340 =  ( n93 ) & ( n20047 )  ;
assign n21341 =  ( n93 ) & ( n20049 )  ;
assign n21342 =  ( n93 ) & ( n20051 )  ;
assign n21343 =  ( n94 ) & ( n20021 )  ;
assign n21344 =  ( n94 ) & ( n20023 )  ;
assign n21345 =  ( n94 ) & ( n20025 )  ;
assign n21346 =  ( n94 ) & ( n20027 )  ;
assign n21347 =  ( n94 ) & ( n20029 )  ;
assign n21348 =  ( n94 ) & ( n20031 )  ;
assign n21349 =  ( n94 ) & ( n20033 )  ;
assign n21350 =  ( n94 ) & ( n20035 )  ;
assign n21351 =  ( n94 ) & ( n20037 )  ;
assign n21352 =  ( n94 ) & ( n20039 )  ;
assign n21353 =  ( n94 ) & ( n20041 )  ;
assign n21354 =  ( n94 ) & ( n20043 )  ;
assign n21355 =  ( n94 ) & ( n20045 )  ;
assign n21356 =  ( n94 ) & ( n20047 )  ;
assign n21357 =  ( n94 ) & ( n20049 )  ;
assign n21358 =  ( n94 ) & ( n20051 )  ;
assign n21359 =  ( n95 ) & ( n20021 )  ;
assign n21360 =  ( n95 ) & ( n20023 )  ;
assign n21361 =  ( n95 ) & ( n20025 )  ;
assign n21362 =  ( n95 ) & ( n20027 )  ;
assign n21363 =  ( n95 ) & ( n20029 )  ;
assign n21364 =  ( n95 ) & ( n20031 )  ;
assign n21365 =  ( n95 ) & ( n20033 )  ;
assign n21366 =  ( n95 ) & ( n20035 )  ;
assign n21367 =  ( n95 ) & ( n20037 )  ;
assign n21368 =  ( n95 ) & ( n20039 )  ;
assign n21369 =  ( n95 ) & ( n20041 )  ;
assign n21370 =  ( n95 ) & ( n20043 )  ;
assign n21371 =  ( n95 ) & ( n20045 )  ;
assign n21372 =  ( n95 ) & ( n20047 )  ;
assign n21373 =  ( n95 ) & ( n20049 )  ;
assign n21374 =  ( n95 ) & ( n20051 )  ;
assign n21375 =  ( n96 ) & ( n20021 )  ;
assign n21376 =  ( n96 ) & ( n20023 )  ;
assign n21377 =  ( n96 ) & ( n20025 )  ;
assign n21378 =  ( n96 ) & ( n20027 )  ;
assign n21379 =  ( n96 ) & ( n20029 )  ;
assign n21380 =  ( n96 ) & ( n20031 )  ;
assign n21381 =  ( n96 ) & ( n20033 )  ;
assign n21382 =  ( n96 ) & ( n20035 )  ;
assign n21383 =  ( n96 ) & ( n20037 )  ;
assign n21384 =  ( n96 ) & ( n20039 )  ;
assign n21385 =  ( n96 ) & ( n20041 )  ;
assign n21386 =  ( n96 ) & ( n20043 )  ;
assign n21387 =  ( n96 ) & ( n20045 )  ;
assign n21388 =  ( n96 ) & ( n20047 )  ;
assign n21389 =  ( n96 ) & ( n20049 )  ;
assign n21390 =  ( n96 ) & ( n20051 )  ;
assign n21391 =  ( n97 ) & ( n20021 )  ;
assign n21392 =  ( n97 ) & ( n20023 )  ;
assign n21393 =  ( n97 ) & ( n20025 )  ;
assign n21394 =  ( n97 ) & ( n20027 )  ;
assign n21395 =  ( n97 ) & ( n20029 )  ;
assign n21396 =  ( n97 ) & ( n20031 )  ;
assign n21397 =  ( n97 ) & ( n20033 )  ;
assign n21398 =  ( n97 ) & ( n20035 )  ;
assign n21399 =  ( n97 ) & ( n20037 )  ;
assign n21400 =  ( n97 ) & ( n20039 )  ;
assign n21401 =  ( n97 ) & ( n20041 )  ;
assign n21402 =  ( n97 ) & ( n20043 )  ;
assign n21403 =  ( n97 ) & ( n20045 )  ;
assign n21404 =  ( n97 ) & ( n20047 )  ;
assign n21405 =  ( n97 ) & ( n20049 )  ;
assign n21406 =  ( n97 ) & ( n20051 )  ;
assign n21407 =  ( n98 ) & ( n20021 )  ;
assign n21408 =  ( n98 ) & ( n20023 )  ;
assign n21409 =  ( n98 ) & ( n20025 )  ;
assign n21410 =  ( n98 ) & ( n20027 )  ;
assign n21411 =  ( n98 ) & ( n20029 )  ;
assign n21412 =  ( n98 ) & ( n20031 )  ;
assign n21413 =  ( n98 ) & ( n20033 )  ;
assign n21414 =  ( n98 ) & ( n20035 )  ;
assign n21415 =  ( n98 ) & ( n20037 )  ;
assign n21416 =  ( n98 ) & ( n20039 )  ;
assign n21417 =  ( n98 ) & ( n20041 )  ;
assign n21418 =  ( n98 ) & ( n20043 )  ;
assign n21419 =  ( n98 ) & ( n20045 )  ;
assign n21420 =  ( n98 ) & ( n20047 )  ;
assign n21421 =  ( n98 ) & ( n20049 )  ;
assign n21422 =  ( n98 ) & ( n20051 )  ;
assign n21423 =  ( n99 ) & ( n20021 )  ;
assign n21424 =  ( n99 ) & ( n20023 )  ;
assign n21425 =  ( n99 ) & ( n20025 )  ;
assign n21426 =  ( n99 ) & ( n20027 )  ;
assign n21427 =  ( n99 ) & ( n20029 )  ;
assign n21428 =  ( n99 ) & ( n20031 )  ;
assign n21429 =  ( n99 ) & ( n20033 )  ;
assign n21430 =  ( n99 ) & ( n20035 )  ;
assign n21431 =  ( n99 ) & ( n20037 )  ;
assign n21432 =  ( n99 ) & ( n20039 )  ;
assign n21433 =  ( n99 ) & ( n20041 )  ;
assign n21434 =  ( n99 ) & ( n20043 )  ;
assign n21435 =  ( n99 ) & ( n20045 )  ;
assign n21436 =  ( n99 ) & ( n20047 )  ;
assign n21437 =  ( n99 ) & ( n20049 )  ;
assign n21438 =  ( n99 ) & ( n20051 )  ;
assign n21439 =  ( n100 ) & ( n20021 )  ;
assign n21440 =  ( n100 ) & ( n20023 )  ;
assign n21441 =  ( n100 ) & ( n20025 )  ;
assign n21442 =  ( n100 ) & ( n20027 )  ;
assign n21443 =  ( n100 ) & ( n20029 )  ;
assign n21444 =  ( n100 ) & ( n20031 )  ;
assign n21445 =  ( n100 ) & ( n20033 )  ;
assign n21446 =  ( n100 ) & ( n20035 )  ;
assign n21447 =  ( n100 ) & ( n20037 )  ;
assign n21448 =  ( n100 ) & ( n20039 )  ;
assign n21449 =  ( n100 ) & ( n20041 )  ;
assign n21450 =  ( n100 ) & ( n20043 )  ;
assign n21451 =  ( n100 ) & ( n20045 )  ;
assign n21452 =  ( n100 ) & ( n20047 )  ;
assign n21453 =  ( n100 ) & ( n20049 )  ;
assign n21454 =  ( n100 ) & ( n20051 )  ;
assign n21455 =  ( n101 ) & ( n20021 )  ;
assign n21456 =  ( n101 ) & ( n20023 )  ;
assign n21457 =  ( n101 ) & ( n20025 )  ;
assign n21458 =  ( n101 ) & ( n20027 )  ;
assign n21459 =  ( n101 ) & ( n20029 )  ;
assign n21460 =  ( n101 ) & ( n20031 )  ;
assign n21461 =  ( n101 ) & ( n20033 )  ;
assign n21462 =  ( n101 ) & ( n20035 )  ;
assign n21463 =  ( n101 ) & ( n20037 )  ;
assign n21464 =  ( n101 ) & ( n20039 )  ;
assign n21465 =  ( n101 ) & ( n20041 )  ;
assign n21466 =  ( n101 ) & ( n20043 )  ;
assign n21467 =  ( n101 ) & ( n20045 )  ;
assign n21468 =  ( n101 ) & ( n20047 )  ;
assign n21469 =  ( n101 ) & ( n20049 )  ;
assign n21470 =  ( n101 ) & ( n20051 )  ;
assign n21471 =  ( n102 ) & ( n20021 )  ;
assign n21472 =  ( n102 ) & ( n20023 )  ;
assign n21473 =  ( n102 ) & ( n20025 )  ;
assign n21474 =  ( n102 ) & ( n20027 )  ;
assign n21475 =  ( n102 ) & ( n20029 )  ;
assign n21476 =  ( n102 ) & ( n20031 )  ;
assign n21477 =  ( n102 ) & ( n20033 )  ;
assign n21478 =  ( n102 ) & ( n20035 )  ;
assign n21479 =  ( n102 ) & ( n20037 )  ;
assign n21480 =  ( n102 ) & ( n20039 )  ;
assign n21481 =  ( n102 ) & ( n20041 )  ;
assign n21482 =  ( n102 ) & ( n20043 )  ;
assign n21483 =  ( n102 ) & ( n20045 )  ;
assign n21484 =  ( n102 ) & ( n20047 )  ;
assign n21485 =  ( n102 ) & ( n20049 )  ;
assign n21486 =  ( n102 ) & ( n20051 )  ;
assign n21487 =  ( n103 ) & ( n20021 )  ;
assign n21488 =  ( n103 ) & ( n20023 )  ;
assign n21489 =  ( n103 ) & ( n20025 )  ;
assign n21490 =  ( n103 ) & ( n20027 )  ;
assign n21491 =  ( n103 ) & ( n20029 )  ;
assign n21492 =  ( n103 ) & ( n20031 )  ;
assign n21493 =  ( n103 ) & ( n20033 )  ;
assign n21494 =  ( n103 ) & ( n20035 )  ;
assign n21495 =  ( n103 ) & ( n20037 )  ;
assign n21496 =  ( n103 ) & ( n20039 )  ;
assign n21497 =  ( n103 ) & ( n20041 )  ;
assign n21498 =  ( n103 ) & ( n20043 )  ;
assign n21499 =  ( n103 ) & ( n20045 )  ;
assign n21500 =  ( n103 ) & ( n20047 )  ;
assign n21501 =  ( n103 ) & ( n20049 )  ;
assign n21502 =  ( n103 ) & ( n20051 )  ;
assign n21503 =  ( n104 ) & ( n20021 )  ;
assign n21504 =  ( n104 ) & ( n20023 )  ;
assign n21505 =  ( n104 ) & ( n20025 )  ;
assign n21506 =  ( n104 ) & ( n20027 )  ;
assign n21507 =  ( n104 ) & ( n20029 )  ;
assign n21508 =  ( n104 ) & ( n20031 )  ;
assign n21509 =  ( n104 ) & ( n20033 )  ;
assign n21510 =  ( n104 ) & ( n20035 )  ;
assign n21511 =  ( n104 ) & ( n20037 )  ;
assign n21512 =  ( n104 ) & ( n20039 )  ;
assign n21513 =  ( n104 ) & ( n20041 )  ;
assign n21514 =  ( n104 ) & ( n20043 )  ;
assign n21515 =  ( n104 ) & ( n20045 )  ;
assign n21516 =  ( n104 ) & ( n20047 )  ;
assign n21517 =  ( n104 ) & ( n20049 )  ;
assign n21518 =  ( n104 ) & ( n20051 )  ;
assign n21519 =  ( n105 ) & ( n20021 )  ;
assign n21520 =  ( n105 ) & ( n20023 )  ;
assign n21521 =  ( n105 ) & ( n20025 )  ;
assign n21522 =  ( n105 ) & ( n20027 )  ;
assign n21523 =  ( n105 ) & ( n20029 )  ;
assign n21524 =  ( n105 ) & ( n20031 )  ;
assign n21525 =  ( n105 ) & ( n20033 )  ;
assign n21526 =  ( n105 ) & ( n20035 )  ;
assign n21527 =  ( n105 ) & ( n20037 )  ;
assign n21528 =  ( n105 ) & ( n20039 )  ;
assign n21529 =  ( n105 ) & ( n20041 )  ;
assign n21530 =  ( n105 ) & ( n20043 )  ;
assign n21531 =  ( n105 ) & ( n20045 )  ;
assign n21532 =  ( n105 ) & ( n20047 )  ;
assign n21533 =  ( n105 ) & ( n20049 )  ;
assign n21534 =  ( n105 ) & ( n20051 )  ;
assign n21535 =  ( n106 ) & ( n20021 )  ;
assign n21536 =  ( n106 ) & ( n20023 )  ;
assign n21537 =  ( n106 ) & ( n20025 )  ;
assign n21538 =  ( n106 ) & ( n20027 )  ;
assign n21539 =  ( n106 ) & ( n20029 )  ;
assign n21540 =  ( n106 ) & ( n20031 )  ;
assign n21541 =  ( n106 ) & ( n20033 )  ;
assign n21542 =  ( n106 ) & ( n20035 )  ;
assign n21543 =  ( n106 ) & ( n20037 )  ;
assign n21544 =  ( n106 ) & ( n20039 )  ;
assign n21545 =  ( n106 ) & ( n20041 )  ;
assign n21546 =  ( n106 ) & ( n20043 )  ;
assign n21547 =  ( n106 ) & ( n20045 )  ;
assign n21548 =  ( n106 ) & ( n20047 )  ;
assign n21549 =  ( n106 ) & ( n20049 )  ;
assign n21550 =  ( n106 ) & ( n20051 )  ;
assign n21551 =  ( n107 ) & ( n20021 )  ;
assign n21552 =  ( n107 ) & ( n20023 )  ;
assign n21553 =  ( n107 ) & ( n20025 )  ;
assign n21554 =  ( n107 ) & ( n20027 )  ;
assign n21555 =  ( n107 ) & ( n20029 )  ;
assign n21556 =  ( n107 ) & ( n20031 )  ;
assign n21557 =  ( n107 ) & ( n20033 )  ;
assign n21558 =  ( n107 ) & ( n20035 )  ;
assign n21559 =  ( n107 ) & ( n20037 )  ;
assign n21560 =  ( n107 ) & ( n20039 )  ;
assign n21561 =  ( n107 ) & ( n20041 )  ;
assign n21562 =  ( n107 ) & ( n20043 )  ;
assign n21563 =  ( n107 ) & ( n20045 )  ;
assign n21564 =  ( n107 ) & ( n20047 )  ;
assign n21565 =  ( n107 ) & ( n20049 )  ;
assign n21566 =  ( n107 ) & ( n20051 )  ;
assign n21567 =  ( n108 ) & ( n20021 )  ;
assign n21568 =  ( n108 ) & ( n20023 )  ;
assign n21569 =  ( n108 ) & ( n20025 )  ;
assign n21570 =  ( n108 ) & ( n20027 )  ;
assign n21571 =  ( n108 ) & ( n20029 )  ;
assign n21572 =  ( n108 ) & ( n20031 )  ;
assign n21573 =  ( n108 ) & ( n20033 )  ;
assign n21574 =  ( n108 ) & ( n20035 )  ;
assign n21575 =  ( n108 ) & ( n20037 )  ;
assign n21576 =  ( n108 ) & ( n20039 )  ;
assign n21577 =  ( n108 ) & ( n20041 )  ;
assign n21578 =  ( n108 ) & ( n20043 )  ;
assign n21579 =  ( n108 ) & ( n20045 )  ;
assign n21580 =  ( n108 ) & ( n20047 )  ;
assign n21581 =  ( n108 ) & ( n20049 )  ;
assign n21582 =  ( n108 ) & ( n20051 )  ;
assign n21583 =  ( n21582 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n21584 =  ( n21581 ) ? ( VREG_0_1 ) : ( n21583 ) ;
assign n21585 =  ( n21580 ) ? ( VREG_0_2 ) : ( n21584 ) ;
assign n21586 =  ( n21579 ) ? ( VREG_0_3 ) : ( n21585 ) ;
assign n21587 =  ( n21578 ) ? ( VREG_0_4 ) : ( n21586 ) ;
assign n21588 =  ( n21577 ) ? ( VREG_0_5 ) : ( n21587 ) ;
assign n21589 =  ( n21576 ) ? ( VREG_0_6 ) : ( n21588 ) ;
assign n21590 =  ( n21575 ) ? ( VREG_0_7 ) : ( n21589 ) ;
assign n21591 =  ( n21574 ) ? ( VREG_0_8 ) : ( n21590 ) ;
assign n21592 =  ( n21573 ) ? ( VREG_0_9 ) : ( n21591 ) ;
assign n21593 =  ( n21572 ) ? ( VREG_0_10 ) : ( n21592 ) ;
assign n21594 =  ( n21571 ) ? ( VREG_0_11 ) : ( n21593 ) ;
assign n21595 =  ( n21570 ) ? ( VREG_0_12 ) : ( n21594 ) ;
assign n21596 =  ( n21569 ) ? ( VREG_0_13 ) : ( n21595 ) ;
assign n21597 =  ( n21568 ) ? ( VREG_0_14 ) : ( n21596 ) ;
assign n21598 =  ( n21567 ) ? ( VREG_0_15 ) : ( n21597 ) ;
assign n21599 =  ( n21566 ) ? ( VREG_1_0 ) : ( n21598 ) ;
assign n21600 =  ( n21565 ) ? ( VREG_1_1 ) : ( n21599 ) ;
assign n21601 =  ( n21564 ) ? ( VREG_1_2 ) : ( n21600 ) ;
assign n21602 =  ( n21563 ) ? ( VREG_1_3 ) : ( n21601 ) ;
assign n21603 =  ( n21562 ) ? ( VREG_1_4 ) : ( n21602 ) ;
assign n21604 =  ( n21561 ) ? ( VREG_1_5 ) : ( n21603 ) ;
assign n21605 =  ( n21560 ) ? ( VREG_1_6 ) : ( n21604 ) ;
assign n21606 =  ( n21559 ) ? ( VREG_1_7 ) : ( n21605 ) ;
assign n21607 =  ( n21558 ) ? ( VREG_1_8 ) : ( n21606 ) ;
assign n21608 =  ( n21557 ) ? ( VREG_1_9 ) : ( n21607 ) ;
assign n21609 =  ( n21556 ) ? ( VREG_1_10 ) : ( n21608 ) ;
assign n21610 =  ( n21555 ) ? ( VREG_1_11 ) : ( n21609 ) ;
assign n21611 =  ( n21554 ) ? ( VREG_1_12 ) : ( n21610 ) ;
assign n21612 =  ( n21553 ) ? ( VREG_1_13 ) : ( n21611 ) ;
assign n21613 =  ( n21552 ) ? ( VREG_1_14 ) : ( n21612 ) ;
assign n21614 =  ( n21551 ) ? ( VREG_1_15 ) : ( n21613 ) ;
assign n21615 =  ( n21550 ) ? ( VREG_2_0 ) : ( n21614 ) ;
assign n21616 =  ( n21549 ) ? ( VREG_2_1 ) : ( n21615 ) ;
assign n21617 =  ( n21548 ) ? ( VREG_2_2 ) : ( n21616 ) ;
assign n21618 =  ( n21547 ) ? ( VREG_2_3 ) : ( n21617 ) ;
assign n21619 =  ( n21546 ) ? ( VREG_2_4 ) : ( n21618 ) ;
assign n21620 =  ( n21545 ) ? ( VREG_2_5 ) : ( n21619 ) ;
assign n21621 =  ( n21544 ) ? ( VREG_2_6 ) : ( n21620 ) ;
assign n21622 =  ( n21543 ) ? ( VREG_2_7 ) : ( n21621 ) ;
assign n21623 =  ( n21542 ) ? ( VREG_2_8 ) : ( n21622 ) ;
assign n21624 =  ( n21541 ) ? ( VREG_2_9 ) : ( n21623 ) ;
assign n21625 =  ( n21540 ) ? ( VREG_2_10 ) : ( n21624 ) ;
assign n21626 =  ( n21539 ) ? ( VREG_2_11 ) : ( n21625 ) ;
assign n21627 =  ( n21538 ) ? ( VREG_2_12 ) : ( n21626 ) ;
assign n21628 =  ( n21537 ) ? ( VREG_2_13 ) : ( n21627 ) ;
assign n21629 =  ( n21536 ) ? ( VREG_2_14 ) : ( n21628 ) ;
assign n21630 =  ( n21535 ) ? ( VREG_2_15 ) : ( n21629 ) ;
assign n21631 =  ( n21534 ) ? ( VREG_3_0 ) : ( n21630 ) ;
assign n21632 =  ( n21533 ) ? ( VREG_3_1 ) : ( n21631 ) ;
assign n21633 =  ( n21532 ) ? ( VREG_3_2 ) : ( n21632 ) ;
assign n21634 =  ( n21531 ) ? ( VREG_3_3 ) : ( n21633 ) ;
assign n21635 =  ( n21530 ) ? ( VREG_3_4 ) : ( n21634 ) ;
assign n21636 =  ( n21529 ) ? ( VREG_3_5 ) : ( n21635 ) ;
assign n21637 =  ( n21528 ) ? ( VREG_3_6 ) : ( n21636 ) ;
assign n21638 =  ( n21527 ) ? ( VREG_3_7 ) : ( n21637 ) ;
assign n21639 =  ( n21526 ) ? ( VREG_3_8 ) : ( n21638 ) ;
assign n21640 =  ( n21525 ) ? ( VREG_3_9 ) : ( n21639 ) ;
assign n21641 =  ( n21524 ) ? ( VREG_3_10 ) : ( n21640 ) ;
assign n21642 =  ( n21523 ) ? ( VREG_3_11 ) : ( n21641 ) ;
assign n21643 =  ( n21522 ) ? ( VREG_3_12 ) : ( n21642 ) ;
assign n21644 =  ( n21521 ) ? ( VREG_3_13 ) : ( n21643 ) ;
assign n21645 =  ( n21520 ) ? ( VREG_3_14 ) : ( n21644 ) ;
assign n21646 =  ( n21519 ) ? ( VREG_3_15 ) : ( n21645 ) ;
assign n21647 =  ( n21518 ) ? ( VREG_4_0 ) : ( n21646 ) ;
assign n21648 =  ( n21517 ) ? ( VREG_4_1 ) : ( n21647 ) ;
assign n21649 =  ( n21516 ) ? ( VREG_4_2 ) : ( n21648 ) ;
assign n21650 =  ( n21515 ) ? ( VREG_4_3 ) : ( n21649 ) ;
assign n21651 =  ( n21514 ) ? ( VREG_4_4 ) : ( n21650 ) ;
assign n21652 =  ( n21513 ) ? ( VREG_4_5 ) : ( n21651 ) ;
assign n21653 =  ( n21512 ) ? ( VREG_4_6 ) : ( n21652 ) ;
assign n21654 =  ( n21511 ) ? ( VREG_4_7 ) : ( n21653 ) ;
assign n21655 =  ( n21510 ) ? ( VREG_4_8 ) : ( n21654 ) ;
assign n21656 =  ( n21509 ) ? ( VREG_4_9 ) : ( n21655 ) ;
assign n21657 =  ( n21508 ) ? ( VREG_4_10 ) : ( n21656 ) ;
assign n21658 =  ( n21507 ) ? ( VREG_4_11 ) : ( n21657 ) ;
assign n21659 =  ( n21506 ) ? ( VREG_4_12 ) : ( n21658 ) ;
assign n21660 =  ( n21505 ) ? ( VREG_4_13 ) : ( n21659 ) ;
assign n21661 =  ( n21504 ) ? ( VREG_4_14 ) : ( n21660 ) ;
assign n21662 =  ( n21503 ) ? ( VREG_4_15 ) : ( n21661 ) ;
assign n21663 =  ( n21502 ) ? ( VREG_5_0 ) : ( n21662 ) ;
assign n21664 =  ( n21501 ) ? ( VREG_5_1 ) : ( n21663 ) ;
assign n21665 =  ( n21500 ) ? ( VREG_5_2 ) : ( n21664 ) ;
assign n21666 =  ( n21499 ) ? ( VREG_5_3 ) : ( n21665 ) ;
assign n21667 =  ( n21498 ) ? ( VREG_5_4 ) : ( n21666 ) ;
assign n21668 =  ( n21497 ) ? ( VREG_5_5 ) : ( n21667 ) ;
assign n21669 =  ( n21496 ) ? ( VREG_5_6 ) : ( n21668 ) ;
assign n21670 =  ( n21495 ) ? ( VREG_5_7 ) : ( n21669 ) ;
assign n21671 =  ( n21494 ) ? ( VREG_5_8 ) : ( n21670 ) ;
assign n21672 =  ( n21493 ) ? ( VREG_5_9 ) : ( n21671 ) ;
assign n21673 =  ( n21492 ) ? ( VREG_5_10 ) : ( n21672 ) ;
assign n21674 =  ( n21491 ) ? ( VREG_5_11 ) : ( n21673 ) ;
assign n21675 =  ( n21490 ) ? ( VREG_5_12 ) : ( n21674 ) ;
assign n21676 =  ( n21489 ) ? ( VREG_5_13 ) : ( n21675 ) ;
assign n21677 =  ( n21488 ) ? ( VREG_5_14 ) : ( n21676 ) ;
assign n21678 =  ( n21487 ) ? ( VREG_5_15 ) : ( n21677 ) ;
assign n21679 =  ( n21486 ) ? ( VREG_6_0 ) : ( n21678 ) ;
assign n21680 =  ( n21485 ) ? ( VREG_6_1 ) : ( n21679 ) ;
assign n21681 =  ( n21484 ) ? ( VREG_6_2 ) : ( n21680 ) ;
assign n21682 =  ( n21483 ) ? ( VREG_6_3 ) : ( n21681 ) ;
assign n21683 =  ( n21482 ) ? ( VREG_6_4 ) : ( n21682 ) ;
assign n21684 =  ( n21481 ) ? ( VREG_6_5 ) : ( n21683 ) ;
assign n21685 =  ( n21480 ) ? ( VREG_6_6 ) : ( n21684 ) ;
assign n21686 =  ( n21479 ) ? ( VREG_6_7 ) : ( n21685 ) ;
assign n21687 =  ( n21478 ) ? ( VREG_6_8 ) : ( n21686 ) ;
assign n21688 =  ( n21477 ) ? ( VREG_6_9 ) : ( n21687 ) ;
assign n21689 =  ( n21476 ) ? ( VREG_6_10 ) : ( n21688 ) ;
assign n21690 =  ( n21475 ) ? ( VREG_6_11 ) : ( n21689 ) ;
assign n21691 =  ( n21474 ) ? ( VREG_6_12 ) : ( n21690 ) ;
assign n21692 =  ( n21473 ) ? ( VREG_6_13 ) : ( n21691 ) ;
assign n21693 =  ( n21472 ) ? ( VREG_6_14 ) : ( n21692 ) ;
assign n21694 =  ( n21471 ) ? ( VREG_6_15 ) : ( n21693 ) ;
assign n21695 =  ( n21470 ) ? ( VREG_7_0 ) : ( n21694 ) ;
assign n21696 =  ( n21469 ) ? ( VREG_7_1 ) : ( n21695 ) ;
assign n21697 =  ( n21468 ) ? ( VREG_7_2 ) : ( n21696 ) ;
assign n21698 =  ( n21467 ) ? ( VREG_7_3 ) : ( n21697 ) ;
assign n21699 =  ( n21466 ) ? ( VREG_7_4 ) : ( n21698 ) ;
assign n21700 =  ( n21465 ) ? ( VREG_7_5 ) : ( n21699 ) ;
assign n21701 =  ( n21464 ) ? ( VREG_7_6 ) : ( n21700 ) ;
assign n21702 =  ( n21463 ) ? ( VREG_7_7 ) : ( n21701 ) ;
assign n21703 =  ( n21462 ) ? ( VREG_7_8 ) : ( n21702 ) ;
assign n21704 =  ( n21461 ) ? ( VREG_7_9 ) : ( n21703 ) ;
assign n21705 =  ( n21460 ) ? ( VREG_7_10 ) : ( n21704 ) ;
assign n21706 =  ( n21459 ) ? ( VREG_7_11 ) : ( n21705 ) ;
assign n21707 =  ( n21458 ) ? ( VREG_7_12 ) : ( n21706 ) ;
assign n21708 =  ( n21457 ) ? ( VREG_7_13 ) : ( n21707 ) ;
assign n21709 =  ( n21456 ) ? ( VREG_7_14 ) : ( n21708 ) ;
assign n21710 =  ( n21455 ) ? ( VREG_7_15 ) : ( n21709 ) ;
assign n21711 =  ( n21454 ) ? ( VREG_8_0 ) : ( n21710 ) ;
assign n21712 =  ( n21453 ) ? ( VREG_8_1 ) : ( n21711 ) ;
assign n21713 =  ( n21452 ) ? ( VREG_8_2 ) : ( n21712 ) ;
assign n21714 =  ( n21451 ) ? ( VREG_8_3 ) : ( n21713 ) ;
assign n21715 =  ( n21450 ) ? ( VREG_8_4 ) : ( n21714 ) ;
assign n21716 =  ( n21449 ) ? ( VREG_8_5 ) : ( n21715 ) ;
assign n21717 =  ( n21448 ) ? ( VREG_8_6 ) : ( n21716 ) ;
assign n21718 =  ( n21447 ) ? ( VREG_8_7 ) : ( n21717 ) ;
assign n21719 =  ( n21446 ) ? ( VREG_8_8 ) : ( n21718 ) ;
assign n21720 =  ( n21445 ) ? ( VREG_8_9 ) : ( n21719 ) ;
assign n21721 =  ( n21444 ) ? ( VREG_8_10 ) : ( n21720 ) ;
assign n21722 =  ( n21443 ) ? ( VREG_8_11 ) : ( n21721 ) ;
assign n21723 =  ( n21442 ) ? ( VREG_8_12 ) : ( n21722 ) ;
assign n21724 =  ( n21441 ) ? ( VREG_8_13 ) : ( n21723 ) ;
assign n21725 =  ( n21440 ) ? ( VREG_8_14 ) : ( n21724 ) ;
assign n21726 =  ( n21439 ) ? ( VREG_8_15 ) : ( n21725 ) ;
assign n21727 =  ( n21438 ) ? ( VREG_9_0 ) : ( n21726 ) ;
assign n21728 =  ( n21437 ) ? ( VREG_9_1 ) : ( n21727 ) ;
assign n21729 =  ( n21436 ) ? ( VREG_9_2 ) : ( n21728 ) ;
assign n21730 =  ( n21435 ) ? ( VREG_9_3 ) : ( n21729 ) ;
assign n21731 =  ( n21434 ) ? ( VREG_9_4 ) : ( n21730 ) ;
assign n21732 =  ( n21433 ) ? ( VREG_9_5 ) : ( n21731 ) ;
assign n21733 =  ( n21432 ) ? ( VREG_9_6 ) : ( n21732 ) ;
assign n21734 =  ( n21431 ) ? ( VREG_9_7 ) : ( n21733 ) ;
assign n21735 =  ( n21430 ) ? ( VREG_9_8 ) : ( n21734 ) ;
assign n21736 =  ( n21429 ) ? ( VREG_9_9 ) : ( n21735 ) ;
assign n21737 =  ( n21428 ) ? ( VREG_9_10 ) : ( n21736 ) ;
assign n21738 =  ( n21427 ) ? ( VREG_9_11 ) : ( n21737 ) ;
assign n21739 =  ( n21426 ) ? ( VREG_9_12 ) : ( n21738 ) ;
assign n21740 =  ( n21425 ) ? ( VREG_9_13 ) : ( n21739 ) ;
assign n21741 =  ( n21424 ) ? ( VREG_9_14 ) : ( n21740 ) ;
assign n21742 =  ( n21423 ) ? ( VREG_9_15 ) : ( n21741 ) ;
assign n21743 =  ( n21422 ) ? ( VREG_10_0 ) : ( n21742 ) ;
assign n21744 =  ( n21421 ) ? ( VREG_10_1 ) : ( n21743 ) ;
assign n21745 =  ( n21420 ) ? ( VREG_10_2 ) : ( n21744 ) ;
assign n21746 =  ( n21419 ) ? ( VREG_10_3 ) : ( n21745 ) ;
assign n21747 =  ( n21418 ) ? ( VREG_10_4 ) : ( n21746 ) ;
assign n21748 =  ( n21417 ) ? ( VREG_10_5 ) : ( n21747 ) ;
assign n21749 =  ( n21416 ) ? ( VREG_10_6 ) : ( n21748 ) ;
assign n21750 =  ( n21415 ) ? ( VREG_10_7 ) : ( n21749 ) ;
assign n21751 =  ( n21414 ) ? ( VREG_10_8 ) : ( n21750 ) ;
assign n21752 =  ( n21413 ) ? ( VREG_10_9 ) : ( n21751 ) ;
assign n21753 =  ( n21412 ) ? ( VREG_10_10 ) : ( n21752 ) ;
assign n21754 =  ( n21411 ) ? ( VREG_10_11 ) : ( n21753 ) ;
assign n21755 =  ( n21410 ) ? ( VREG_10_12 ) : ( n21754 ) ;
assign n21756 =  ( n21409 ) ? ( VREG_10_13 ) : ( n21755 ) ;
assign n21757 =  ( n21408 ) ? ( VREG_10_14 ) : ( n21756 ) ;
assign n21758 =  ( n21407 ) ? ( VREG_10_15 ) : ( n21757 ) ;
assign n21759 =  ( n21406 ) ? ( VREG_11_0 ) : ( n21758 ) ;
assign n21760 =  ( n21405 ) ? ( VREG_11_1 ) : ( n21759 ) ;
assign n21761 =  ( n21404 ) ? ( VREG_11_2 ) : ( n21760 ) ;
assign n21762 =  ( n21403 ) ? ( VREG_11_3 ) : ( n21761 ) ;
assign n21763 =  ( n21402 ) ? ( VREG_11_4 ) : ( n21762 ) ;
assign n21764 =  ( n21401 ) ? ( VREG_11_5 ) : ( n21763 ) ;
assign n21765 =  ( n21400 ) ? ( VREG_11_6 ) : ( n21764 ) ;
assign n21766 =  ( n21399 ) ? ( VREG_11_7 ) : ( n21765 ) ;
assign n21767 =  ( n21398 ) ? ( VREG_11_8 ) : ( n21766 ) ;
assign n21768 =  ( n21397 ) ? ( VREG_11_9 ) : ( n21767 ) ;
assign n21769 =  ( n21396 ) ? ( VREG_11_10 ) : ( n21768 ) ;
assign n21770 =  ( n21395 ) ? ( VREG_11_11 ) : ( n21769 ) ;
assign n21771 =  ( n21394 ) ? ( VREG_11_12 ) : ( n21770 ) ;
assign n21772 =  ( n21393 ) ? ( VREG_11_13 ) : ( n21771 ) ;
assign n21773 =  ( n21392 ) ? ( VREG_11_14 ) : ( n21772 ) ;
assign n21774 =  ( n21391 ) ? ( VREG_11_15 ) : ( n21773 ) ;
assign n21775 =  ( n21390 ) ? ( VREG_12_0 ) : ( n21774 ) ;
assign n21776 =  ( n21389 ) ? ( VREG_12_1 ) : ( n21775 ) ;
assign n21777 =  ( n21388 ) ? ( VREG_12_2 ) : ( n21776 ) ;
assign n21778 =  ( n21387 ) ? ( VREG_12_3 ) : ( n21777 ) ;
assign n21779 =  ( n21386 ) ? ( VREG_12_4 ) : ( n21778 ) ;
assign n21780 =  ( n21385 ) ? ( VREG_12_5 ) : ( n21779 ) ;
assign n21781 =  ( n21384 ) ? ( VREG_12_6 ) : ( n21780 ) ;
assign n21782 =  ( n21383 ) ? ( VREG_12_7 ) : ( n21781 ) ;
assign n21783 =  ( n21382 ) ? ( VREG_12_8 ) : ( n21782 ) ;
assign n21784 =  ( n21381 ) ? ( VREG_12_9 ) : ( n21783 ) ;
assign n21785 =  ( n21380 ) ? ( VREG_12_10 ) : ( n21784 ) ;
assign n21786 =  ( n21379 ) ? ( VREG_12_11 ) : ( n21785 ) ;
assign n21787 =  ( n21378 ) ? ( VREG_12_12 ) : ( n21786 ) ;
assign n21788 =  ( n21377 ) ? ( VREG_12_13 ) : ( n21787 ) ;
assign n21789 =  ( n21376 ) ? ( VREG_12_14 ) : ( n21788 ) ;
assign n21790 =  ( n21375 ) ? ( VREG_12_15 ) : ( n21789 ) ;
assign n21791 =  ( n21374 ) ? ( VREG_13_0 ) : ( n21790 ) ;
assign n21792 =  ( n21373 ) ? ( VREG_13_1 ) : ( n21791 ) ;
assign n21793 =  ( n21372 ) ? ( VREG_13_2 ) : ( n21792 ) ;
assign n21794 =  ( n21371 ) ? ( VREG_13_3 ) : ( n21793 ) ;
assign n21795 =  ( n21370 ) ? ( VREG_13_4 ) : ( n21794 ) ;
assign n21796 =  ( n21369 ) ? ( VREG_13_5 ) : ( n21795 ) ;
assign n21797 =  ( n21368 ) ? ( VREG_13_6 ) : ( n21796 ) ;
assign n21798 =  ( n21367 ) ? ( VREG_13_7 ) : ( n21797 ) ;
assign n21799 =  ( n21366 ) ? ( VREG_13_8 ) : ( n21798 ) ;
assign n21800 =  ( n21365 ) ? ( VREG_13_9 ) : ( n21799 ) ;
assign n21801 =  ( n21364 ) ? ( VREG_13_10 ) : ( n21800 ) ;
assign n21802 =  ( n21363 ) ? ( VREG_13_11 ) : ( n21801 ) ;
assign n21803 =  ( n21362 ) ? ( VREG_13_12 ) : ( n21802 ) ;
assign n21804 =  ( n21361 ) ? ( VREG_13_13 ) : ( n21803 ) ;
assign n21805 =  ( n21360 ) ? ( VREG_13_14 ) : ( n21804 ) ;
assign n21806 =  ( n21359 ) ? ( VREG_13_15 ) : ( n21805 ) ;
assign n21807 =  ( n21358 ) ? ( VREG_14_0 ) : ( n21806 ) ;
assign n21808 =  ( n21357 ) ? ( VREG_14_1 ) : ( n21807 ) ;
assign n21809 =  ( n21356 ) ? ( VREG_14_2 ) : ( n21808 ) ;
assign n21810 =  ( n21355 ) ? ( VREG_14_3 ) : ( n21809 ) ;
assign n21811 =  ( n21354 ) ? ( VREG_14_4 ) : ( n21810 ) ;
assign n21812 =  ( n21353 ) ? ( VREG_14_5 ) : ( n21811 ) ;
assign n21813 =  ( n21352 ) ? ( VREG_14_6 ) : ( n21812 ) ;
assign n21814 =  ( n21351 ) ? ( VREG_14_7 ) : ( n21813 ) ;
assign n21815 =  ( n21350 ) ? ( VREG_14_8 ) : ( n21814 ) ;
assign n21816 =  ( n21349 ) ? ( VREG_14_9 ) : ( n21815 ) ;
assign n21817 =  ( n21348 ) ? ( VREG_14_10 ) : ( n21816 ) ;
assign n21818 =  ( n21347 ) ? ( VREG_14_11 ) : ( n21817 ) ;
assign n21819 =  ( n21346 ) ? ( VREG_14_12 ) : ( n21818 ) ;
assign n21820 =  ( n21345 ) ? ( VREG_14_13 ) : ( n21819 ) ;
assign n21821 =  ( n21344 ) ? ( VREG_14_14 ) : ( n21820 ) ;
assign n21822 =  ( n21343 ) ? ( VREG_14_15 ) : ( n21821 ) ;
assign n21823 =  ( n21342 ) ? ( VREG_15_0 ) : ( n21822 ) ;
assign n21824 =  ( n21341 ) ? ( VREG_15_1 ) : ( n21823 ) ;
assign n21825 =  ( n21340 ) ? ( VREG_15_2 ) : ( n21824 ) ;
assign n21826 =  ( n21339 ) ? ( VREG_15_3 ) : ( n21825 ) ;
assign n21827 =  ( n21338 ) ? ( VREG_15_4 ) : ( n21826 ) ;
assign n21828 =  ( n21337 ) ? ( VREG_15_5 ) : ( n21827 ) ;
assign n21829 =  ( n21336 ) ? ( VREG_15_6 ) : ( n21828 ) ;
assign n21830 =  ( n21335 ) ? ( VREG_15_7 ) : ( n21829 ) ;
assign n21831 =  ( n21334 ) ? ( VREG_15_8 ) : ( n21830 ) ;
assign n21832 =  ( n21333 ) ? ( VREG_15_9 ) : ( n21831 ) ;
assign n21833 =  ( n21332 ) ? ( VREG_15_10 ) : ( n21832 ) ;
assign n21834 =  ( n21331 ) ? ( VREG_15_11 ) : ( n21833 ) ;
assign n21835 =  ( n21330 ) ? ( VREG_15_12 ) : ( n21834 ) ;
assign n21836 =  ( n21329 ) ? ( VREG_15_13 ) : ( n21835 ) ;
assign n21837 =  ( n21328 ) ? ( VREG_15_14 ) : ( n21836 ) ;
assign n21838 =  ( n21327 ) ? ( VREG_15_15 ) : ( n21837 ) ;
assign n21839 =  ( n21326 ) ? ( VREG_16_0 ) : ( n21838 ) ;
assign n21840 =  ( n21325 ) ? ( VREG_16_1 ) : ( n21839 ) ;
assign n21841 =  ( n21324 ) ? ( VREG_16_2 ) : ( n21840 ) ;
assign n21842 =  ( n21323 ) ? ( VREG_16_3 ) : ( n21841 ) ;
assign n21843 =  ( n21322 ) ? ( VREG_16_4 ) : ( n21842 ) ;
assign n21844 =  ( n21321 ) ? ( VREG_16_5 ) : ( n21843 ) ;
assign n21845 =  ( n21320 ) ? ( VREG_16_6 ) : ( n21844 ) ;
assign n21846 =  ( n21319 ) ? ( VREG_16_7 ) : ( n21845 ) ;
assign n21847 =  ( n21318 ) ? ( VREG_16_8 ) : ( n21846 ) ;
assign n21848 =  ( n21317 ) ? ( VREG_16_9 ) : ( n21847 ) ;
assign n21849 =  ( n21316 ) ? ( VREG_16_10 ) : ( n21848 ) ;
assign n21850 =  ( n21315 ) ? ( VREG_16_11 ) : ( n21849 ) ;
assign n21851 =  ( n21314 ) ? ( VREG_16_12 ) : ( n21850 ) ;
assign n21852 =  ( n21313 ) ? ( VREG_16_13 ) : ( n21851 ) ;
assign n21853 =  ( n21312 ) ? ( VREG_16_14 ) : ( n21852 ) ;
assign n21854 =  ( n21311 ) ? ( VREG_16_15 ) : ( n21853 ) ;
assign n21855 =  ( n21310 ) ? ( VREG_17_0 ) : ( n21854 ) ;
assign n21856 =  ( n21309 ) ? ( VREG_17_1 ) : ( n21855 ) ;
assign n21857 =  ( n21308 ) ? ( VREG_17_2 ) : ( n21856 ) ;
assign n21858 =  ( n21307 ) ? ( VREG_17_3 ) : ( n21857 ) ;
assign n21859 =  ( n21306 ) ? ( VREG_17_4 ) : ( n21858 ) ;
assign n21860 =  ( n21305 ) ? ( VREG_17_5 ) : ( n21859 ) ;
assign n21861 =  ( n21304 ) ? ( VREG_17_6 ) : ( n21860 ) ;
assign n21862 =  ( n21303 ) ? ( VREG_17_7 ) : ( n21861 ) ;
assign n21863 =  ( n21302 ) ? ( VREG_17_8 ) : ( n21862 ) ;
assign n21864 =  ( n21301 ) ? ( VREG_17_9 ) : ( n21863 ) ;
assign n21865 =  ( n21300 ) ? ( VREG_17_10 ) : ( n21864 ) ;
assign n21866 =  ( n21299 ) ? ( VREG_17_11 ) : ( n21865 ) ;
assign n21867 =  ( n21298 ) ? ( VREG_17_12 ) : ( n21866 ) ;
assign n21868 =  ( n21297 ) ? ( VREG_17_13 ) : ( n21867 ) ;
assign n21869 =  ( n21296 ) ? ( VREG_17_14 ) : ( n21868 ) ;
assign n21870 =  ( n21295 ) ? ( VREG_17_15 ) : ( n21869 ) ;
assign n21871 =  ( n21294 ) ? ( VREG_18_0 ) : ( n21870 ) ;
assign n21872 =  ( n21293 ) ? ( VREG_18_1 ) : ( n21871 ) ;
assign n21873 =  ( n21292 ) ? ( VREG_18_2 ) : ( n21872 ) ;
assign n21874 =  ( n21291 ) ? ( VREG_18_3 ) : ( n21873 ) ;
assign n21875 =  ( n21290 ) ? ( VREG_18_4 ) : ( n21874 ) ;
assign n21876 =  ( n21289 ) ? ( VREG_18_5 ) : ( n21875 ) ;
assign n21877 =  ( n21288 ) ? ( VREG_18_6 ) : ( n21876 ) ;
assign n21878 =  ( n21287 ) ? ( VREG_18_7 ) : ( n21877 ) ;
assign n21879 =  ( n21286 ) ? ( VREG_18_8 ) : ( n21878 ) ;
assign n21880 =  ( n21285 ) ? ( VREG_18_9 ) : ( n21879 ) ;
assign n21881 =  ( n21284 ) ? ( VREG_18_10 ) : ( n21880 ) ;
assign n21882 =  ( n21283 ) ? ( VREG_18_11 ) : ( n21881 ) ;
assign n21883 =  ( n21282 ) ? ( VREG_18_12 ) : ( n21882 ) ;
assign n21884 =  ( n21281 ) ? ( VREG_18_13 ) : ( n21883 ) ;
assign n21885 =  ( n21280 ) ? ( VREG_18_14 ) : ( n21884 ) ;
assign n21886 =  ( n21279 ) ? ( VREG_18_15 ) : ( n21885 ) ;
assign n21887 =  ( n21278 ) ? ( VREG_19_0 ) : ( n21886 ) ;
assign n21888 =  ( n21277 ) ? ( VREG_19_1 ) : ( n21887 ) ;
assign n21889 =  ( n21276 ) ? ( VREG_19_2 ) : ( n21888 ) ;
assign n21890 =  ( n21275 ) ? ( VREG_19_3 ) : ( n21889 ) ;
assign n21891 =  ( n21274 ) ? ( VREG_19_4 ) : ( n21890 ) ;
assign n21892 =  ( n21273 ) ? ( VREG_19_5 ) : ( n21891 ) ;
assign n21893 =  ( n21272 ) ? ( VREG_19_6 ) : ( n21892 ) ;
assign n21894 =  ( n21271 ) ? ( VREG_19_7 ) : ( n21893 ) ;
assign n21895 =  ( n21270 ) ? ( VREG_19_8 ) : ( n21894 ) ;
assign n21896 =  ( n21269 ) ? ( VREG_19_9 ) : ( n21895 ) ;
assign n21897 =  ( n21268 ) ? ( VREG_19_10 ) : ( n21896 ) ;
assign n21898 =  ( n21267 ) ? ( VREG_19_11 ) : ( n21897 ) ;
assign n21899 =  ( n21266 ) ? ( VREG_19_12 ) : ( n21898 ) ;
assign n21900 =  ( n21265 ) ? ( VREG_19_13 ) : ( n21899 ) ;
assign n21901 =  ( n21264 ) ? ( VREG_19_14 ) : ( n21900 ) ;
assign n21902 =  ( n21263 ) ? ( VREG_19_15 ) : ( n21901 ) ;
assign n21903 =  ( n21262 ) ? ( VREG_20_0 ) : ( n21902 ) ;
assign n21904 =  ( n21261 ) ? ( VREG_20_1 ) : ( n21903 ) ;
assign n21905 =  ( n21260 ) ? ( VREG_20_2 ) : ( n21904 ) ;
assign n21906 =  ( n21259 ) ? ( VREG_20_3 ) : ( n21905 ) ;
assign n21907 =  ( n21258 ) ? ( VREG_20_4 ) : ( n21906 ) ;
assign n21908 =  ( n21257 ) ? ( VREG_20_5 ) : ( n21907 ) ;
assign n21909 =  ( n21256 ) ? ( VREG_20_6 ) : ( n21908 ) ;
assign n21910 =  ( n21255 ) ? ( VREG_20_7 ) : ( n21909 ) ;
assign n21911 =  ( n21254 ) ? ( VREG_20_8 ) : ( n21910 ) ;
assign n21912 =  ( n21253 ) ? ( VREG_20_9 ) : ( n21911 ) ;
assign n21913 =  ( n21252 ) ? ( VREG_20_10 ) : ( n21912 ) ;
assign n21914 =  ( n21251 ) ? ( VREG_20_11 ) : ( n21913 ) ;
assign n21915 =  ( n21250 ) ? ( VREG_20_12 ) : ( n21914 ) ;
assign n21916 =  ( n21249 ) ? ( VREG_20_13 ) : ( n21915 ) ;
assign n21917 =  ( n21248 ) ? ( VREG_20_14 ) : ( n21916 ) ;
assign n21918 =  ( n21247 ) ? ( VREG_20_15 ) : ( n21917 ) ;
assign n21919 =  ( n21246 ) ? ( VREG_21_0 ) : ( n21918 ) ;
assign n21920 =  ( n21245 ) ? ( VREG_21_1 ) : ( n21919 ) ;
assign n21921 =  ( n21244 ) ? ( VREG_21_2 ) : ( n21920 ) ;
assign n21922 =  ( n21243 ) ? ( VREG_21_3 ) : ( n21921 ) ;
assign n21923 =  ( n21242 ) ? ( VREG_21_4 ) : ( n21922 ) ;
assign n21924 =  ( n21241 ) ? ( VREG_21_5 ) : ( n21923 ) ;
assign n21925 =  ( n21240 ) ? ( VREG_21_6 ) : ( n21924 ) ;
assign n21926 =  ( n21239 ) ? ( VREG_21_7 ) : ( n21925 ) ;
assign n21927 =  ( n21238 ) ? ( VREG_21_8 ) : ( n21926 ) ;
assign n21928 =  ( n21237 ) ? ( VREG_21_9 ) : ( n21927 ) ;
assign n21929 =  ( n21236 ) ? ( VREG_21_10 ) : ( n21928 ) ;
assign n21930 =  ( n21235 ) ? ( VREG_21_11 ) : ( n21929 ) ;
assign n21931 =  ( n21234 ) ? ( VREG_21_12 ) : ( n21930 ) ;
assign n21932 =  ( n21233 ) ? ( VREG_21_13 ) : ( n21931 ) ;
assign n21933 =  ( n21232 ) ? ( VREG_21_14 ) : ( n21932 ) ;
assign n21934 =  ( n21231 ) ? ( VREG_21_15 ) : ( n21933 ) ;
assign n21935 =  ( n21230 ) ? ( VREG_22_0 ) : ( n21934 ) ;
assign n21936 =  ( n21229 ) ? ( VREG_22_1 ) : ( n21935 ) ;
assign n21937 =  ( n21228 ) ? ( VREG_22_2 ) : ( n21936 ) ;
assign n21938 =  ( n21227 ) ? ( VREG_22_3 ) : ( n21937 ) ;
assign n21939 =  ( n21226 ) ? ( VREG_22_4 ) : ( n21938 ) ;
assign n21940 =  ( n21225 ) ? ( VREG_22_5 ) : ( n21939 ) ;
assign n21941 =  ( n21224 ) ? ( VREG_22_6 ) : ( n21940 ) ;
assign n21942 =  ( n21223 ) ? ( VREG_22_7 ) : ( n21941 ) ;
assign n21943 =  ( n21222 ) ? ( VREG_22_8 ) : ( n21942 ) ;
assign n21944 =  ( n21221 ) ? ( VREG_22_9 ) : ( n21943 ) ;
assign n21945 =  ( n21220 ) ? ( VREG_22_10 ) : ( n21944 ) ;
assign n21946 =  ( n21219 ) ? ( VREG_22_11 ) : ( n21945 ) ;
assign n21947 =  ( n21218 ) ? ( VREG_22_12 ) : ( n21946 ) ;
assign n21948 =  ( n21217 ) ? ( VREG_22_13 ) : ( n21947 ) ;
assign n21949 =  ( n21216 ) ? ( VREG_22_14 ) : ( n21948 ) ;
assign n21950 =  ( n21215 ) ? ( VREG_22_15 ) : ( n21949 ) ;
assign n21951 =  ( n21214 ) ? ( VREG_23_0 ) : ( n21950 ) ;
assign n21952 =  ( n21213 ) ? ( VREG_23_1 ) : ( n21951 ) ;
assign n21953 =  ( n21212 ) ? ( VREG_23_2 ) : ( n21952 ) ;
assign n21954 =  ( n21211 ) ? ( VREG_23_3 ) : ( n21953 ) ;
assign n21955 =  ( n21210 ) ? ( VREG_23_4 ) : ( n21954 ) ;
assign n21956 =  ( n21209 ) ? ( VREG_23_5 ) : ( n21955 ) ;
assign n21957 =  ( n21208 ) ? ( VREG_23_6 ) : ( n21956 ) ;
assign n21958 =  ( n21207 ) ? ( VREG_23_7 ) : ( n21957 ) ;
assign n21959 =  ( n21206 ) ? ( VREG_23_8 ) : ( n21958 ) ;
assign n21960 =  ( n21205 ) ? ( VREG_23_9 ) : ( n21959 ) ;
assign n21961 =  ( n21204 ) ? ( VREG_23_10 ) : ( n21960 ) ;
assign n21962 =  ( n21203 ) ? ( VREG_23_11 ) : ( n21961 ) ;
assign n21963 =  ( n21202 ) ? ( VREG_23_12 ) : ( n21962 ) ;
assign n21964 =  ( n21201 ) ? ( VREG_23_13 ) : ( n21963 ) ;
assign n21965 =  ( n21200 ) ? ( VREG_23_14 ) : ( n21964 ) ;
assign n21966 =  ( n21199 ) ? ( VREG_23_15 ) : ( n21965 ) ;
assign n21967 =  ( n21198 ) ? ( VREG_24_0 ) : ( n21966 ) ;
assign n21968 =  ( n21197 ) ? ( VREG_24_1 ) : ( n21967 ) ;
assign n21969 =  ( n21196 ) ? ( VREG_24_2 ) : ( n21968 ) ;
assign n21970 =  ( n21195 ) ? ( VREG_24_3 ) : ( n21969 ) ;
assign n21971 =  ( n21194 ) ? ( VREG_24_4 ) : ( n21970 ) ;
assign n21972 =  ( n21193 ) ? ( VREG_24_5 ) : ( n21971 ) ;
assign n21973 =  ( n21192 ) ? ( VREG_24_6 ) : ( n21972 ) ;
assign n21974 =  ( n21191 ) ? ( VREG_24_7 ) : ( n21973 ) ;
assign n21975 =  ( n21190 ) ? ( VREG_24_8 ) : ( n21974 ) ;
assign n21976 =  ( n21189 ) ? ( VREG_24_9 ) : ( n21975 ) ;
assign n21977 =  ( n21188 ) ? ( VREG_24_10 ) : ( n21976 ) ;
assign n21978 =  ( n21187 ) ? ( VREG_24_11 ) : ( n21977 ) ;
assign n21979 =  ( n21186 ) ? ( VREG_24_12 ) : ( n21978 ) ;
assign n21980 =  ( n21185 ) ? ( VREG_24_13 ) : ( n21979 ) ;
assign n21981 =  ( n21184 ) ? ( VREG_24_14 ) : ( n21980 ) ;
assign n21982 =  ( n21183 ) ? ( VREG_24_15 ) : ( n21981 ) ;
assign n21983 =  ( n21182 ) ? ( VREG_25_0 ) : ( n21982 ) ;
assign n21984 =  ( n21181 ) ? ( VREG_25_1 ) : ( n21983 ) ;
assign n21985 =  ( n21180 ) ? ( VREG_25_2 ) : ( n21984 ) ;
assign n21986 =  ( n21179 ) ? ( VREG_25_3 ) : ( n21985 ) ;
assign n21987 =  ( n21178 ) ? ( VREG_25_4 ) : ( n21986 ) ;
assign n21988 =  ( n21177 ) ? ( VREG_25_5 ) : ( n21987 ) ;
assign n21989 =  ( n21176 ) ? ( VREG_25_6 ) : ( n21988 ) ;
assign n21990 =  ( n21175 ) ? ( VREG_25_7 ) : ( n21989 ) ;
assign n21991 =  ( n21174 ) ? ( VREG_25_8 ) : ( n21990 ) ;
assign n21992 =  ( n21173 ) ? ( VREG_25_9 ) : ( n21991 ) ;
assign n21993 =  ( n21172 ) ? ( VREG_25_10 ) : ( n21992 ) ;
assign n21994 =  ( n21171 ) ? ( VREG_25_11 ) : ( n21993 ) ;
assign n21995 =  ( n21170 ) ? ( VREG_25_12 ) : ( n21994 ) ;
assign n21996 =  ( n21169 ) ? ( VREG_25_13 ) : ( n21995 ) ;
assign n21997 =  ( n21168 ) ? ( VREG_25_14 ) : ( n21996 ) ;
assign n21998 =  ( n21167 ) ? ( VREG_25_15 ) : ( n21997 ) ;
assign n21999 =  ( n21166 ) ? ( VREG_26_0 ) : ( n21998 ) ;
assign n22000 =  ( n21165 ) ? ( VREG_26_1 ) : ( n21999 ) ;
assign n22001 =  ( n21164 ) ? ( VREG_26_2 ) : ( n22000 ) ;
assign n22002 =  ( n21163 ) ? ( VREG_26_3 ) : ( n22001 ) ;
assign n22003 =  ( n21162 ) ? ( VREG_26_4 ) : ( n22002 ) ;
assign n22004 =  ( n21161 ) ? ( VREG_26_5 ) : ( n22003 ) ;
assign n22005 =  ( n21160 ) ? ( VREG_26_6 ) : ( n22004 ) ;
assign n22006 =  ( n21159 ) ? ( VREG_26_7 ) : ( n22005 ) ;
assign n22007 =  ( n21158 ) ? ( VREG_26_8 ) : ( n22006 ) ;
assign n22008 =  ( n21157 ) ? ( VREG_26_9 ) : ( n22007 ) ;
assign n22009 =  ( n21156 ) ? ( VREG_26_10 ) : ( n22008 ) ;
assign n22010 =  ( n21155 ) ? ( VREG_26_11 ) : ( n22009 ) ;
assign n22011 =  ( n21154 ) ? ( VREG_26_12 ) : ( n22010 ) ;
assign n22012 =  ( n21153 ) ? ( VREG_26_13 ) : ( n22011 ) ;
assign n22013 =  ( n21152 ) ? ( VREG_26_14 ) : ( n22012 ) ;
assign n22014 =  ( n21151 ) ? ( VREG_26_15 ) : ( n22013 ) ;
assign n22015 =  ( n21150 ) ? ( VREG_27_0 ) : ( n22014 ) ;
assign n22016 =  ( n21149 ) ? ( VREG_27_1 ) : ( n22015 ) ;
assign n22017 =  ( n21148 ) ? ( VREG_27_2 ) : ( n22016 ) ;
assign n22018 =  ( n21147 ) ? ( VREG_27_3 ) : ( n22017 ) ;
assign n22019 =  ( n21146 ) ? ( VREG_27_4 ) : ( n22018 ) ;
assign n22020 =  ( n21145 ) ? ( VREG_27_5 ) : ( n22019 ) ;
assign n22021 =  ( n21144 ) ? ( VREG_27_6 ) : ( n22020 ) ;
assign n22022 =  ( n21143 ) ? ( VREG_27_7 ) : ( n22021 ) ;
assign n22023 =  ( n21142 ) ? ( VREG_27_8 ) : ( n22022 ) ;
assign n22024 =  ( n21141 ) ? ( VREG_27_9 ) : ( n22023 ) ;
assign n22025 =  ( n21140 ) ? ( VREG_27_10 ) : ( n22024 ) ;
assign n22026 =  ( n21139 ) ? ( VREG_27_11 ) : ( n22025 ) ;
assign n22027 =  ( n21138 ) ? ( VREG_27_12 ) : ( n22026 ) ;
assign n22028 =  ( n21137 ) ? ( VREG_27_13 ) : ( n22027 ) ;
assign n22029 =  ( n21136 ) ? ( VREG_27_14 ) : ( n22028 ) ;
assign n22030 =  ( n21135 ) ? ( VREG_27_15 ) : ( n22029 ) ;
assign n22031 =  ( n21134 ) ? ( VREG_28_0 ) : ( n22030 ) ;
assign n22032 =  ( n21133 ) ? ( VREG_28_1 ) : ( n22031 ) ;
assign n22033 =  ( n21132 ) ? ( VREG_28_2 ) : ( n22032 ) ;
assign n22034 =  ( n21131 ) ? ( VREG_28_3 ) : ( n22033 ) ;
assign n22035 =  ( n21130 ) ? ( VREG_28_4 ) : ( n22034 ) ;
assign n22036 =  ( n21129 ) ? ( VREG_28_5 ) : ( n22035 ) ;
assign n22037 =  ( n21128 ) ? ( VREG_28_6 ) : ( n22036 ) ;
assign n22038 =  ( n21127 ) ? ( VREG_28_7 ) : ( n22037 ) ;
assign n22039 =  ( n21126 ) ? ( VREG_28_8 ) : ( n22038 ) ;
assign n22040 =  ( n21125 ) ? ( VREG_28_9 ) : ( n22039 ) ;
assign n22041 =  ( n21124 ) ? ( VREG_28_10 ) : ( n22040 ) ;
assign n22042 =  ( n21123 ) ? ( VREG_28_11 ) : ( n22041 ) ;
assign n22043 =  ( n21122 ) ? ( VREG_28_12 ) : ( n22042 ) ;
assign n22044 =  ( n21121 ) ? ( VREG_28_13 ) : ( n22043 ) ;
assign n22045 =  ( n21120 ) ? ( VREG_28_14 ) : ( n22044 ) ;
assign n22046 =  ( n21119 ) ? ( VREG_28_15 ) : ( n22045 ) ;
assign n22047 =  ( n21118 ) ? ( VREG_29_0 ) : ( n22046 ) ;
assign n22048 =  ( n21117 ) ? ( VREG_29_1 ) : ( n22047 ) ;
assign n22049 =  ( n21116 ) ? ( VREG_29_2 ) : ( n22048 ) ;
assign n22050 =  ( n21115 ) ? ( VREG_29_3 ) : ( n22049 ) ;
assign n22051 =  ( n21114 ) ? ( VREG_29_4 ) : ( n22050 ) ;
assign n22052 =  ( n21113 ) ? ( VREG_29_5 ) : ( n22051 ) ;
assign n22053 =  ( n21112 ) ? ( VREG_29_6 ) : ( n22052 ) ;
assign n22054 =  ( n21111 ) ? ( VREG_29_7 ) : ( n22053 ) ;
assign n22055 =  ( n21110 ) ? ( VREG_29_8 ) : ( n22054 ) ;
assign n22056 =  ( n21109 ) ? ( VREG_29_9 ) : ( n22055 ) ;
assign n22057 =  ( n21108 ) ? ( VREG_29_10 ) : ( n22056 ) ;
assign n22058 =  ( n21107 ) ? ( VREG_29_11 ) : ( n22057 ) ;
assign n22059 =  ( n21106 ) ? ( VREG_29_12 ) : ( n22058 ) ;
assign n22060 =  ( n21105 ) ? ( VREG_29_13 ) : ( n22059 ) ;
assign n22061 =  ( n21104 ) ? ( VREG_29_14 ) : ( n22060 ) ;
assign n22062 =  ( n21103 ) ? ( VREG_29_15 ) : ( n22061 ) ;
assign n22063 =  ( n21102 ) ? ( VREG_30_0 ) : ( n22062 ) ;
assign n22064 =  ( n21101 ) ? ( VREG_30_1 ) : ( n22063 ) ;
assign n22065 =  ( n21100 ) ? ( VREG_30_2 ) : ( n22064 ) ;
assign n22066 =  ( n21099 ) ? ( VREG_30_3 ) : ( n22065 ) ;
assign n22067 =  ( n21098 ) ? ( VREG_30_4 ) : ( n22066 ) ;
assign n22068 =  ( n21097 ) ? ( VREG_30_5 ) : ( n22067 ) ;
assign n22069 =  ( n21096 ) ? ( VREG_30_6 ) : ( n22068 ) ;
assign n22070 =  ( n21095 ) ? ( VREG_30_7 ) : ( n22069 ) ;
assign n22071 =  ( n21094 ) ? ( VREG_30_8 ) : ( n22070 ) ;
assign n22072 =  ( n21093 ) ? ( VREG_30_9 ) : ( n22071 ) ;
assign n22073 =  ( n21092 ) ? ( VREG_30_10 ) : ( n22072 ) ;
assign n22074 =  ( n21091 ) ? ( VREG_30_11 ) : ( n22073 ) ;
assign n22075 =  ( n21090 ) ? ( VREG_30_12 ) : ( n22074 ) ;
assign n22076 =  ( n21089 ) ? ( VREG_30_13 ) : ( n22075 ) ;
assign n22077 =  ( n21088 ) ? ( VREG_30_14 ) : ( n22076 ) ;
assign n22078 =  ( n21087 ) ? ( VREG_30_15 ) : ( n22077 ) ;
assign n22079 =  ( n21086 ) ? ( VREG_31_0 ) : ( n22078 ) ;
assign n22080 =  ( n21085 ) ? ( VREG_31_1 ) : ( n22079 ) ;
assign n22081 =  ( n21084 ) ? ( VREG_31_2 ) : ( n22080 ) ;
assign n22082 =  ( n21083 ) ? ( VREG_31_3 ) : ( n22081 ) ;
assign n22083 =  ( n21082 ) ? ( VREG_31_4 ) : ( n22082 ) ;
assign n22084 =  ( n21081 ) ? ( VREG_31_5 ) : ( n22083 ) ;
assign n22085 =  ( n21080 ) ? ( VREG_31_6 ) : ( n22084 ) ;
assign n22086 =  ( n21079 ) ? ( VREG_31_7 ) : ( n22085 ) ;
assign n22087 =  ( n21078 ) ? ( VREG_31_8 ) : ( n22086 ) ;
assign n22088 =  ( n21077 ) ? ( VREG_31_9 ) : ( n22087 ) ;
assign n22089 =  ( n21076 ) ? ( VREG_31_10 ) : ( n22088 ) ;
assign n22090 =  ( n21075 ) ? ( VREG_31_11 ) : ( n22089 ) ;
assign n22091 =  ( n21074 ) ? ( VREG_31_12 ) : ( n22090 ) ;
assign n22092 =  ( n21073 ) ? ( VREG_31_13 ) : ( n22091 ) ;
assign n22093 =  ( n21072 ) ? ( VREG_31_14 ) : ( n22092 ) ;
assign n22094 =  ( n21071 ) ? ( VREG_31_15 ) : ( n22093 ) ;
assign n22095 =  ( n21060 ) + ( n22094 )  ;
assign n22096 =  ( n21060 ) - ( n22094 )  ;
assign n22097 =  ( n21060 ) & ( n22094 )  ;
assign n22098 =  ( n21060 ) | ( n22094 )  ;
assign n22099 =  ( ( n21060 ) * ( n22094 ))  ;
assign n22100 =  ( n148 ) ? ( n22099 ) : ( VREG_0_3 ) ;
assign n22101 =  ( n146 ) ? ( n22098 ) : ( n22100 ) ;
assign n22102 =  ( n144 ) ? ( n22097 ) : ( n22101 ) ;
assign n22103 =  ( n142 ) ? ( n22096 ) : ( n22102 ) ;
assign n22104 =  ( n10 ) ? ( n22095 ) : ( n22103 ) ;
assign n22105 = n3030[3:3] ;
assign n22106 =  ( n22105 ) == ( 1'd0 )  ;
assign n22107 =  ( n22106 ) ? ( VREG_0_3 ) : ( n21070 ) ;
assign n22108 =  ( n22106 ) ? ( VREG_0_3 ) : ( n22104 ) ;
assign n22109 =  ( n3034 ) ? ( n22108 ) : ( VREG_0_3 ) ;
assign n22110 =  ( n2965 ) ? ( n22107 ) : ( n22109 ) ;
assign n22111 =  ( n1930 ) ? ( n22104 ) : ( n22110 ) ;
assign n22112 =  ( n879 ) ? ( n21070 ) : ( n22111 ) ;
assign n22113 =  ( n21060 ) + ( n164 )  ;
assign n22114 =  ( n21060 ) - ( n164 )  ;
assign n22115 =  ( n21060 ) & ( n164 )  ;
assign n22116 =  ( n21060 ) | ( n164 )  ;
assign n22117 =  ( ( n21060 ) * ( n164 ))  ;
assign n22118 =  ( n172 ) ? ( n22117 ) : ( VREG_0_3 ) ;
assign n22119 =  ( n170 ) ? ( n22116 ) : ( n22118 ) ;
assign n22120 =  ( n168 ) ? ( n22115 ) : ( n22119 ) ;
assign n22121 =  ( n166 ) ? ( n22114 ) : ( n22120 ) ;
assign n22122 =  ( n162 ) ? ( n22113 ) : ( n22121 ) ;
assign n22123 =  ( n21060 ) + ( n180 )  ;
assign n22124 =  ( n21060 ) - ( n180 )  ;
assign n22125 =  ( n21060 ) & ( n180 )  ;
assign n22126 =  ( n21060 ) | ( n180 )  ;
assign n22127 =  ( ( n21060 ) * ( n180 ))  ;
assign n22128 =  ( n172 ) ? ( n22127 ) : ( VREG_0_3 ) ;
assign n22129 =  ( n170 ) ? ( n22126 ) : ( n22128 ) ;
assign n22130 =  ( n168 ) ? ( n22125 ) : ( n22129 ) ;
assign n22131 =  ( n166 ) ? ( n22124 ) : ( n22130 ) ;
assign n22132 =  ( n162 ) ? ( n22123 ) : ( n22131 ) ;
assign n22133 =  ( n22106 ) ? ( VREG_0_3 ) : ( n22132 ) ;
assign n22134 =  ( n3051 ) ? ( n22133 ) : ( VREG_0_3 ) ;
assign n22135 =  ( n3040 ) ? ( n22122 ) : ( n22134 ) ;
assign n22136 =  ( n192 ) ? ( VREG_0_3 ) : ( VREG_0_3 ) ;
assign n22137 =  ( n157 ) ? ( n22135 ) : ( n22136 ) ;
assign n22138 =  ( n6 ) ? ( n22112 ) : ( n22137 ) ;
assign n22139 =  ( n4 ) ? ( n22138 ) : ( VREG_0_3 ) ;
assign n22140 =  ( 32'd4 ) == ( 32'd15 )  ;
assign n22141 =  ( n12 ) & ( n22140 )  ;
assign n22142 =  ( 32'd4 ) == ( 32'd14 )  ;
assign n22143 =  ( n12 ) & ( n22142 )  ;
assign n22144 =  ( 32'd4 ) == ( 32'd13 )  ;
assign n22145 =  ( n12 ) & ( n22144 )  ;
assign n22146 =  ( 32'd4 ) == ( 32'd12 )  ;
assign n22147 =  ( n12 ) & ( n22146 )  ;
assign n22148 =  ( 32'd4 ) == ( 32'd11 )  ;
assign n22149 =  ( n12 ) & ( n22148 )  ;
assign n22150 =  ( 32'd4 ) == ( 32'd10 )  ;
assign n22151 =  ( n12 ) & ( n22150 )  ;
assign n22152 =  ( 32'd4 ) == ( 32'd9 )  ;
assign n22153 =  ( n12 ) & ( n22152 )  ;
assign n22154 =  ( 32'd4 ) == ( 32'd8 )  ;
assign n22155 =  ( n12 ) & ( n22154 )  ;
assign n22156 =  ( 32'd4 ) == ( 32'd7 )  ;
assign n22157 =  ( n12 ) & ( n22156 )  ;
assign n22158 =  ( 32'd4 ) == ( 32'd6 )  ;
assign n22159 =  ( n12 ) & ( n22158 )  ;
assign n22160 =  ( 32'd4 ) == ( 32'd5 )  ;
assign n22161 =  ( n12 ) & ( n22160 )  ;
assign n22162 =  ( 32'd4 ) == ( 32'd4 )  ;
assign n22163 =  ( n12 ) & ( n22162 )  ;
assign n22164 =  ( 32'd4 ) == ( 32'd3 )  ;
assign n22165 =  ( n12 ) & ( n22164 )  ;
assign n22166 =  ( 32'd4 ) == ( 32'd2 )  ;
assign n22167 =  ( n12 ) & ( n22166 )  ;
assign n22168 =  ( 32'd4 ) == ( 32'd1 )  ;
assign n22169 =  ( n12 ) & ( n22168 )  ;
assign n22170 =  ( 32'd4 ) == ( 32'd0 )  ;
assign n22171 =  ( n12 ) & ( n22170 )  ;
assign n22172 =  ( n13 ) & ( n22140 )  ;
assign n22173 =  ( n13 ) & ( n22142 )  ;
assign n22174 =  ( n13 ) & ( n22144 )  ;
assign n22175 =  ( n13 ) & ( n22146 )  ;
assign n22176 =  ( n13 ) & ( n22148 )  ;
assign n22177 =  ( n13 ) & ( n22150 )  ;
assign n22178 =  ( n13 ) & ( n22152 )  ;
assign n22179 =  ( n13 ) & ( n22154 )  ;
assign n22180 =  ( n13 ) & ( n22156 )  ;
assign n22181 =  ( n13 ) & ( n22158 )  ;
assign n22182 =  ( n13 ) & ( n22160 )  ;
assign n22183 =  ( n13 ) & ( n22162 )  ;
assign n22184 =  ( n13 ) & ( n22164 )  ;
assign n22185 =  ( n13 ) & ( n22166 )  ;
assign n22186 =  ( n13 ) & ( n22168 )  ;
assign n22187 =  ( n13 ) & ( n22170 )  ;
assign n22188 =  ( n14 ) & ( n22140 )  ;
assign n22189 =  ( n14 ) & ( n22142 )  ;
assign n22190 =  ( n14 ) & ( n22144 )  ;
assign n22191 =  ( n14 ) & ( n22146 )  ;
assign n22192 =  ( n14 ) & ( n22148 )  ;
assign n22193 =  ( n14 ) & ( n22150 )  ;
assign n22194 =  ( n14 ) & ( n22152 )  ;
assign n22195 =  ( n14 ) & ( n22154 )  ;
assign n22196 =  ( n14 ) & ( n22156 )  ;
assign n22197 =  ( n14 ) & ( n22158 )  ;
assign n22198 =  ( n14 ) & ( n22160 )  ;
assign n22199 =  ( n14 ) & ( n22162 )  ;
assign n22200 =  ( n14 ) & ( n22164 )  ;
assign n22201 =  ( n14 ) & ( n22166 )  ;
assign n22202 =  ( n14 ) & ( n22168 )  ;
assign n22203 =  ( n14 ) & ( n22170 )  ;
assign n22204 =  ( n15 ) & ( n22140 )  ;
assign n22205 =  ( n15 ) & ( n22142 )  ;
assign n22206 =  ( n15 ) & ( n22144 )  ;
assign n22207 =  ( n15 ) & ( n22146 )  ;
assign n22208 =  ( n15 ) & ( n22148 )  ;
assign n22209 =  ( n15 ) & ( n22150 )  ;
assign n22210 =  ( n15 ) & ( n22152 )  ;
assign n22211 =  ( n15 ) & ( n22154 )  ;
assign n22212 =  ( n15 ) & ( n22156 )  ;
assign n22213 =  ( n15 ) & ( n22158 )  ;
assign n22214 =  ( n15 ) & ( n22160 )  ;
assign n22215 =  ( n15 ) & ( n22162 )  ;
assign n22216 =  ( n15 ) & ( n22164 )  ;
assign n22217 =  ( n15 ) & ( n22166 )  ;
assign n22218 =  ( n15 ) & ( n22168 )  ;
assign n22219 =  ( n15 ) & ( n22170 )  ;
assign n22220 =  ( n16 ) & ( n22140 )  ;
assign n22221 =  ( n16 ) & ( n22142 )  ;
assign n22222 =  ( n16 ) & ( n22144 )  ;
assign n22223 =  ( n16 ) & ( n22146 )  ;
assign n22224 =  ( n16 ) & ( n22148 )  ;
assign n22225 =  ( n16 ) & ( n22150 )  ;
assign n22226 =  ( n16 ) & ( n22152 )  ;
assign n22227 =  ( n16 ) & ( n22154 )  ;
assign n22228 =  ( n16 ) & ( n22156 )  ;
assign n22229 =  ( n16 ) & ( n22158 )  ;
assign n22230 =  ( n16 ) & ( n22160 )  ;
assign n22231 =  ( n16 ) & ( n22162 )  ;
assign n22232 =  ( n16 ) & ( n22164 )  ;
assign n22233 =  ( n16 ) & ( n22166 )  ;
assign n22234 =  ( n16 ) & ( n22168 )  ;
assign n22235 =  ( n16 ) & ( n22170 )  ;
assign n22236 =  ( n17 ) & ( n22140 )  ;
assign n22237 =  ( n17 ) & ( n22142 )  ;
assign n22238 =  ( n17 ) & ( n22144 )  ;
assign n22239 =  ( n17 ) & ( n22146 )  ;
assign n22240 =  ( n17 ) & ( n22148 )  ;
assign n22241 =  ( n17 ) & ( n22150 )  ;
assign n22242 =  ( n17 ) & ( n22152 )  ;
assign n22243 =  ( n17 ) & ( n22154 )  ;
assign n22244 =  ( n17 ) & ( n22156 )  ;
assign n22245 =  ( n17 ) & ( n22158 )  ;
assign n22246 =  ( n17 ) & ( n22160 )  ;
assign n22247 =  ( n17 ) & ( n22162 )  ;
assign n22248 =  ( n17 ) & ( n22164 )  ;
assign n22249 =  ( n17 ) & ( n22166 )  ;
assign n22250 =  ( n17 ) & ( n22168 )  ;
assign n22251 =  ( n17 ) & ( n22170 )  ;
assign n22252 =  ( n18 ) & ( n22140 )  ;
assign n22253 =  ( n18 ) & ( n22142 )  ;
assign n22254 =  ( n18 ) & ( n22144 )  ;
assign n22255 =  ( n18 ) & ( n22146 )  ;
assign n22256 =  ( n18 ) & ( n22148 )  ;
assign n22257 =  ( n18 ) & ( n22150 )  ;
assign n22258 =  ( n18 ) & ( n22152 )  ;
assign n22259 =  ( n18 ) & ( n22154 )  ;
assign n22260 =  ( n18 ) & ( n22156 )  ;
assign n22261 =  ( n18 ) & ( n22158 )  ;
assign n22262 =  ( n18 ) & ( n22160 )  ;
assign n22263 =  ( n18 ) & ( n22162 )  ;
assign n22264 =  ( n18 ) & ( n22164 )  ;
assign n22265 =  ( n18 ) & ( n22166 )  ;
assign n22266 =  ( n18 ) & ( n22168 )  ;
assign n22267 =  ( n18 ) & ( n22170 )  ;
assign n22268 =  ( n19 ) & ( n22140 )  ;
assign n22269 =  ( n19 ) & ( n22142 )  ;
assign n22270 =  ( n19 ) & ( n22144 )  ;
assign n22271 =  ( n19 ) & ( n22146 )  ;
assign n22272 =  ( n19 ) & ( n22148 )  ;
assign n22273 =  ( n19 ) & ( n22150 )  ;
assign n22274 =  ( n19 ) & ( n22152 )  ;
assign n22275 =  ( n19 ) & ( n22154 )  ;
assign n22276 =  ( n19 ) & ( n22156 )  ;
assign n22277 =  ( n19 ) & ( n22158 )  ;
assign n22278 =  ( n19 ) & ( n22160 )  ;
assign n22279 =  ( n19 ) & ( n22162 )  ;
assign n22280 =  ( n19 ) & ( n22164 )  ;
assign n22281 =  ( n19 ) & ( n22166 )  ;
assign n22282 =  ( n19 ) & ( n22168 )  ;
assign n22283 =  ( n19 ) & ( n22170 )  ;
assign n22284 =  ( n20 ) & ( n22140 )  ;
assign n22285 =  ( n20 ) & ( n22142 )  ;
assign n22286 =  ( n20 ) & ( n22144 )  ;
assign n22287 =  ( n20 ) & ( n22146 )  ;
assign n22288 =  ( n20 ) & ( n22148 )  ;
assign n22289 =  ( n20 ) & ( n22150 )  ;
assign n22290 =  ( n20 ) & ( n22152 )  ;
assign n22291 =  ( n20 ) & ( n22154 )  ;
assign n22292 =  ( n20 ) & ( n22156 )  ;
assign n22293 =  ( n20 ) & ( n22158 )  ;
assign n22294 =  ( n20 ) & ( n22160 )  ;
assign n22295 =  ( n20 ) & ( n22162 )  ;
assign n22296 =  ( n20 ) & ( n22164 )  ;
assign n22297 =  ( n20 ) & ( n22166 )  ;
assign n22298 =  ( n20 ) & ( n22168 )  ;
assign n22299 =  ( n20 ) & ( n22170 )  ;
assign n22300 =  ( n21 ) & ( n22140 )  ;
assign n22301 =  ( n21 ) & ( n22142 )  ;
assign n22302 =  ( n21 ) & ( n22144 )  ;
assign n22303 =  ( n21 ) & ( n22146 )  ;
assign n22304 =  ( n21 ) & ( n22148 )  ;
assign n22305 =  ( n21 ) & ( n22150 )  ;
assign n22306 =  ( n21 ) & ( n22152 )  ;
assign n22307 =  ( n21 ) & ( n22154 )  ;
assign n22308 =  ( n21 ) & ( n22156 )  ;
assign n22309 =  ( n21 ) & ( n22158 )  ;
assign n22310 =  ( n21 ) & ( n22160 )  ;
assign n22311 =  ( n21 ) & ( n22162 )  ;
assign n22312 =  ( n21 ) & ( n22164 )  ;
assign n22313 =  ( n21 ) & ( n22166 )  ;
assign n22314 =  ( n21 ) & ( n22168 )  ;
assign n22315 =  ( n21 ) & ( n22170 )  ;
assign n22316 =  ( n22 ) & ( n22140 )  ;
assign n22317 =  ( n22 ) & ( n22142 )  ;
assign n22318 =  ( n22 ) & ( n22144 )  ;
assign n22319 =  ( n22 ) & ( n22146 )  ;
assign n22320 =  ( n22 ) & ( n22148 )  ;
assign n22321 =  ( n22 ) & ( n22150 )  ;
assign n22322 =  ( n22 ) & ( n22152 )  ;
assign n22323 =  ( n22 ) & ( n22154 )  ;
assign n22324 =  ( n22 ) & ( n22156 )  ;
assign n22325 =  ( n22 ) & ( n22158 )  ;
assign n22326 =  ( n22 ) & ( n22160 )  ;
assign n22327 =  ( n22 ) & ( n22162 )  ;
assign n22328 =  ( n22 ) & ( n22164 )  ;
assign n22329 =  ( n22 ) & ( n22166 )  ;
assign n22330 =  ( n22 ) & ( n22168 )  ;
assign n22331 =  ( n22 ) & ( n22170 )  ;
assign n22332 =  ( n23 ) & ( n22140 )  ;
assign n22333 =  ( n23 ) & ( n22142 )  ;
assign n22334 =  ( n23 ) & ( n22144 )  ;
assign n22335 =  ( n23 ) & ( n22146 )  ;
assign n22336 =  ( n23 ) & ( n22148 )  ;
assign n22337 =  ( n23 ) & ( n22150 )  ;
assign n22338 =  ( n23 ) & ( n22152 )  ;
assign n22339 =  ( n23 ) & ( n22154 )  ;
assign n22340 =  ( n23 ) & ( n22156 )  ;
assign n22341 =  ( n23 ) & ( n22158 )  ;
assign n22342 =  ( n23 ) & ( n22160 )  ;
assign n22343 =  ( n23 ) & ( n22162 )  ;
assign n22344 =  ( n23 ) & ( n22164 )  ;
assign n22345 =  ( n23 ) & ( n22166 )  ;
assign n22346 =  ( n23 ) & ( n22168 )  ;
assign n22347 =  ( n23 ) & ( n22170 )  ;
assign n22348 =  ( n24 ) & ( n22140 )  ;
assign n22349 =  ( n24 ) & ( n22142 )  ;
assign n22350 =  ( n24 ) & ( n22144 )  ;
assign n22351 =  ( n24 ) & ( n22146 )  ;
assign n22352 =  ( n24 ) & ( n22148 )  ;
assign n22353 =  ( n24 ) & ( n22150 )  ;
assign n22354 =  ( n24 ) & ( n22152 )  ;
assign n22355 =  ( n24 ) & ( n22154 )  ;
assign n22356 =  ( n24 ) & ( n22156 )  ;
assign n22357 =  ( n24 ) & ( n22158 )  ;
assign n22358 =  ( n24 ) & ( n22160 )  ;
assign n22359 =  ( n24 ) & ( n22162 )  ;
assign n22360 =  ( n24 ) & ( n22164 )  ;
assign n22361 =  ( n24 ) & ( n22166 )  ;
assign n22362 =  ( n24 ) & ( n22168 )  ;
assign n22363 =  ( n24 ) & ( n22170 )  ;
assign n22364 =  ( n25 ) & ( n22140 )  ;
assign n22365 =  ( n25 ) & ( n22142 )  ;
assign n22366 =  ( n25 ) & ( n22144 )  ;
assign n22367 =  ( n25 ) & ( n22146 )  ;
assign n22368 =  ( n25 ) & ( n22148 )  ;
assign n22369 =  ( n25 ) & ( n22150 )  ;
assign n22370 =  ( n25 ) & ( n22152 )  ;
assign n22371 =  ( n25 ) & ( n22154 )  ;
assign n22372 =  ( n25 ) & ( n22156 )  ;
assign n22373 =  ( n25 ) & ( n22158 )  ;
assign n22374 =  ( n25 ) & ( n22160 )  ;
assign n22375 =  ( n25 ) & ( n22162 )  ;
assign n22376 =  ( n25 ) & ( n22164 )  ;
assign n22377 =  ( n25 ) & ( n22166 )  ;
assign n22378 =  ( n25 ) & ( n22168 )  ;
assign n22379 =  ( n25 ) & ( n22170 )  ;
assign n22380 =  ( n26 ) & ( n22140 )  ;
assign n22381 =  ( n26 ) & ( n22142 )  ;
assign n22382 =  ( n26 ) & ( n22144 )  ;
assign n22383 =  ( n26 ) & ( n22146 )  ;
assign n22384 =  ( n26 ) & ( n22148 )  ;
assign n22385 =  ( n26 ) & ( n22150 )  ;
assign n22386 =  ( n26 ) & ( n22152 )  ;
assign n22387 =  ( n26 ) & ( n22154 )  ;
assign n22388 =  ( n26 ) & ( n22156 )  ;
assign n22389 =  ( n26 ) & ( n22158 )  ;
assign n22390 =  ( n26 ) & ( n22160 )  ;
assign n22391 =  ( n26 ) & ( n22162 )  ;
assign n22392 =  ( n26 ) & ( n22164 )  ;
assign n22393 =  ( n26 ) & ( n22166 )  ;
assign n22394 =  ( n26 ) & ( n22168 )  ;
assign n22395 =  ( n26 ) & ( n22170 )  ;
assign n22396 =  ( n27 ) & ( n22140 )  ;
assign n22397 =  ( n27 ) & ( n22142 )  ;
assign n22398 =  ( n27 ) & ( n22144 )  ;
assign n22399 =  ( n27 ) & ( n22146 )  ;
assign n22400 =  ( n27 ) & ( n22148 )  ;
assign n22401 =  ( n27 ) & ( n22150 )  ;
assign n22402 =  ( n27 ) & ( n22152 )  ;
assign n22403 =  ( n27 ) & ( n22154 )  ;
assign n22404 =  ( n27 ) & ( n22156 )  ;
assign n22405 =  ( n27 ) & ( n22158 )  ;
assign n22406 =  ( n27 ) & ( n22160 )  ;
assign n22407 =  ( n27 ) & ( n22162 )  ;
assign n22408 =  ( n27 ) & ( n22164 )  ;
assign n22409 =  ( n27 ) & ( n22166 )  ;
assign n22410 =  ( n27 ) & ( n22168 )  ;
assign n22411 =  ( n27 ) & ( n22170 )  ;
assign n22412 =  ( n28 ) & ( n22140 )  ;
assign n22413 =  ( n28 ) & ( n22142 )  ;
assign n22414 =  ( n28 ) & ( n22144 )  ;
assign n22415 =  ( n28 ) & ( n22146 )  ;
assign n22416 =  ( n28 ) & ( n22148 )  ;
assign n22417 =  ( n28 ) & ( n22150 )  ;
assign n22418 =  ( n28 ) & ( n22152 )  ;
assign n22419 =  ( n28 ) & ( n22154 )  ;
assign n22420 =  ( n28 ) & ( n22156 )  ;
assign n22421 =  ( n28 ) & ( n22158 )  ;
assign n22422 =  ( n28 ) & ( n22160 )  ;
assign n22423 =  ( n28 ) & ( n22162 )  ;
assign n22424 =  ( n28 ) & ( n22164 )  ;
assign n22425 =  ( n28 ) & ( n22166 )  ;
assign n22426 =  ( n28 ) & ( n22168 )  ;
assign n22427 =  ( n28 ) & ( n22170 )  ;
assign n22428 =  ( n29 ) & ( n22140 )  ;
assign n22429 =  ( n29 ) & ( n22142 )  ;
assign n22430 =  ( n29 ) & ( n22144 )  ;
assign n22431 =  ( n29 ) & ( n22146 )  ;
assign n22432 =  ( n29 ) & ( n22148 )  ;
assign n22433 =  ( n29 ) & ( n22150 )  ;
assign n22434 =  ( n29 ) & ( n22152 )  ;
assign n22435 =  ( n29 ) & ( n22154 )  ;
assign n22436 =  ( n29 ) & ( n22156 )  ;
assign n22437 =  ( n29 ) & ( n22158 )  ;
assign n22438 =  ( n29 ) & ( n22160 )  ;
assign n22439 =  ( n29 ) & ( n22162 )  ;
assign n22440 =  ( n29 ) & ( n22164 )  ;
assign n22441 =  ( n29 ) & ( n22166 )  ;
assign n22442 =  ( n29 ) & ( n22168 )  ;
assign n22443 =  ( n29 ) & ( n22170 )  ;
assign n22444 =  ( n30 ) & ( n22140 )  ;
assign n22445 =  ( n30 ) & ( n22142 )  ;
assign n22446 =  ( n30 ) & ( n22144 )  ;
assign n22447 =  ( n30 ) & ( n22146 )  ;
assign n22448 =  ( n30 ) & ( n22148 )  ;
assign n22449 =  ( n30 ) & ( n22150 )  ;
assign n22450 =  ( n30 ) & ( n22152 )  ;
assign n22451 =  ( n30 ) & ( n22154 )  ;
assign n22452 =  ( n30 ) & ( n22156 )  ;
assign n22453 =  ( n30 ) & ( n22158 )  ;
assign n22454 =  ( n30 ) & ( n22160 )  ;
assign n22455 =  ( n30 ) & ( n22162 )  ;
assign n22456 =  ( n30 ) & ( n22164 )  ;
assign n22457 =  ( n30 ) & ( n22166 )  ;
assign n22458 =  ( n30 ) & ( n22168 )  ;
assign n22459 =  ( n30 ) & ( n22170 )  ;
assign n22460 =  ( n31 ) & ( n22140 )  ;
assign n22461 =  ( n31 ) & ( n22142 )  ;
assign n22462 =  ( n31 ) & ( n22144 )  ;
assign n22463 =  ( n31 ) & ( n22146 )  ;
assign n22464 =  ( n31 ) & ( n22148 )  ;
assign n22465 =  ( n31 ) & ( n22150 )  ;
assign n22466 =  ( n31 ) & ( n22152 )  ;
assign n22467 =  ( n31 ) & ( n22154 )  ;
assign n22468 =  ( n31 ) & ( n22156 )  ;
assign n22469 =  ( n31 ) & ( n22158 )  ;
assign n22470 =  ( n31 ) & ( n22160 )  ;
assign n22471 =  ( n31 ) & ( n22162 )  ;
assign n22472 =  ( n31 ) & ( n22164 )  ;
assign n22473 =  ( n31 ) & ( n22166 )  ;
assign n22474 =  ( n31 ) & ( n22168 )  ;
assign n22475 =  ( n31 ) & ( n22170 )  ;
assign n22476 =  ( n32 ) & ( n22140 )  ;
assign n22477 =  ( n32 ) & ( n22142 )  ;
assign n22478 =  ( n32 ) & ( n22144 )  ;
assign n22479 =  ( n32 ) & ( n22146 )  ;
assign n22480 =  ( n32 ) & ( n22148 )  ;
assign n22481 =  ( n32 ) & ( n22150 )  ;
assign n22482 =  ( n32 ) & ( n22152 )  ;
assign n22483 =  ( n32 ) & ( n22154 )  ;
assign n22484 =  ( n32 ) & ( n22156 )  ;
assign n22485 =  ( n32 ) & ( n22158 )  ;
assign n22486 =  ( n32 ) & ( n22160 )  ;
assign n22487 =  ( n32 ) & ( n22162 )  ;
assign n22488 =  ( n32 ) & ( n22164 )  ;
assign n22489 =  ( n32 ) & ( n22166 )  ;
assign n22490 =  ( n32 ) & ( n22168 )  ;
assign n22491 =  ( n32 ) & ( n22170 )  ;
assign n22492 =  ( n33 ) & ( n22140 )  ;
assign n22493 =  ( n33 ) & ( n22142 )  ;
assign n22494 =  ( n33 ) & ( n22144 )  ;
assign n22495 =  ( n33 ) & ( n22146 )  ;
assign n22496 =  ( n33 ) & ( n22148 )  ;
assign n22497 =  ( n33 ) & ( n22150 )  ;
assign n22498 =  ( n33 ) & ( n22152 )  ;
assign n22499 =  ( n33 ) & ( n22154 )  ;
assign n22500 =  ( n33 ) & ( n22156 )  ;
assign n22501 =  ( n33 ) & ( n22158 )  ;
assign n22502 =  ( n33 ) & ( n22160 )  ;
assign n22503 =  ( n33 ) & ( n22162 )  ;
assign n22504 =  ( n33 ) & ( n22164 )  ;
assign n22505 =  ( n33 ) & ( n22166 )  ;
assign n22506 =  ( n33 ) & ( n22168 )  ;
assign n22507 =  ( n33 ) & ( n22170 )  ;
assign n22508 =  ( n34 ) & ( n22140 )  ;
assign n22509 =  ( n34 ) & ( n22142 )  ;
assign n22510 =  ( n34 ) & ( n22144 )  ;
assign n22511 =  ( n34 ) & ( n22146 )  ;
assign n22512 =  ( n34 ) & ( n22148 )  ;
assign n22513 =  ( n34 ) & ( n22150 )  ;
assign n22514 =  ( n34 ) & ( n22152 )  ;
assign n22515 =  ( n34 ) & ( n22154 )  ;
assign n22516 =  ( n34 ) & ( n22156 )  ;
assign n22517 =  ( n34 ) & ( n22158 )  ;
assign n22518 =  ( n34 ) & ( n22160 )  ;
assign n22519 =  ( n34 ) & ( n22162 )  ;
assign n22520 =  ( n34 ) & ( n22164 )  ;
assign n22521 =  ( n34 ) & ( n22166 )  ;
assign n22522 =  ( n34 ) & ( n22168 )  ;
assign n22523 =  ( n34 ) & ( n22170 )  ;
assign n22524 =  ( n35 ) & ( n22140 )  ;
assign n22525 =  ( n35 ) & ( n22142 )  ;
assign n22526 =  ( n35 ) & ( n22144 )  ;
assign n22527 =  ( n35 ) & ( n22146 )  ;
assign n22528 =  ( n35 ) & ( n22148 )  ;
assign n22529 =  ( n35 ) & ( n22150 )  ;
assign n22530 =  ( n35 ) & ( n22152 )  ;
assign n22531 =  ( n35 ) & ( n22154 )  ;
assign n22532 =  ( n35 ) & ( n22156 )  ;
assign n22533 =  ( n35 ) & ( n22158 )  ;
assign n22534 =  ( n35 ) & ( n22160 )  ;
assign n22535 =  ( n35 ) & ( n22162 )  ;
assign n22536 =  ( n35 ) & ( n22164 )  ;
assign n22537 =  ( n35 ) & ( n22166 )  ;
assign n22538 =  ( n35 ) & ( n22168 )  ;
assign n22539 =  ( n35 ) & ( n22170 )  ;
assign n22540 =  ( n36 ) & ( n22140 )  ;
assign n22541 =  ( n36 ) & ( n22142 )  ;
assign n22542 =  ( n36 ) & ( n22144 )  ;
assign n22543 =  ( n36 ) & ( n22146 )  ;
assign n22544 =  ( n36 ) & ( n22148 )  ;
assign n22545 =  ( n36 ) & ( n22150 )  ;
assign n22546 =  ( n36 ) & ( n22152 )  ;
assign n22547 =  ( n36 ) & ( n22154 )  ;
assign n22548 =  ( n36 ) & ( n22156 )  ;
assign n22549 =  ( n36 ) & ( n22158 )  ;
assign n22550 =  ( n36 ) & ( n22160 )  ;
assign n22551 =  ( n36 ) & ( n22162 )  ;
assign n22552 =  ( n36 ) & ( n22164 )  ;
assign n22553 =  ( n36 ) & ( n22166 )  ;
assign n22554 =  ( n36 ) & ( n22168 )  ;
assign n22555 =  ( n36 ) & ( n22170 )  ;
assign n22556 =  ( n37 ) & ( n22140 )  ;
assign n22557 =  ( n37 ) & ( n22142 )  ;
assign n22558 =  ( n37 ) & ( n22144 )  ;
assign n22559 =  ( n37 ) & ( n22146 )  ;
assign n22560 =  ( n37 ) & ( n22148 )  ;
assign n22561 =  ( n37 ) & ( n22150 )  ;
assign n22562 =  ( n37 ) & ( n22152 )  ;
assign n22563 =  ( n37 ) & ( n22154 )  ;
assign n22564 =  ( n37 ) & ( n22156 )  ;
assign n22565 =  ( n37 ) & ( n22158 )  ;
assign n22566 =  ( n37 ) & ( n22160 )  ;
assign n22567 =  ( n37 ) & ( n22162 )  ;
assign n22568 =  ( n37 ) & ( n22164 )  ;
assign n22569 =  ( n37 ) & ( n22166 )  ;
assign n22570 =  ( n37 ) & ( n22168 )  ;
assign n22571 =  ( n37 ) & ( n22170 )  ;
assign n22572 =  ( n38 ) & ( n22140 )  ;
assign n22573 =  ( n38 ) & ( n22142 )  ;
assign n22574 =  ( n38 ) & ( n22144 )  ;
assign n22575 =  ( n38 ) & ( n22146 )  ;
assign n22576 =  ( n38 ) & ( n22148 )  ;
assign n22577 =  ( n38 ) & ( n22150 )  ;
assign n22578 =  ( n38 ) & ( n22152 )  ;
assign n22579 =  ( n38 ) & ( n22154 )  ;
assign n22580 =  ( n38 ) & ( n22156 )  ;
assign n22581 =  ( n38 ) & ( n22158 )  ;
assign n22582 =  ( n38 ) & ( n22160 )  ;
assign n22583 =  ( n38 ) & ( n22162 )  ;
assign n22584 =  ( n38 ) & ( n22164 )  ;
assign n22585 =  ( n38 ) & ( n22166 )  ;
assign n22586 =  ( n38 ) & ( n22168 )  ;
assign n22587 =  ( n38 ) & ( n22170 )  ;
assign n22588 =  ( n39 ) & ( n22140 )  ;
assign n22589 =  ( n39 ) & ( n22142 )  ;
assign n22590 =  ( n39 ) & ( n22144 )  ;
assign n22591 =  ( n39 ) & ( n22146 )  ;
assign n22592 =  ( n39 ) & ( n22148 )  ;
assign n22593 =  ( n39 ) & ( n22150 )  ;
assign n22594 =  ( n39 ) & ( n22152 )  ;
assign n22595 =  ( n39 ) & ( n22154 )  ;
assign n22596 =  ( n39 ) & ( n22156 )  ;
assign n22597 =  ( n39 ) & ( n22158 )  ;
assign n22598 =  ( n39 ) & ( n22160 )  ;
assign n22599 =  ( n39 ) & ( n22162 )  ;
assign n22600 =  ( n39 ) & ( n22164 )  ;
assign n22601 =  ( n39 ) & ( n22166 )  ;
assign n22602 =  ( n39 ) & ( n22168 )  ;
assign n22603 =  ( n39 ) & ( n22170 )  ;
assign n22604 =  ( n40 ) & ( n22140 )  ;
assign n22605 =  ( n40 ) & ( n22142 )  ;
assign n22606 =  ( n40 ) & ( n22144 )  ;
assign n22607 =  ( n40 ) & ( n22146 )  ;
assign n22608 =  ( n40 ) & ( n22148 )  ;
assign n22609 =  ( n40 ) & ( n22150 )  ;
assign n22610 =  ( n40 ) & ( n22152 )  ;
assign n22611 =  ( n40 ) & ( n22154 )  ;
assign n22612 =  ( n40 ) & ( n22156 )  ;
assign n22613 =  ( n40 ) & ( n22158 )  ;
assign n22614 =  ( n40 ) & ( n22160 )  ;
assign n22615 =  ( n40 ) & ( n22162 )  ;
assign n22616 =  ( n40 ) & ( n22164 )  ;
assign n22617 =  ( n40 ) & ( n22166 )  ;
assign n22618 =  ( n40 ) & ( n22168 )  ;
assign n22619 =  ( n40 ) & ( n22170 )  ;
assign n22620 =  ( n41 ) & ( n22140 )  ;
assign n22621 =  ( n41 ) & ( n22142 )  ;
assign n22622 =  ( n41 ) & ( n22144 )  ;
assign n22623 =  ( n41 ) & ( n22146 )  ;
assign n22624 =  ( n41 ) & ( n22148 )  ;
assign n22625 =  ( n41 ) & ( n22150 )  ;
assign n22626 =  ( n41 ) & ( n22152 )  ;
assign n22627 =  ( n41 ) & ( n22154 )  ;
assign n22628 =  ( n41 ) & ( n22156 )  ;
assign n22629 =  ( n41 ) & ( n22158 )  ;
assign n22630 =  ( n41 ) & ( n22160 )  ;
assign n22631 =  ( n41 ) & ( n22162 )  ;
assign n22632 =  ( n41 ) & ( n22164 )  ;
assign n22633 =  ( n41 ) & ( n22166 )  ;
assign n22634 =  ( n41 ) & ( n22168 )  ;
assign n22635 =  ( n41 ) & ( n22170 )  ;
assign n22636 =  ( n42 ) & ( n22140 )  ;
assign n22637 =  ( n42 ) & ( n22142 )  ;
assign n22638 =  ( n42 ) & ( n22144 )  ;
assign n22639 =  ( n42 ) & ( n22146 )  ;
assign n22640 =  ( n42 ) & ( n22148 )  ;
assign n22641 =  ( n42 ) & ( n22150 )  ;
assign n22642 =  ( n42 ) & ( n22152 )  ;
assign n22643 =  ( n42 ) & ( n22154 )  ;
assign n22644 =  ( n42 ) & ( n22156 )  ;
assign n22645 =  ( n42 ) & ( n22158 )  ;
assign n22646 =  ( n42 ) & ( n22160 )  ;
assign n22647 =  ( n42 ) & ( n22162 )  ;
assign n22648 =  ( n42 ) & ( n22164 )  ;
assign n22649 =  ( n42 ) & ( n22166 )  ;
assign n22650 =  ( n42 ) & ( n22168 )  ;
assign n22651 =  ( n42 ) & ( n22170 )  ;
assign n22652 =  ( n43 ) & ( n22140 )  ;
assign n22653 =  ( n43 ) & ( n22142 )  ;
assign n22654 =  ( n43 ) & ( n22144 )  ;
assign n22655 =  ( n43 ) & ( n22146 )  ;
assign n22656 =  ( n43 ) & ( n22148 )  ;
assign n22657 =  ( n43 ) & ( n22150 )  ;
assign n22658 =  ( n43 ) & ( n22152 )  ;
assign n22659 =  ( n43 ) & ( n22154 )  ;
assign n22660 =  ( n43 ) & ( n22156 )  ;
assign n22661 =  ( n43 ) & ( n22158 )  ;
assign n22662 =  ( n43 ) & ( n22160 )  ;
assign n22663 =  ( n43 ) & ( n22162 )  ;
assign n22664 =  ( n43 ) & ( n22164 )  ;
assign n22665 =  ( n43 ) & ( n22166 )  ;
assign n22666 =  ( n43 ) & ( n22168 )  ;
assign n22667 =  ( n43 ) & ( n22170 )  ;
assign n22668 =  ( n22667 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n22669 =  ( n22666 ) ? ( VREG_0_1 ) : ( n22668 ) ;
assign n22670 =  ( n22665 ) ? ( VREG_0_2 ) : ( n22669 ) ;
assign n22671 =  ( n22664 ) ? ( VREG_0_3 ) : ( n22670 ) ;
assign n22672 =  ( n22663 ) ? ( VREG_0_4 ) : ( n22671 ) ;
assign n22673 =  ( n22662 ) ? ( VREG_0_5 ) : ( n22672 ) ;
assign n22674 =  ( n22661 ) ? ( VREG_0_6 ) : ( n22673 ) ;
assign n22675 =  ( n22660 ) ? ( VREG_0_7 ) : ( n22674 ) ;
assign n22676 =  ( n22659 ) ? ( VREG_0_8 ) : ( n22675 ) ;
assign n22677 =  ( n22658 ) ? ( VREG_0_9 ) : ( n22676 ) ;
assign n22678 =  ( n22657 ) ? ( VREG_0_10 ) : ( n22677 ) ;
assign n22679 =  ( n22656 ) ? ( VREG_0_11 ) : ( n22678 ) ;
assign n22680 =  ( n22655 ) ? ( VREG_0_12 ) : ( n22679 ) ;
assign n22681 =  ( n22654 ) ? ( VREG_0_13 ) : ( n22680 ) ;
assign n22682 =  ( n22653 ) ? ( VREG_0_14 ) : ( n22681 ) ;
assign n22683 =  ( n22652 ) ? ( VREG_0_15 ) : ( n22682 ) ;
assign n22684 =  ( n22651 ) ? ( VREG_1_0 ) : ( n22683 ) ;
assign n22685 =  ( n22650 ) ? ( VREG_1_1 ) : ( n22684 ) ;
assign n22686 =  ( n22649 ) ? ( VREG_1_2 ) : ( n22685 ) ;
assign n22687 =  ( n22648 ) ? ( VREG_1_3 ) : ( n22686 ) ;
assign n22688 =  ( n22647 ) ? ( VREG_1_4 ) : ( n22687 ) ;
assign n22689 =  ( n22646 ) ? ( VREG_1_5 ) : ( n22688 ) ;
assign n22690 =  ( n22645 ) ? ( VREG_1_6 ) : ( n22689 ) ;
assign n22691 =  ( n22644 ) ? ( VREG_1_7 ) : ( n22690 ) ;
assign n22692 =  ( n22643 ) ? ( VREG_1_8 ) : ( n22691 ) ;
assign n22693 =  ( n22642 ) ? ( VREG_1_9 ) : ( n22692 ) ;
assign n22694 =  ( n22641 ) ? ( VREG_1_10 ) : ( n22693 ) ;
assign n22695 =  ( n22640 ) ? ( VREG_1_11 ) : ( n22694 ) ;
assign n22696 =  ( n22639 ) ? ( VREG_1_12 ) : ( n22695 ) ;
assign n22697 =  ( n22638 ) ? ( VREG_1_13 ) : ( n22696 ) ;
assign n22698 =  ( n22637 ) ? ( VREG_1_14 ) : ( n22697 ) ;
assign n22699 =  ( n22636 ) ? ( VREG_1_15 ) : ( n22698 ) ;
assign n22700 =  ( n22635 ) ? ( VREG_2_0 ) : ( n22699 ) ;
assign n22701 =  ( n22634 ) ? ( VREG_2_1 ) : ( n22700 ) ;
assign n22702 =  ( n22633 ) ? ( VREG_2_2 ) : ( n22701 ) ;
assign n22703 =  ( n22632 ) ? ( VREG_2_3 ) : ( n22702 ) ;
assign n22704 =  ( n22631 ) ? ( VREG_2_4 ) : ( n22703 ) ;
assign n22705 =  ( n22630 ) ? ( VREG_2_5 ) : ( n22704 ) ;
assign n22706 =  ( n22629 ) ? ( VREG_2_6 ) : ( n22705 ) ;
assign n22707 =  ( n22628 ) ? ( VREG_2_7 ) : ( n22706 ) ;
assign n22708 =  ( n22627 ) ? ( VREG_2_8 ) : ( n22707 ) ;
assign n22709 =  ( n22626 ) ? ( VREG_2_9 ) : ( n22708 ) ;
assign n22710 =  ( n22625 ) ? ( VREG_2_10 ) : ( n22709 ) ;
assign n22711 =  ( n22624 ) ? ( VREG_2_11 ) : ( n22710 ) ;
assign n22712 =  ( n22623 ) ? ( VREG_2_12 ) : ( n22711 ) ;
assign n22713 =  ( n22622 ) ? ( VREG_2_13 ) : ( n22712 ) ;
assign n22714 =  ( n22621 ) ? ( VREG_2_14 ) : ( n22713 ) ;
assign n22715 =  ( n22620 ) ? ( VREG_2_15 ) : ( n22714 ) ;
assign n22716 =  ( n22619 ) ? ( VREG_3_0 ) : ( n22715 ) ;
assign n22717 =  ( n22618 ) ? ( VREG_3_1 ) : ( n22716 ) ;
assign n22718 =  ( n22617 ) ? ( VREG_3_2 ) : ( n22717 ) ;
assign n22719 =  ( n22616 ) ? ( VREG_3_3 ) : ( n22718 ) ;
assign n22720 =  ( n22615 ) ? ( VREG_3_4 ) : ( n22719 ) ;
assign n22721 =  ( n22614 ) ? ( VREG_3_5 ) : ( n22720 ) ;
assign n22722 =  ( n22613 ) ? ( VREG_3_6 ) : ( n22721 ) ;
assign n22723 =  ( n22612 ) ? ( VREG_3_7 ) : ( n22722 ) ;
assign n22724 =  ( n22611 ) ? ( VREG_3_8 ) : ( n22723 ) ;
assign n22725 =  ( n22610 ) ? ( VREG_3_9 ) : ( n22724 ) ;
assign n22726 =  ( n22609 ) ? ( VREG_3_10 ) : ( n22725 ) ;
assign n22727 =  ( n22608 ) ? ( VREG_3_11 ) : ( n22726 ) ;
assign n22728 =  ( n22607 ) ? ( VREG_3_12 ) : ( n22727 ) ;
assign n22729 =  ( n22606 ) ? ( VREG_3_13 ) : ( n22728 ) ;
assign n22730 =  ( n22605 ) ? ( VREG_3_14 ) : ( n22729 ) ;
assign n22731 =  ( n22604 ) ? ( VREG_3_15 ) : ( n22730 ) ;
assign n22732 =  ( n22603 ) ? ( VREG_4_0 ) : ( n22731 ) ;
assign n22733 =  ( n22602 ) ? ( VREG_4_1 ) : ( n22732 ) ;
assign n22734 =  ( n22601 ) ? ( VREG_4_2 ) : ( n22733 ) ;
assign n22735 =  ( n22600 ) ? ( VREG_4_3 ) : ( n22734 ) ;
assign n22736 =  ( n22599 ) ? ( VREG_4_4 ) : ( n22735 ) ;
assign n22737 =  ( n22598 ) ? ( VREG_4_5 ) : ( n22736 ) ;
assign n22738 =  ( n22597 ) ? ( VREG_4_6 ) : ( n22737 ) ;
assign n22739 =  ( n22596 ) ? ( VREG_4_7 ) : ( n22738 ) ;
assign n22740 =  ( n22595 ) ? ( VREG_4_8 ) : ( n22739 ) ;
assign n22741 =  ( n22594 ) ? ( VREG_4_9 ) : ( n22740 ) ;
assign n22742 =  ( n22593 ) ? ( VREG_4_10 ) : ( n22741 ) ;
assign n22743 =  ( n22592 ) ? ( VREG_4_11 ) : ( n22742 ) ;
assign n22744 =  ( n22591 ) ? ( VREG_4_12 ) : ( n22743 ) ;
assign n22745 =  ( n22590 ) ? ( VREG_4_13 ) : ( n22744 ) ;
assign n22746 =  ( n22589 ) ? ( VREG_4_14 ) : ( n22745 ) ;
assign n22747 =  ( n22588 ) ? ( VREG_4_15 ) : ( n22746 ) ;
assign n22748 =  ( n22587 ) ? ( VREG_5_0 ) : ( n22747 ) ;
assign n22749 =  ( n22586 ) ? ( VREG_5_1 ) : ( n22748 ) ;
assign n22750 =  ( n22585 ) ? ( VREG_5_2 ) : ( n22749 ) ;
assign n22751 =  ( n22584 ) ? ( VREG_5_3 ) : ( n22750 ) ;
assign n22752 =  ( n22583 ) ? ( VREG_5_4 ) : ( n22751 ) ;
assign n22753 =  ( n22582 ) ? ( VREG_5_5 ) : ( n22752 ) ;
assign n22754 =  ( n22581 ) ? ( VREG_5_6 ) : ( n22753 ) ;
assign n22755 =  ( n22580 ) ? ( VREG_5_7 ) : ( n22754 ) ;
assign n22756 =  ( n22579 ) ? ( VREG_5_8 ) : ( n22755 ) ;
assign n22757 =  ( n22578 ) ? ( VREG_5_9 ) : ( n22756 ) ;
assign n22758 =  ( n22577 ) ? ( VREG_5_10 ) : ( n22757 ) ;
assign n22759 =  ( n22576 ) ? ( VREG_5_11 ) : ( n22758 ) ;
assign n22760 =  ( n22575 ) ? ( VREG_5_12 ) : ( n22759 ) ;
assign n22761 =  ( n22574 ) ? ( VREG_5_13 ) : ( n22760 ) ;
assign n22762 =  ( n22573 ) ? ( VREG_5_14 ) : ( n22761 ) ;
assign n22763 =  ( n22572 ) ? ( VREG_5_15 ) : ( n22762 ) ;
assign n22764 =  ( n22571 ) ? ( VREG_6_0 ) : ( n22763 ) ;
assign n22765 =  ( n22570 ) ? ( VREG_6_1 ) : ( n22764 ) ;
assign n22766 =  ( n22569 ) ? ( VREG_6_2 ) : ( n22765 ) ;
assign n22767 =  ( n22568 ) ? ( VREG_6_3 ) : ( n22766 ) ;
assign n22768 =  ( n22567 ) ? ( VREG_6_4 ) : ( n22767 ) ;
assign n22769 =  ( n22566 ) ? ( VREG_6_5 ) : ( n22768 ) ;
assign n22770 =  ( n22565 ) ? ( VREG_6_6 ) : ( n22769 ) ;
assign n22771 =  ( n22564 ) ? ( VREG_6_7 ) : ( n22770 ) ;
assign n22772 =  ( n22563 ) ? ( VREG_6_8 ) : ( n22771 ) ;
assign n22773 =  ( n22562 ) ? ( VREG_6_9 ) : ( n22772 ) ;
assign n22774 =  ( n22561 ) ? ( VREG_6_10 ) : ( n22773 ) ;
assign n22775 =  ( n22560 ) ? ( VREG_6_11 ) : ( n22774 ) ;
assign n22776 =  ( n22559 ) ? ( VREG_6_12 ) : ( n22775 ) ;
assign n22777 =  ( n22558 ) ? ( VREG_6_13 ) : ( n22776 ) ;
assign n22778 =  ( n22557 ) ? ( VREG_6_14 ) : ( n22777 ) ;
assign n22779 =  ( n22556 ) ? ( VREG_6_15 ) : ( n22778 ) ;
assign n22780 =  ( n22555 ) ? ( VREG_7_0 ) : ( n22779 ) ;
assign n22781 =  ( n22554 ) ? ( VREG_7_1 ) : ( n22780 ) ;
assign n22782 =  ( n22553 ) ? ( VREG_7_2 ) : ( n22781 ) ;
assign n22783 =  ( n22552 ) ? ( VREG_7_3 ) : ( n22782 ) ;
assign n22784 =  ( n22551 ) ? ( VREG_7_4 ) : ( n22783 ) ;
assign n22785 =  ( n22550 ) ? ( VREG_7_5 ) : ( n22784 ) ;
assign n22786 =  ( n22549 ) ? ( VREG_7_6 ) : ( n22785 ) ;
assign n22787 =  ( n22548 ) ? ( VREG_7_7 ) : ( n22786 ) ;
assign n22788 =  ( n22547 ) ? ( VREG_7_8 ) : ( n22787 ) ;
assign n22789 =  ( n22546 ) ? ( VREG_7_9 ) : ( n22788 ) ;
assign n22790 =  ( n22545 ) ? ( VREG_7_10 ) : ( n22789 ) ;
assign n22791 =  ( n22544 ) ? ( VREG_7_11 ) : ( n22790 ) ;
assign n22792 =  ( n22543 ) ? ( VREG_7_12 ) : ( n22791 ) ;
assign n22793 =  ( n22542 ) ? ( VREG_7_13 ) : ( n22792 ) ;
assign n22794 =  ( n22541 ) ? ( VREG_7_14 ) : ( n22793 ) ;
assign n22795 =  ( n22540 ) ? ( VREG_7_15 ) : ( n22794 ) ;
assign n22796 =  ( n22539 ) ? ( VREG_8_0 ) : ( n22795 ) ;
assign n22797 =  ( n22538 ) ? ( VREG_8_1 ) : ( n22796 ) ;
assign n22798 =  ( n22537 ) ? ( VREG_8_2 ) : ( n22797 ) ;
assign n22799 =  ( n22536 ) ? ( VREG_8_3 ) : ( n22798 ) ;
assign n22800 =  ( n22535 ) ? ( VREG_8_4 ) : ( n22799 ) ;
assign n22801 =  ( n22534 ) ? ( VREG_8_5 ) : ( n22800 ) ;
assign n22802 =  ( n22533 ) ? ( VREG_8_6 ) : ( n22801 ) ;
assign n22803 =  ( n22532 ) ? ( VREG_8_7 ) : ( n22802 ) ;
assign n22804 =  ( n22531 ) ? ( VREG_8_8 ) : ( n22803 ) ;
assign n22805 =  ( n22530 ) ? ( VREG_8_9 ) : ( n22804 ) ;
assign n22806 =  ( n22529 ) ? ( VREG_8_10 ) : ( n22805 ) ;
assign n22807 =  ( n22528 ) ? ( VREG_8_11 ) : ( n22806 ) ;
assign n22808 =  ( n22527 ) ? ( VREG_8_12 ) : ( n22807 ) ;
assign n22809 =  ( n22526 ) ? ( VREG_8_13 ) : ( n22808 ) ;
assign n22810 =  ( n22525 ) ? ( VREG_8_14 ) : ( n22809 ) ;
assign n22811 =  ( n22524 ) ? ( VREG_8_15 ) : ( n22810 ) ;
assign n22812 =  ( n22523 ) ? ( VREG_9_0 ) : ( n22811 ) ;
assign n22813 =  ( n22522 ) ? ( VREG_9_1 ) : ( n22812 ) ;
assign n22814 =  ( n22521 ) ? ( VREG_9_2 ) : ( n22813 ) ;
assign n22815 =  ( n22520 ) ? ( VREG_9_3 ) : ( n22814 ) ;
assign n22816 =  ( n22519 ) ? ( VREG_9_4 ) : ( n22815 ) ;
assign n22817 =  ( n22518 ) ? ( VREG_9_5 ) : ( n22816 ) ;
assign n22818 =  ( n22517 ) ? ( VREG_9_6 ) : ( n22817 ) ;
assign n22819 =  ( n22516 ) ? ( VREG_9_7 ) : ( n22818 ) ;
assign n22820 =  ( n22515 ) ? ( VREG_9_8 ) : ( n22819 ) ;
assign n22821 =  ( n22514 ) ? ( VREG_9_9 ) : ( n22820 ) ;
assign n22822 =  ( n22513 ) ? ( VREG_9_10 ) : ( n22821 ) ;
assign n22823 =  ( n22512 ) ? ( VREG_9_11 ) : ( n22822 ) ;
assign n22824 =  ( n22511 ) ? ( VREG_9_12 ) : ( n22823 ) ;
assign n22825 =  ( n22510 ) ? ( VREG_9_13 ) : ( n22824 ) ;
assign n22826 =  ( n22509 ) ? ( VREG_9_14 ) : ( n22825 ) ;
assign n22827 =  ( n22508 ) ? ( VREG_9_15 ) : ( n22826 ) ;
assign n22828 =  ( n22507 ) ? ( VREG_10_0 ) : ( n22827 ) ;
assign n22829 =  ( n22506 ) ? ( VREG_10_1 ) : ( n22828 ) ;
assign n22830 =  ( n22505 ) ? ( VREG_10_2 ) : ( n22829 ) ;
assign n22831 =  ( n22504 ) ? ( VREG_10_3 ) : ( n22830 ) ;
assign n22832 =  ( n22503 ) ? ( VREG_10_4 ) : ( n22831 ) ;
assign n22833 =  ( n22502 ) ? ( VREG_10_5 ) : ( n22832 ) ;
assign n22834 =  ( n22501 ) ? ( VREG_10_6 ) : ( n22833 ) ;
assign n22835 =  ( n22500 ) ? ( VREG_10_7 ) : ( n22834 ) ;
assign n22836 =  ( n22499 ) ? ( VREG_10_8 ) : ( n22835 ) ;
assign n22837 =  ( n22498 ) ? ( VREG_10_9 ) : ( n22836 ) ;
assign n22838 =  ( n22497 ) ? ( VREG_10_10 ) : ( n22837 ) ;
assign n22839 =  ( n22496 ) ? ( VREG_10_11 ) : ( n22838 ) ;
assign n22840 =  ( n22495 ) ? ( VREG_10_12 ) : ( n22839 ) ;
assign n22841 =  ( n22494 ) ? ( VREG_10_13 ) : ( n22840 ) ;
assign n22842 =  ( n22493 ) ? ( VREG_10_14 ) : ( n22841 ) ;
assign n22843 =  ( n22492 ) ? ( VREG_10_15 ) : ( n22842 ) ;
assign n22844 =  ( n22491 ) ? ( VREG_11_0 ) : ( n22843 ) ;
assign n22845 =  ( n22490 ) ? ( VREG_11_1 ) : ( n22844 ) ;
assign n22846 =  ( n22489 ) ? ( VREG_11_2 ) : ( n22845 ) ;
assign n22847 =  ( n22488 ) ? ( VREG_11_3 ) : ( n22846 ) ;
assign n22848 =  ( n22487 ) ? ( VREG_11_4 ) : ( n22847 ) ;
assign n22849 =  ( n22486 ) ? ( VREG_11_5 ) : ( n22848 ) ;
assign n22850 =  ( n22485 ) ? ( VREG_11_6 ) : ( n22849 ) ;
assign n22851 =  ( n22484 ) ? ( VREG_11_7 ) : ( n22850 ) ;
assign n22852 =  ( n22483 ) ? ( VREG_11_8 ) : ( n22851 ) ;
assign n22853 =  ( n22482 ) ? ( VREG_11_9 ) : ( n22852 ) ;
assign n22854 =  ( n22481 ) ? ( VREG_11_10 ) : ( n22853 ) ;
assign n22855 =  ( n22480 ) ? ( VREG_11_11 ) : ( n22854 ) ;
assign n22856 =  ( n22479 ) ? ( VREG_11_12 ) : ( n22855 ) ;
assign n22857 =  ( n22478 ) ? ( VREG_11_13 ) : ( n22856 ) ;
assign n22858 =  ( n22477 ) ? ( VREG_11_14 ) : ( n22857 ) ;
assign n22859 =  ( n22476 ) ? ( VREG_11_15 ) : ( n22858 ) ;
assign n22860 =  ( n22475 ) ? ( VREG_12_0 ) : ( n22859 ) ;
assign n22861 =  ( n22474 ) ? ( VREG_12_1 ) : ( n22860 ) ;
assign n22862 =  ( n22473 ) ? ( VREG_12_2 ) : ( n22861 ) ;
assign n22863 =  ( n22472 ) ? ( VREG_12_3 ) : ( n22862 ) ;
assign n22864 =  ( n22471 ) ? ( VREG_12_4 ) : ( n22863 ) ;
assign n22865 =  ( n22470 ) ? ( VREG_12_5 ) : ( n22864 ) ;
assign n22866 =  ( n22469 ) ? ( VREG_12_6 ) : ( n22865 ) ;
assign n22867 =  ( n22468 ) ? ( VREG_12_7 ) : ( n22866 ) ;
assign n22868 =  ( n22467 ) ? ( VREG_12_8 ) : ( n22867 ) ;
assign n22869 =  ( n22466 ) ? ( VREG_12_9 ) : ( n22868 ) ;
assign n22870 =  ( n22465 ) ? ( VREG_12_10 ) : ( n22869 ) ;
assign n22871 =  ( n22464 ) ? ( VREG_12_11 ) : ( n22870 ) ;
assign n22872 =  ( n22463 ) ? ( VREG_12_12 ) : ( n22871 ) ;
assign n22873 =  ( n22462 ) ? ( VREG_12_13 ) : ( n22872 ) ;
assign n22874 =  ( n22461 ) ? ( VREG_12_14 ) : ( n22873 ) ;
assign n22875 =  ( n22460 ) ? ( VREG_12_15 ) : ( n22874 ) ;
assign n22876 =  ( n22459 ) ? ( VREG_13_0 ) : ( n22875 ) ;
assign n22877 =  ( n22458 ) ? ( VREG_13_1 ) : ( n22876 ) ;
assign n22878 =  ( n22457 ) ? ( VREG_13_2 ) : ( n22877 ) ;
assign n22879 =  ( n22456 ) ? ( VREG_13_3 ) : ( n22878 ) ;
assign n22880 =  ( n22455 ) ? ( VREG_13_4 ) : ( n22879 ) ;
assign n22881 =  ( n22454 ) ? ( VREG_13_5 ) : ( n22880 ) ;
assign n22882 =  ( n22453 ) ? ( VREG_13_6 ) : ( n22881 ) ;
assign n22883 =  ( n22452 ) ? ( VREG_13_7 ) : ( n22882 ) ;
assign n22884 =  ( n22451 ) ? ( VREG_13_8 ) : ( n22883 ) ;
assign n22885 =  ( n22450 ) ? ( VREG_13_9 ) : ( n22884 ) ;
assign n22886 =  ( n22449 ) ? ( VREG_13_10 ) : ( n22885 ) ;
assign n22887 =  ( n22448 ) ? ( VREG_13_11 ) : ( n22886 ) ;
assign n22888 =  ( n22447 ) ? ( VREG_13_12 ) : ( n22887 ) ;
assign n22889 =  ( n22446 ) ? ( VREG_13_13 ) : ( n22888 ) ;
assign n22890 =  ( n22445 ) ? ( VREG_13_14 ) : ( n22889 ) ;
assign n22891 =  ( n22444 ) ? ( VREG_13_15 ) : ( n22890 ) ;
assign n22892 =  ( n22443 ) ? ( VREG_14_0 ) : ( n22891 ) ;
assign n22893 =  ( n22442 ) ? ( VREG_14_1 ) : ( n22892 ) ;
assign n22894 =  ( n22441 ) ? ( VREG_14_2 ) : ( n22893 ) ;
assign n22895 =  ( n22440 ) ? ( VREG_14_3 ) : ( n22894 ) ;
assign n22896 =  ( n22439 ) ? ( VREG_14_4 ) : ( n22895 ) ;
assign n22897 =  ( n22438 ) ? ( VREG_14_5 ) : ( n22896 ) ;
assign n22898 =  ( n22437 ) ? ( VREG_14_6 ) : ( n22897 ) ;
assign n22899 =  ( n22436 ) ? ( VREG_14_7 ) : ( n22898 ) ;
assign n22900 =  ( n22435 ) ? ( VREG_14_8 ) : ( n22899 ) ;
assign n22901 =  ( n22434 ) ? ( VREG_14_9 ) : ( n22900 ) ;
assign n22902 =  ( n22433 ) ? ( VREG_14_10 ) : ( n22901 ) ;
assign n22903 =  ( n22432 ) ? ( VREG_14_11 ) : ( n22902 ) ;
assign n22904 =  ( n22431 ) ? ( VREG_14_12 ) : ( n22903 ) ;
assign n22905 =  ( n22430 ) ? ( VREG_14_13 ) : ( n22904 ) ;
assign n22906 =  ( n22429 ) ? ( VREG_14_14 ) : ( n22905 ) ;
assign n22907 =  ( n22428 ) ? ( VREG_14_15 ) : ( n22906 ) ;
assign n22908 =  ( n22427 ) ? ( VREG_15_0 ) : ( n22907 ) ;
assign n22909 =  ( n22426 ) ? ( VREG_15_1 ) : ( n22908 ) ;
assign n22910 =  ( n22425 ) ? ( VREG_15_2 ) : ( n22909 ) ;
assign n22911 =  ( n22424 ) ? ( VREG_15_3 ) : ( n22910 ) ;
assign n22912 =  ( n22423 ) ? ( VREG_15_4 ) : ( n22911 ) ;
assign n22913 =  ( n22422 ) ? ( VREG_15_5 ) : ( n22912 ) ;
assign n22914 =  ( n22421 ) ? ( VREG_15_6 ) : ( n22913 ) ;
assign n22915 =  ( n22420 ) ? ( VREG_15_7 ) : ( n22914 ) ;
assign n22916 =  ( n22419 ) ? ( VREG_15_8 ) : ( n22915 ) ;
assign n22917 =  ( n22418 ) ? ( VREG_15_9 ) : ( n22916 ) ;
assign n22918 =  ( n22417 ) ? ( VREG_15_10 ) : ( n22917 ) ;
assign n22919 =  ( n22416 ) ? ( VREG_15_11 ) : ( n22918 ) ;
assign n22920 =  ( n22415 ) ? ( VREG_15_12 ) : ( n22919 ) ;
assign n22921 =  ( n22414 ) ? ( VREG_15_13 ) : ( n22920 ) ;
assign n22922 =  ( n22413 ) ? ( VREG_15_14 ) : ( n22921 ) ;
assign n22923 =  ( n22412 ) ? ( VREG_15_15 ) : ( n22922 ) ;
assign n22924 =  ( n22411 ) ? ( VREG_16_0 ) : ( n22923 ) ;
assign n22925 =  ( n22410 ) ? ( VREG_16_1 ) : ( n22924 ) ;
assign n22926 =  ( n22409 ) ? ( VREG_16_2 ) : ( n22925 ) ;
assign n22927 =  ( n22408 ) ? ( VREG_16_3 ) : ( n22926 ) ;
assign n22928 =  ( n22407 ) ? ( VREG_16_4 ) : ( n22927 ) ;
assign n22929 =  ( n22406 ) ? ( VREG_16_5 ) : ( n22928 ) ;
assign n22930 =  ( n22405 ) ? ( VREG_16_6 ) : ( n22929 ) ;
assign n22931 =  ( n22404 ) ? ( VREG_16_7 ) : ( n22930 ) ;
assign n22932 =  ( n22403 ) ? ( VREG_16_8 ) : ( n22931 ) ;
assign n22933 =  ( n22402 ) ? ( VREG_16_9 ) : ( n22932 ) ;
assign n22934 =  ( n22401 ) ? ( VREG_16_10 ) : ( n22933 ) ;
assign n22935 =  ( n22400 ) ? ( VREG_16_11 ) : ( n22934 ) ;
assign n22936 =  ( n22399 ) ? ( VREG_16_12 ) : ( n22935 ) ;
assign n22937 =  ( n22398 ) ? ( VREG_16_13 ) : ( n22936 ) ;
assign n22938 =  ( n22397 ) ? ( VREG_16_14 ) : ( n22937 ) ;
assign n22939 =  ( n22396 ) ? ( VREG_16_15 ) : ( n22938 ) ;
assign n22940 =  ( n22395 ) ? ( VREG_17_0 ) : ( n22939 ) ;
assign n22941 =  ( n22394 ) ? ( VREG_17_1 ) : ( n22940 ) ;
assign n22942 =  ( n22393 ) ? ( VREG_17_2 ) : ( n22941 ) ;
assign n22943 =  ( n22392 ) ? ( VREG_17_3 ) : ( n22942 ) ;
assign n22944 =  ( n22391 ) ? ( VREG_17_4 ) : ( n22943 ) ;
assign n22945 =  ( n22390 ) ? ( VREG_17_5 ) : ( n22944 ) ;
assign n22946 =  ( n22389 ) ? ( VREG_17_6 ) : ( n22945 ) ;
assign n22947 =  ( n22388 ) ? ( VREG_17_7 ) : ( n22946 ) ;
assign n22948 =  ( n22387 ) ? ( VREG_17_8 ) : ( n22947 ) ;
assign n22949 =  ( n22386 ) ? ( VREG_17_9 ) : ( n22948 ) ;
assign n22950 =  ( n22385 ) ? ( VREG_17_10 ) : ( n22949 ) ;
assign n22951 =  ( n22384 ) ? ( VREG_17_11 ) : ( n22950 ) ;
assign n22952 =  ( n22383 ) ? ( VREG_17_12 ) : ( n22951 ) ;
assign n22953 =  ( n22382 ) ? ( VREG_17_13 ) : ( n22952 ) ;
assign n22954 =  ( n22381 ) ? ( VREG_17_14 ) : ( n22953 ) ;
assign n22955 =  ( n22380 ) ? ( VREG_17_15 ) : ( n22954 ) ;
assign n22956 =  ( n22379 ) ? ( VREG_18_0 ) : ( n22955 ) ;
assign n22957 =  ( n22378 ) ? ( VREG_18_1 ) : ( n22956 ) ;
assign n22958 =  ( n22377 ) ? ( VREG_18_2 ) : ( n22957 ) ;
assign n22959 =  ( n22376 ) ? ( VREG_18_3 ) : ( n22958 ) ;
assign n22960 =  ( n22375 ) ? ( VREG_18_4 ) : ( n22959 ) ;
assign n22961 =  ( n22374 ) ? ( VREG_18_5 ) : ( n22960 ) ;
assign n22962 =  ( n22373 ) ? ( VREG_18_6 ) : ( n22961 ) ;
assign n22963 =  ( n22372 ) ? ( VREG_18_7 ) : ( n22962 ) ;
assign n22964 =  ( n22371 ) ? ( VREG_18_8 ) : ( n22963 ) ;
assign n22965 =  ( n22370 ) ? ( VREG_18_9 ) : ( n22964 ) ;
assign n22966 =  ( n22369 ) ? ( VREG_18_10 ) : ( n22965 ) ;
assign n22967 =  ( n22368 ) ? ( VREG_18_11 ) : ( n22966 ) ;
assign n22968 =  ( n22367 ) ? ( VREG_18_12 ) : ( n22967 ) ;
assign n22969 =  ( n22366 ) ? ( VREG_18_13 ) : ( n22968 ) ;
assign n22970 =  ( n22365 ) ? ( VREG_18_14 ) : ( n22969 ) ;
assign n22971 =  ( n22364 ) ? ( VREG_18_15 ) : ( n22970 ) ;
assign n22972 =  ( n22363 ) ? ( VREG_19_0 ) : ( n22971 ) ;
assign n22973 =  ( n22362 ) ? ( VREG_19_1 ) : ( n22972 ) ;
assign n22974 =  ( n22361 ) ? ( VREG_19_2 ) : ( n22973 ) ;
assign n22975 =  ( n22360 ) ? ( VREG_19_3 ) : ( n22974 ) ;
assign n22976 =  ( n22359 ) ? ( VREG_19_4 ) : ( n22975 ) ;
assign n22977 =  ( n22358 ) ? ( VREG_19_5 ) : ( n22976 ) ;
assign n22978 =  ( n22357 ) ? ( VREG_19_6 ) : ( n22977 ) ;
assign n22979 =  ( n22356 ) ? ( VREG_19_7 ) : ( n22978 ) ;
assign n22980 =  ( n22355 ) ? ( VREG_19_8 ) : ( n22979 ) ;
assign n22981 =  ( n22354 ) ? ( VREG_19_9 ) : ( n22980 ) ;
assign n22982 =  ( n22353 ) ? ( VREG_19_10 ) : ( n22981 ) ;
assign n22983 =  ( n22352 ) ? ( VREG_19_11 ) : ( n22982 ) ;
assign n22984 =  ( n22351 ) ? ( VREG_19_12 ) : ( n22983 ) ;
assign n22985 =  ( n22350 ) ? ( VREG_19_13 ) : ( n22984 ) ;
assign n22986 =  ( n22349 ) ? ( VREG_19_14 ) : ( n22985 ) ;
assign n22987 =  ( n22348 ) ? ( VREG_19_15 ) : ( n22986 ) ;
assign n22988 =  ( n22347 ) ? ( VREG_20_0 ) : ( n22987 ) ;
assign n22989 =  ( n22346 ) ? ( VREG_20_1 ) : ( n22988 ) ;
assign n22990 =  ( n22345 ) ? ( VREG_20_2 ) : ( n22989 ) ;
assign n22991 =  ( n22344 ) ? ( VREG_20_3 ) : ( n22990 ) ;
assign n22992 =  ( n22343 ) ? ( VREG_20_4 ) : ( n22991 ) ;
assign n22993 =  ( n22342 ) ? ( VREG_20_5 ) : ( n22992 ) ;
assign n22994 =  ( n22341 ) ? ( VREG_20_6 ) : ( n22993 ) ;
assign n22995 =  ( n22340 ) ? ( VREG_20_7 ) : ( n22994 ) ;
assign n22996 =  ( n22339 ) ? ( VREG_20_8 ) : ( n22995 ) ;
assign n22997 =  ( n22338 ) ? ( VREG_20_9 ) : ( n22996 ) ;
assign n22998 =  ( n22337 ) ? ( VREG_20_10 ) : ( n22997 ) ;
assign n22999 =  ( n22336 ) ? ( VREG_20_11 ) : ( n22998 ) ;
assign n23000 =  ( n22335 ) ? ( VREG_20_12 ) : ( n22999 ) ;
assign n23001 =  ( n22334 ) ? ( VREG_20_13 ) : ( n23000 ) ;
assign n23002 =  ( n22333 ) ? ( VREG_20_14 ) : ( n23001 ) ;
assign n23003 =  ( n22332 ) ? ( VREG_20_15 ) : ( n23002 ) ;
assign n23004 =  ( n22331 ) ? ( VREG_21_0 ) : ( n23003 ) ;
assign n23005 =  ( n22330 ) ? ( VREG_21_1 ) : ( n23004 ) ;
assign n23006 =  ( n22329 ) ? ( VREG_21_2 ) : ( n23005 ) ;
assign n23007 =  ( n22328 ) ? ( VREG_21_3 ) : ( n23006 ) ;
assign n23008 =  ( n22327 ) ? ( VREG_21_4 ) : ( n23007 ) ;
assign n23009 =  ( n22326 ) ? ( VREG_21_5 ) : ( n23008 ) ;
assign n23010 =  ( n22325 ) ? ( VREG_21_6 ) : ( n23009 ) ;
assign n23011 =  ( n22324 ) ? ( VREG_21_7 ) : ( n23010 ) ;
assign n23012 =  ( n22323 ) ? ( VREG_21_8 ) : ( n23011 ) ;
assign n23013 =  ( n22322 ) ? ( VREG_21_9 ) : ( n23012 ) ;
assign n23014 =  ( n22321 ) ? ( VREG_21_10 ) : ( n23013 ) ;
assign n23015 =  ( n22320 ) ? ( VREG_21_11 ) : ( n23014 ) ;
assign n23016 =  ( n22319 ) ? ( VREG_21_12 ) : ( n23015 ) ;
assign n23017 =  ( n22318 ) ? ( VREG_21_13 ) : ( n23016 ) ;
assign n23018 =  ( n22317 ) ? ( VREG_21_14 ) : ( n23017 ) ;
assign n23019 =  ( n22316 ) ? ( VREG_21_15 ) : ( n23018 ) ;
assign n23020 =  ( n22315 ) ? ( VREG_22_0 ) : ( n23019 ) ;
assign n23021 =  ( n22314 ) ? ( VREG_22_1 ) : ( n23020 ) ;
assign n23022 =  ( n22313 ) ? ( VREG_22_2 ) : ( n23021 ) ;
assign n23023 =  ( n22312 ) ? ( VREG_22_3 ) : ( n23022 ) ;
assign n23024 =  ( n22311 ) ? ( VREG_22_4 ) : ( n23023 ) ;
assign n23025 =  ( n22310 ) ? ( VREG_22_5 ) : ( n23024 ) ;
assign n23026 =  ( n22309 ) ? ( VREG_22_6 ) : ( n23025 ) ;
assign n23027 =  ( n22308 ) ? ( VREG_22_7 ) : ( n23026 ) ;
assign n23028 =  ( n22307 ) ? ( VREG_22_8 ) : ( n23027 ) ;
assign n23029 =  ( n22306 ) ? ( VREG_22_9 ) : ( n23028 ) ;
assign n23030 =  ( n22305 ) ? ( VREG_22_10 ) : ( n23029 ) ;
assign n23031 =  ( n22304 ) ? ( VREG_22_11 ) : ( n23030 ) ;
assign n23032 =  ( n22303 ) ? ( VREG_22_12 ) : ( n23031 ) ;
assign n23033 =  ( n22302 ) ? ( VREG_22_13 ) : ( n23032 ) ;
assign n23034 =  ( n22301 ) ? ( VREG_22_14 ) : ( n23033 ) ;
assign n23035 =  ( n22300 ) ? ( VREG_22_15 ) : ( n23034 ) ;
assign n23036 =  ( n22299 ) ? ( VREG_23_0 ) : ( n23035 ) ;
assign n23037 =  ( n22298 ) ? ( VREG_23_1 ) : ( n23036 ) ;
assign n23038 =  ( n22297 ) ? ( VREG_23_2 ) : ( n23037 ) ;
assign n23039 =  ( n22296 ) ? ( VREG_23_3 ) : ( n23038 ) ;
assign n23040 =  ( n22295 ) ? ( VREG_23_4 ) : ( n23039 ) ;
assign n23041 =  ( n22294 ) ? ( VREG_23_5 ) : ( n23040 ) ;
assign n23042 =  ( n22293 ) ? ( VREG_23_6 ) : ( n23041 ) ;
assign n23043 =  ( n22292 ) ? ( VREG_23_7 ) : ( n23042 ) ;
assign n23044 =  ( n22291 ) ? ( VREG_23_8 ) : ( n23043 ) ;
assign n23045 =  ( n22290 ) ? ( VREG_23_9 ) : ( n23044 ) ;
assign n23046 =  ( n22289 ) ? ( VREG_23_10 ) : ( n23045 ) ;
assign n23047 =  ( n22288 ) ? ( VREG_23_11 ) : ( n23046 ) ;
assign n23048 =  ( n22287 ) ? ( VREG_23_12 ) : ( n23047 ) ;
assign n23049 =  ( n22286 ) ? ( VREG_23_13 ) : ( n23048 ) ;
assign n23050 =  ( n22285 ) ? ( VREG_23_14 ) : ( n23049 ) ;
assign n23051 =  ( n22284 ) ? ( VREG_23_15 ) : ( n23050 ) ;
assign n23052 =  ( n22283 ) ? ( VREG_24_0 ) : ( n23051 ) ;
assign n23053 =  ( n22282 ) ? ( VREG_24_1 ) : ( n23052 ) ;
assign n23054 =  ( n22281 ) ? ( VREG_24_2 ) : ( n23053 ) ;
assign n23055 =  ( n22280 ) ? ( VREG_24_3 ) : ( n23054 ) ;
assign n23056 =  ( n22279 ) ? ( VREG_24_4 ) : ( n23055 ) ;
assign n23057 =  ( n22278 ) ? ( VREG_24_5 ) : ( n23056 ) ;
assign n23058 =  ( n22277 ) ? ( VREG_24_6 ) : ( n23057 ) ;
assign n23059 =  ( n22276 ) ? ( VREG_24_7 ) : ( n23058 ) ;
assign n23060 =  ( n22275 ) ? ( VREG_24_8 ) : ( n23059 ) ;
assign n23061 =  ( n22274 ) ? ( VREG_24_9 ) : ( n23060 ) ;
assign n23062 =  ( n22273 ) ? ( VREG_24_10 ) : ( n23061 ) ;
assign n23063 =  ( n22272 ) ? ( VREG_24_11 ) : ( n23062 ) ;
assign n23064 =  ( n22271 ) ? ( VREG_24_12 ) : ( n23063 ) ;
assign n23065 =  ( n22270 ) ? ( VREG_24_13 ) : ( n23064 ) ;
assign n23066 =  ( n22269 ) ? ( VREG_24_14 ) : ( n23065 ) ;
assign n23067 =  ( n22268 ) ? ( VREG_24_15 ) : ( n23066 ) ;
assign n23068 =  ( n22267 ) ? ( VREG_25_0 ) : ( n23067 ) ;
assign n23069 =  ( n22266 ) ? ( VREG_25_1 ) : ( n23068 ) ;
assign n23070 =  ( n22265 ) ? ( VREG_25_2 ) : ( n23069 ) ;
assign n23071 =  ( n22264 ) ? ( VREG_25_3 ) : ( n23070 ) ;
assign n23072 =  ( n22263 ) ? ( VREG_25_4 ) : ( n23071 ) ;
assign n23073 =  ( n22262 ) ? ( VREG_25_5 ) : ( n23072 ) ;
assign n23074 =  ( n22261 ) ? ( VREG_25_6 ) : ( n23073 ) ;
assign n23075 =  ( n22260 ) ? ( VREG_25_7 ) : ( n23074 ) ;
assign n23076 =  ( n22259 ) ? ( VREG_25_8 ) : ( n23075 ) ;
assign n23077 =  ( n22258 ) ? ( VREG_25_9 ) : ( n23076 ) ;
assign n23078 =  ( n22257 ) ? ( VREG_25_10 ) : ( n23077 ) ;
assign n23079 =  ( n22256 ) ? ( VREG_25_11 ) : ( n23078 ) ;
assign n23080 =  ( n22255 ) ? ( VREG_25_12 ) : ( n23079 ) ;
assign n23081 =  ( n22254 ) ? ( VREG_25_13 ) : ( n23080 ) ;
assign n23082 =  ( n22253 ) ? ( VREG_25_14 ) : ( n23081 ) ;
assign n23083 =  ( n22252 ) ? ( VREG_25_15 ) : ( n23082 ) ;
assign n23084 =  ( n22251 ) ? ( VREG_26_0 ) : ( n23083 ) ;
assign n23085 =  ( n22250 ) ? ( VREG_26_1 ) : ( n23084 ) ;
assign n23086 =  ( n22249 ) ? ( VREG_26_2 ) : ( n23085 ) ;
assign n23087 =  ( n22248 ) ? ( VREG_26_3 ) : ( n23086 ) ;
assign n23088 =  ( n22247 ) ? ( VREG_26_4 ) : ( n23087 ) ;
assign n23089 =  ( n22246 ) ? ( VREG_26_5 ) : ( n23088 ) ;
assign n23090 =  ( n22245 ) ? ( VREG_26_6 ) : ( n23089 ) ;
assign n23091 =  ( n22244 ) ? ( VREG_26_7 ) : ( n23090 ) ;
assign n23092 =  ( n22243 ) ? ( VREG_26_8 ) : ( n23091 ) ;
assign n23093 =  ( n22242 ) ? ( VREG_26_9 ) : ( n23092 ) ;
assign n23094 =  ( n22241 ) ? ( VREG_26_10 ) : ( n23093 ) ;
assign n23095 =  ( n22240 ) ? ( VREG_26_11 ) : ( n23094 ) ;
assign n23096 =  ( n22239 ) ? ( VREG_26_12 ) : ( n23095 ) ;
assign n23097 =  ( n22238 ) ? ( VREG_26_13 ) : ( n23096 ) ;
assign n23098 =  ( n22237 ) ? ( VREG_26_14 ) : ( n23097 ) ;
assign n23099 =  ( n22236 ) ? ( VREG_26_15 ) : ( n23098 ) ;
assign n23100 =  ( n22235 ) ? ( VREG_27_0 ) : ( n23099 ) ;
assign n23101 =  ( n22234 ) ? ( VREG_27_1 ) : ( n23100 ) ;
assign n23102 =  ( n22233 ) ? ( VREG_27_2 ) : ( n23101 ) ;
assign n23103 =  ( n22232 ) ? ( VREG_27_3 ) : ( n23102 ) ;
assign n23104 =  ( n22231 ) ? ( VREG_27_4 ) : ( n23103 ) ;
assign n23105 =  ( n22230 ) ? ( VREG_27_5 ) : ( n23104 ) ;
assign n23106 =  ( n22229 ) ? ( VREG_27_6 ) : ( n23105 ) ;
assign n23107 =  ( n22228 ) ? ( VREG_27_7 ) : ( n23106 ) ;
assign n23108 =  ( n22227 ) ? ( VREG_27_8 ) : ( n23107 ) ;
assign n23109 =  ( n22226 ) ? ( VREG_27_9 ) : ( n23108 ) ;
assign n23110 =  ( n22225 ) ? ( VREG_27_10 ) : ( n23109 ) ;
assign n23111 =  ( n22224 ) ? ( VREG_27_11 ) : ( n23110 ) ;
assign n23112 =  ( n22223 ) ? ( VREG_27_12 ) : ( n23111 ) ;
assign n23113 =  ( n22222 ) ? ( VREG_27_13 ) : ( n23112 ) ;
assign n23114 =  ( n22221 ) ? ( VREG_27_14 ) : ( n23113 ) ;
assign n23115 =  ( n22220 ) ? ( VREG_27_15 ) : ( n23114 ) ;
assign n23116 =  ( n22219 ) ? ( VREG_28_0 ) : ( n23115 ) ;
assign n23117 =  ( n22218 ) ? ( VREG_28_1 ) : ( n23116 ) ;
assign n23118 =  ( n22217 ) ? ( VREG_28_2 ) : ( n23117 ) ;
assign n23119 =  ( n22216 ) ? ( VREG_28_3 ) : ( n23118 ) ;
assign n23120 =  ( n22215 ) ? ( VREG_28_4 ) : ( n23119 ) ;
assign n23121 =  ( n22214 ) ? ( VREG_28_5 ) : ( n23120 ) ;
assign n23122 =  ( n22213 ) ? ( VREG_28_6 ) : ( n23121 ) ;
assign n23123 =  ( n22212 ) ? ( VREG_28_7 ) : ( n23122 ) ;
assign n23124 =  ( n22211 ) ? ( VREG_28_8 ) : ( n23123 ) ;
assign n23125 =  ( n22210 ) ? ( VREG_28_9 ) : ( n23124 ) ;
assign n23126 =  ( n22209 ) ? ( VREG_28_10 ) : ( n23125 ) ;
assign n23127 =  ( n22208 ) ? ( VREG_28_11 ) : ( n23126 ) ;
assign n23128 =  ( n22207 ) ? ( VREG_28_12 ) : ( n23127 ) ;
assign n23129 =  ( n22206 ) ? ( VREG_28_13 ) : ( n23128 ) ;
assign n23130 =  ( n22205 ) ? ( VREG_28_14 ) : ( n23129 ) ;
assign n23131 =  ( n22204 ) ? ( VREG_28_15 ) : ( n23130 ) ;
assign n23132 =  ( n22203 ) ? ( VREG_29_0 ) : ( n23131 ) ;
assign n23133 =  ( n22202 ) ? ( VREG_29_1 ) : ( n23132 ) ;
assign n23134 =  ( n22201 ) ? ( VREG_29_2 ) : ( n23133 ) ;
assign n23135 =  ( n22200 ) ? ( VREG_29_3 ) : ( n23134 ) ;
assign n23136 =  ( n22199 ) ? ( VREG_29_4 ) : ( n23135 ) ;
assign n23137 =  ( n22198 ) ? ( VREG_29_5 ) : ( n23136 ) ;
assign n23138 =  ( n22197 ) ? ( VREG_29_6 ) : ( n23137 ) ;
assign n23139 =  ( n22196 ) ? ( VREG_29_7 ) : ( n23138 ) ;
assign n23140 =  ( n22195 ) ? ( VREG_29_8 ) : ( n23139 ) ;
assign n23141 =  ( n22194 ) ? ( VREG_29_9 ) : ( n23140 ) ;
assign n23142 =  ( n22193 ) ? ( VREG_29_10 ) : ( n23141 ) ;
assign n23143 =  ( n22192 ) ? ( VREG_29_11 ) : ( n23142 ) ;
assign n23144 =  ( n22191 ) ? ( VREG_29_12 ) : ( n23143 ) ;
assign n23145 =  ( n22190 ) ? ( VREG_29_13 ) : ( n23144 ) ;
assign n23146 =  ( n22189 ) ? ( VREG_29_14 ) : ( n23145 ) ;
assign n23147 =  ( n22188 ) ? ( VREG_29_15 ) : ( n23146 ) ;
assign n23148 =  ( n22187 ) ? ( VREG_30_0 ) : ( n23147 ) ;
assign n23149 =  ( n22186 ) ? ( VREG_30_1 ) : ( n23148 ) ;
assign n23150 =  ( n22185 ) ? ( VREG_30_2 ) : ( n23149 ) ;
assign n23151 =  ( n22184 ) ? ( VREG_30_3 ) : ( n23150 ) ;
assign n23152 =  ( n22183 ) ? ( VREG_30_4 ) : ( n23151 ) ;
assign n23153 =  ( n22182 ) ? ( VREG_30_5 ) : ( n23152 ) ;
assign n23154 =  ( n22181 ) ? ( VREG_30_6 ) : ( n23153 ) ;
assign n23155 =  ( n22180 ) ? ( VREG_30_7 ) : ( n23154 ) ;
assign n23156 =  ( n22179 ) ? ( VREG_30_8 ) : ( n23155 ) ;
assign n23157 =  ( n22178 ) ? ( VREG_30_9 ) : ( n23156 ) ;
assign n23158 =  ( n22177 ) ? ( VREG_30_10 ) : ( n23157 ) ;
assign n23159 =  ( n22176 ) ? ( VREG_30_11 ) : ( n23158 ) ;
assign n23160 =  ( n22175 ) ? ( VREG_30_12 ) : ( n23159 ) ;
assign n23161 =  ( n22174 ) ? ( VREG_30_13 ) : ( n23160 ) ;
assign n23162 =  ( n22173 ) ? ( VREG_30_14 ) : ( n23161 ) ;
assign n23163 =  ( n22172 ) ? ( VREG_30_15 ) : ( n23162 ) ;
assign n23164 =  ( n22171 ) ? ( VREG_31_0 ) : ( n23163 ) ;
assign n23165 =  ( n22169 ) ? ( VREG_31_1 ) : ( n23164 ) ;
assign n23166 =  ( n22167 ) ? ( VREG_31_2 ) : ( n23165 ) ;
assign n23167 =  ( n22165 ) ? ( VREG_31_3 ) : ( n23166 ) ;
assign n23168 =  ( n22163 ) ? ( VREG_31_4 ) : ( n23167 ) ;
assign n23169 =  ( n22161 ) ? ( VREG_31_5 ) : ( n23168 ) ;
assign n23170 =  ( n22159 ) ? ( VREG_31_6 ) : ( n23169 ) ;
assign n23171 =  ( n22157 ) ? ( VREG_31_7 ) : ( n23170 ) ;
assign n23172 =  ( n22155 ) ? ( VREG_31_8 ) : ( n23171 ) ;
assign n23173 =  ( n22153 ) ? ( VREG_31_9 ) : ( n23172 ) ;
assign n23174 =  ( n22151 ) ? ( VREG_31_10 ) : ( n23173 ) ;
assign n23175 =  ( n22149 ) ? ( VREG_31_11 ) : ( n23174 ) ;
assign n23176 =  ( n22147 ) ? ( VREG_31_12 ) : ( n23175 ) ;
assign n23177 =  ( n22145 ) ? ( VREG_31_13 ) : ( n23176 ) ;
assign n23178 =  ( n22143 ) ? ( VREG_31_14 ) : ( n23177 ) ;
assign n23179 =  ( n22141 ) ? ( VREG_31_15 ) : ( n23178 ) ;
assign n23180 =  ( n23179 ) + ( n140 )  ;
assign n23181 =  ( n23179 ) - ( n140 )  ;
assign n23182 =  ( n23179 ) & ( n140 )  ;
assign n23183 =  ( n23179 ) | ( n140 )  ;
assign n23184 =  ( ( n23179 ) * ( n140 ))  ;
assign n23185 =  ( n148 ) ? ( n23184 ) : ( VREG_0_4 ) ;
assign n23186 =  ( n146 ) ? ( n23183 ) : ( n23185 ) ;
assign n23187 =  ( n144 ) ? ( n23182 ) : ( n23186 ) ;
assign n23188 =  ( n142 ) ? ( n23181 ) : ( n23187 ) ;
assign n23189 =  ( n10 ) ? ( n23180 ) : ( n23188 ) ;
assign n23190 =  ( n77 ) & ( n22140 )  ;
assign n23191 =  ( n77 ) & ( n22142 )  ;
assign n23192 =  ( n77 ) & ( n22144 )  ;
assign n23193 =  ( n77 ) & ( n22146 )  ;
assign n23194 =  ( n77 ) & ( n22148 )  ;
assign n23195 =  ( n77 ) & ( n22150 )  ;
assign n23196 =  ( n77 ) & ( n22152 )  ;
assign n23197 =  ( n77 ) & ( n22154 )  ;
assign n23198 =  ( n77 ) & ( n22156 )  ;
assign n23199 =  ( n77 ) & ( n22158 )  ;
assign n23200 =  ( n77 ) & ( n22160 )  ;
assign n23201 =  ( n77 ) & ( n22162 )  ;
assign n23202 =  ( n77 ) & ( n22164 )  ;
assign n23203 =  ( n77 ) & ( n22166 )  ;
assign n23204 =  ( n77 ) & ( n22168 )  ;
assign n23205 =  ( n77 ) & ( n22170 )  ;
assign n23206 =  ( n78 ) & ( n22140 )  ;
assign n23207 =  ( n78 ) & ( n22142 )  ;
assign n23208 =  ( n78 ) & ( n22144 )  ;
assign n23209 =  ( n78 ) & ( n22146 )  ;
assign n23210 =  ( n78 ) & ( n22148 )  ;
assign n23211 =  ( n78 ) & ( n22150 )  ;
assign n23212 =  ( n78 ) & ( n22152 )  ;
assign n23213 =  ( n78 ) & ( n22154 )  ;
assign n23214 =  ( n78 ) & ( n22156 )  ;
assign n23215 =  ( n78 ) & ( n22158 )  ;
assign n23216 =  ( n78 ) & ( n22160 )  ;
assign n23217 =  ( n78 ) & ( n22162 )  ;
assign n23218 =  ( n78 ) & ( n22164 )  ;
assign n23219 =  ( n78 ) & ( n22166 )  ;
assign n23220 =  ( n78 ) & ( n22168 )  ;
assign n23221 =  ( n78 ) & ( n22170 )  ;
assign n23222 =  ( n79 ) & ( n22140 )  ;
assign n23223 =  ( n79 ) & ( n22142 )  ;
assign n23224 =  ( n79 ) & ( n22144 )  ;
assign n23225 =  ( n79 ) & ( n22146 )  ;
assign n23226 =  ( n79 ) & ( n22148 )  ;
assign n23227 =  ( n79 ) & ( n22150 )  ;
assign n23228 =  ( n79 ) & ( n22152 )  ;
assign n23229 =  ( n79 ) & ( n22154 )  ;
assign n23230 =  ( n79 ) & ( n22156 )  ;
assign n23231 =  ( n79 ) & ( n22158 )  ;
assign n23232 =  ( n79 ) & ( n22160 )  ;
assign n23233 =  ( n79 ) & ( n22162 )  ;
assign n23234 =  ( n79 ) & ( n22164 )  ;
assign n23235 =  ( n79 ) & ( n22166 )  ;
assign n23236 =  ( n79 ) & ( n22168 )  ;
assign n23237 =  ( n79 ) & ( n22170 )  ;
assign n23238 =  ( n80 ) & ( n22140 )  ;
assign n23239 =  ( n80 ) & ( n22142 )  ;
assign n23240 =  ( n80 ) & ( n22144 )  ;
assign n23241 =  ( n80 ) & ( n22146 )  ;
assign n23242 =  ( n80 ) & ( n22148 )  ;
assign n23243 =  ( n80 ) & ( n22150 )  ;
assign n23244 =  ( n80 ) & ( n22152 )  ;
assign n23245 =  ( n80 ) & ( n22154 )  ;
assign n23246 =  ( n80 ) & ( n22156 )  ;
assign n23247 =  ( n80 ) & ( n22158 )  ;
assign n23248 =  ( n80 ) & ( n22160 )  ;
assign n23249 =  ( n80 ) & ( n22162 )  ;
assign n23250 =  ( n80 ) & ( n22164 )  ;
assign n23251 =  ( n80 ) & ( n22166 )  ;
assign n23252 =  ( n80 ) & ( n22168 )  ;
assign n23253 =  ( n80 ) & ( n22170 )  ;
assign n23254 =  ( n81 ) & ( n22140 )  ;
assign n23255 =  ( n81 ) & ( n22142 )  ;
assign n23256 =  ( n81 ) & ( n22144 )  ;
assign n23257 =  ( n81 ) & ( n22146 )  ;
assign n23258 =  ( n81 ) & ( n22148 )  ;
assign n23259 =  ( n81 ) & ( n22150 )  ;
assign n23260 =  ( n81 ) & ( n22152 )  ;
assign n23261 =  ( n81 ) & ( n22154 )  ;
assign n23262 =  ( n81 ) & ( n22156 )  ;
assign n23263 =  ( n81 ) & ( n22158 )  ;
assign n23264 =  ( n81 ) & ( n22160 )  ;
assign n23265 =  ( n81 ) & ( n22162 )  ;
assign n23266 =  ( n81 ) & ( n22164 )  ;
assign n23267 =  ( n81 ) & ( n22166 )  ;
assign n23268 =  ( n81 ) & ( n22168 )  ;
assign n23269 =  ( n81 ) & ( n22170 )  ;
assign n23270 =  ( n82 ) & ( n22140 )  ;
assign n23271 =  ( n82 ) & ( n22142 )  ;
assign n23272 =  ( n82 ) & ( n22144 )  ;
assign n23273 =  ( n82 ) & ( n22146 )  ;
assign n23274 =  ( n82 ) & ( n22148 )  ;
assign n23275 =  ( n82 ) & ( n22150 )  ;
assign n23276 =  ( n82 ) & ( n22152 )  ;
assign n23277 =  ( n82 ) & ( n22154 )  ;
assign n23278 =  ( n82 ) & ( n22156 )  ;
assign n23279 =  ( n82 ) & ( n22158 )  ;
assign n23280 =  ( n82 ) & ( n22160 )  ;
assign n23281 =  ( n82 ) & ( n22162 )  ;
assign n23282 =  ( n82 ) & ( n22164 )  ;
assign n23283 =  ( n82 ) & ( n22166 )  ;
assign n23284 =  ( n82 ) & ( n22168 )  ;
assign n23285 =  ( n82 ) & ( n22170 )  ;
assign n23286 =  ( n83 ) & ( n22140 )  ;
assign n23287 =  ( n83 ) & ( n22142 )  ;
assign n23288 =  ( n83 ) & ( n22144 )  ;
assign n23289 =  ( n83 ) & ( n22146 )  ;
assign n23290 =  ( n83 ) & ( n22148 )  ;
assign n23291 =  ( n83 ) & ( n22150 )  ;
assign n23292 =  ( n83 ) & ( n22152 )  ;
assign n23293 =  ( n83 ) & ( n22154 )  ;
assign n23294 =  ( n83 ) & ( n22156 )  ;
assign n23295 =  ( n83 ) & ( n22158 )  ;
assign n23296 =  ( n83 ) & ( n22160 )  ;
assign n23297 =  ( n83 ) & ( n22162 )  ;
assign n23298 =  ( n83 ) & ( n22164 )  ;
assign n23299 =  ( n83 ) & ( n22166 )  ;
assign n23300 =  ( n83 ) & ( n22168 )  ;
assign n23301 =  ( n83 ) & ( n22170 )  ;
assign n23302 =  ( n84 ) & ( n22140 )  ;
assign n23303 =  ( n84 ) & ( n22142 )  ;
assign n23304 =  ( n84 ) & ( n22144 )  ;
assign n23305 =  ( n84 ) & ( n22146 )  ;
assign n23306 =  ( n84 ) & ( n22148 )  ;
assign n23307 =  ( n84 ) & ( n22150 )  ;
assign n23308 =  ( n84 ) & ( n22152 )  ;
assign n23309 =  ( n84 ) & ( n22154 )  ;
assign n23310 =  ( n84 ) & ( n22156 )  ;
assign n23311 =  ( n84 ) & ( n22158 )  ;
assign n23312 =  ( n84 ) & ( n22160 )  ;
assign n23313 =  ( n84 ) & ( n22162 )  ;
assign n23314 =  ( n84 ) & ( n22164 )  ;
assign n23315 =  ( n84 ) & ( n22166 )  ;
assign n23316 =  ( n84 ) & ( n22168 )  ;
assign n23317 =  ( n84 ) & ( n22170 )  ;
assign n23318 =  ( n85 ) & ( n22140 )  ;
assign n23319 =  ( n85 ) & ( n22142 )  ;
assign n23320 =  ( n85 ) & ( n22144 )  ;
assign n23321 =  ( n85 ) & ( n22146 )  ;
assign n23322 =  ( n85 ) & ( n22148 )  ;
assign n23323 =  ( n85 ) & ( n22150 )  ;
assign n23324 =  ( n85 ) & ( n22152 )  ;
assign n23325 =  ( n85 ) & ( n22154 )  ;
assign n23326 =  ( n85 ) & ( n22156 )  ;
assign n23327 =  ( n85 ) & ( n22158 )  ;
assign n23328 =  ( n85 ) & ( n22160 )  ;
assign n23329 =  ( n85 ) & ( n22162 )  ;
assign n23330 =  ( n85 ) & ( n22164 )  ;
assign n23331 =  ( n85 ) & ( n22166 )  ;
assign n23332 =  ( n85 ) & ( n22168 )  ;
assign n23333 =  ( n85 ) & ( n22170 )  ;
assign n23334 =  ( n86 ) & ( n22140 )  ;
assign n23335 =  ( n86 ) & ( n22142 )  ;
assign n23336 =  ( n86 ) & ( n22144 )  ;
assign n23337 =  ( n86 ) & ( n22146 )  ;
assign n23338 =  ( n86 ) & ( n22148 )  ;
assign n23339 =  ( n86 ) & ( n22150 )  ;
assign n23340 =  ( n86 ) & ( n22152 )  ;
assign n23341 =  ( n86 ) & ( n22154 )  ;
assign n23342 =  ( n86 ) & ( n22156 )  ;
assign n23343 =  ( n86 ) & ( n22158 )  ;
assign n23344 =  ( n86 ) & ( n22160 )  ;
assign n23345 =  ( n86 ) & ( n22162 )  ;
assign n23346 =  ( n86 ) & ( n22164 )  ;
assign n23347 =  ( n86 ) & ( n22166 )  ;
assign n23348 =  ( n86 ) & ( n22168 )  ;
assign n23349 =  ( n86 ) & ( n22170 )  ;
assign n23350 =  ( n87 ) & ( n22140 )  ;
assign n23351 =  ( n87 ) & ( n22142 )  ;
assign n23352 =  ( n87 ) & ( n22144 )  ;
assign n23353 =  ( n87 ) & ( n22146 )  ;
assign n23354 =  ( n87 ) & ( n22148 )  ;
assign n23355 =  ( n87 ) & ( n22150 )  ;
assign n23356 =  ( n87 ) & ( n22152 )  ;
assign n23357 =  ( n87 ) & ( n22154 )  ;
assign n23358 =  ( n87 ) & ( n22156 )  ;
assign n23359 =  ( n87 ) & ( n22158 )  ;
assign n23360 =  ( n87 ) & ( n22160 )  ;
assign n23361 =  ( n87 ) & ( n22162 )  ;
assign n23362 =  ( n87 ) & ( n22164 )  ;
assign n23363 =  ( n87 ) & ( n22166 )  ;
assign n23364 =  ( n87 ) & ( n22168 )  ;
assign n23365 =  ( n87 ) & ( n22170 )  ;
assign n23366 =  ( n88 ) & ( n22140 )  ;
assign n23367 =  ( n88 ) & ( n22142 )  ;
assign n23368 =  ( n88 ) & ( n22144 )  ;
assign n23369 =  ( n88 ) & ( n22146 )  ;
assign n23370 =  ( n88 ) & ( n22148 )  ;
assign n23371 =  ( n88 ) & ( n22150 )  ;
assign n23372 =  ( n88 ) & ( n22152 )  ;
assign n23373 =  ( n88 ) & ( n22154 )  ;
assign n23374 =  ( n88 ) & ( n22156 )  ;
assign n23375 =  ( n88 ) & ( n22158 )  ;
assign n23376 =  ( n88 ) & ( n22160 )  ;
assign n23377 =  ( n88 ) & ( n22162 )  ;
assign n23378 =  ( n88 ) & ( n22164 )  ;
assign n23379 =  ( n88 ) & ( n22166 )  ;
assign n23380 =  ( n88 ) & ( n22168 )  ;
assign n23381 =  ( n88 ) & ( n22170 )  ;
assign n23382 =  ( n89 ) & ( n22140 )  ;
assign n23383 =  ( n89 ) & ( n22142 )  ;
assign n23384 =  ( n89 ) & ( n22144 )  ;
assign n23385 =  ( n89 ) & ( n22146 )  ;
assign n23386 =  ( n89 ) & ( n22148 )  ;
assign n23387 =  ( n89 ) & ( n22150 )  ;
assign n23388 =  ( n89 ) & ( n22152 )  ;
assign n23389 =  ( n89 ) & ( n22154 )  ;
assign n23390 =  ( n89 ) & ( n22156 )  ;
assign n23391 =  ( n89 ) & ( n22158 )  ;
assign n23392 =  ( n89 ) & ( n22160 )  ;
assign n23393 =  ( n89 ) & ( n22162 )  ;
assign n23394 =  ( n89 ) & ( n22164 )  ;
assign n23395 =  ( n89 ) & ( n22166 )  ;
assign n23396 =  ( n89 ) & ( n22168 )  ;
assign n23397 =  ( n89 ) & ( n22170 )  ;
assign n23398 =  ( n90 ) & ( n22140 )  ;
assign n23399 =  ( n90 ) & ( n22142 )  ;
assign n23400 =  ( n90 ) & ( n22144 )  ;
assign n23401 =  ( n90 ) & ( n22146 )  ;
assign n23402 =  ( n90 ) & ( n22148 )  ;
assign n23403 =  ( n90 ) & ( n22150 )  ;
assign n23404 =  ( n90 ) & ( n22152 )  ;
assign n23405 =  ( n90 ) & ( n22154 )  ;
assign n23406 =  ( n90 ) & ( n22156 )  ;
assign n23407 =  ( n90 ) & ( n22158 )  ;
assign n23408 =  ( n90 ) & ( n22160 )  ;
assign n23409 =  ( n90 ) & ( n22162 )  ;
assign n23410 =  ( n90 ) & ( n22164 )  ;
assign n23411 =  ( n90 ) & ( n22166 )  ;
assign n23412 =  ( n90 ) & ( n22168 )  ;
assign n23413 =  ( n90 ) & ( n22170 )  ;
assign n23414 =  ( n91 ) & ( n22140 )  ;
assign n23415 =  ( n91 ) & ( n22142 )  ;
assign n23416 =  ( n91 ) & ( n22144 )  ;
assign n23417 =  ( n91 ) & ( n22146 )  ;
assign n23418 =  ( n91 ) & ( n22148 )  ;
assign n23419 =  ( n91 ) & ( n22150 )  ;
assign n23420 =  ( n91 ) & ( n22152 )  ;
assign n23421 =  ( n91 ) & ( n22154 )  ;
assign n23422 =  ( n91 ) & ( n22156 )  ;
assign n23423 =  ( n91 ) & ( n22158 )  ;
assign n23424 =  ( n91 ) & ( n22160 )  ;
assign n23425 =  ( n91 ) & ( n22162 )  ;
assign n23426 =  ( n91 ) & ( n22164 )  ;
assign n23427 =  ( n91 ) & ( n22166 )  ;
assign n23428 =  ( n91 ) & ( n22168 )  ;
assign n23429 =  ( n91 ) & ( n22170 )  ;
assign n23430 =  ( n92 ) & ( n22140 )  ;
assign n23431 =  ( n92 ) & ( n22142 )  ;
assign n23432 =  ( n92 ) & ( n22144 )  ;
assign n23433 =  ( n92 ) & ( n22146 )  ;
assign n23434 =  ( n92 ) & ( n22148 )  ;
assign n23435 =  ( n92 ) & ( n22150 )  ;
assign n23436 =  ( n92 ) & ( n22152 )  ;
assign n23437 =  ( n92 ) & ( n22154 )  ;
assign n23438 =  ( n92 ) & ( n22156 )  ;
assign n23439 =  ( n92 ) & ( n22158 )  ;
assign n23440 =  ( n92 ) & ( n22160 )  ;
assign n23441 =  ( n92 ) & ( n22162 )  ;
assign n23442 =  ( n92 ) & ( n22164 )  ;
assign n23443 =  ( n92 ) & ( n22166 )  ;
assign n23444 =  ( n92 ) & ( n22168 )  ;
assign n23445 =  ( n92 ) & ( n22170 )  ;
assign n23446 =  ( n93 ) & ( n22140 )  ;
assign n23447 =  ( n93 ) & ( n22142 )  ;
assign n23448 =  ( n93 ) & ( n22144 )  ;
assign n23449 =  ( n93 ) & ( n22146 )  ;
assign n23450 =  ( n93 ) & ( n22148 )  ;
assign n23451 =  ( n93 ) & ( n22150 )  ;
assign n23452 =  ( n93 ) & ( n22152 )  ;
assign n23453 =  ( n93 ) & ( n22154 )  ;
assign n23454 =  ( n93 ) & ( n22156 )  ;
assign n23455 =  ( n93 ) & ( n22158 )  ;
assign n23456 =  ( n93 ) & ( n22160 )  ;
assign n23457 =  ( n93 ) & ( n22162 )  ;
assign n23458 =  ( n93 ) & ( n22164 )  ;
assign n23459 =  ( n93 ) & ( n22166 )  ;
assign n23460 =  ( n93 ) & ( n22168 )  ;
assign n23461 =  ( n93 ) & ( n22170 )  ;
assign n23462 =  ( n94 ) & ( n22140 )  ;
assign n23463 =  ( n94 ) & ( n22142 )  ;
assign n23464 =  ( n94 ) & ( n22144 )  ;
assign n23465 =  ( n94 ) & ( n22146 )  ;
assign n23466 =  ( n94 ) & ( n22148 )  ;
assign n23467 =  ( n94 ) & ( n22150 )  ;
assign n23468 =  ( n94 ) & ( n22152 )  ;
assign n23469 =  ( n94 ) & ( n22154 )  ;
assign n23470 =  ( n94 ) & ( n22156 )  ;
assign n23471 =  ( n94 ) & ( n22158 )  ;
assign n23472 =  ( n94 ) & ( n22160 )  ;
assign n23473 =  ( n94 ) & ( n22162 )  ;
assign n23474 =  ( n94 ) & ( n22164 )  ;
assign n23475 =  ( n94 ) & ( n22166 )  ;
assign n23476 =  ( n94 ) & ( n22168 )  ;
assign n23477 =  ( n94 ) & ( n22170 )  ;
assign n23478 =  ( n95 ) & ( n22140 )  ;
assign n23479 =  ( n95 ) & ( n22142 )  ;
assign n23480 =  ( n95 ) & ( n22144 )  ;
assign n23481 =  ( n95 ) & ( n22146 )  ;
assign n23482 =  ( n95 ) & ( n22148 )  ;
assign n23483 =  ( n95 ) & ( n22150 )  ;
assign n23484 =  ( n95 ) & ( n22152 )  ;
assign n23485 =  ( n95 ) & ( n22154 )  ;
assign n23486 =  ( n95 ) & ( n22156 )  ;
assign n23487 =  ( n95 ) & ( n22158 )  ;
assign n23488 =  ( n95 ) & ( n22160 )  ;
assign n23489 =  ( n95 ) & ( n22162 )  ;
assign n23490 =  ( n95 ) & ( n22164 )  ;
assign n23491 =  ( n95 ) & ( n22166 )  ;
assign n23492 =  ( n95 ) & ( n22168 )  ;
assign n23493 =  ( n95 ) & ( n22170 )  ;
assign n23494 =  ( n96 ) & ( n22140 )  ;
assign n23495 =  ( n96 ) & ( n22142 )  ;
assign n23496 =  ( n96 ) & ( n22144 )  ;
assign n23497 =  ( n96 ) & ( n22146 )  ;
assign n23498 =  ( n96 ) & ( n22148 )  ;
assign n23499 =  ( n96 ) & ( n22150 )  ;
assign n23500 =  ( n96 ) & ( n22152 )  ;
assign n23501 =  ( n96 ) & ( n22154 )  ;
assign n23502 =  ( n96 ) & ( n22156 )  ;
assign n23503 =  ( n96 ) & ( n22158 )  ;
assign n23504 =  ( n96 ) & ( n22160 )  ;
assign n23505 =  ( n96 ) & ( n22162 )  ;
assign n23506 =  ( n96 ) & ( n22164 )  ;
assign n23507 =  ( n96 ) & ( n22166 )  ;
assign n23508 =  ( n96 ) & ( n22168 )  ;
assign n23509 =  ( n96 ) & ( n22170 )  ;
assign n23510 =  ( n97 ) & ( n22140 )  ;
assign n23511 =  ( n97 ) & ( n22142 )  ;
assign n23512 =  ( n97 ) & ( n22144 )  ;
assign n23513 =  ( n97 ) & ( n22146 )  ;
assign n23514 =  ( n97 ) & ( n22148 )  ;
assign n23515 =  ( n97 ) & ( n22150 )  ;
assign n23516 =  ( n97 ) & ( n22152 )  ;
assign n23517 =  ( n97 ) & ( n22154 )  ;
assign n23518 =  ( n97 ) & ( n22156 )  ;
assign n23519 =  ( n97 ) & ( n22158 )  ;
assign n23520 =  ( n97 ) & ( n22160 )  ;
assign n23521 =  ( n97 ) & ( n22162 )  ;
assign n23522 =  ( n97 ) & ( n22164 )  ;
assign n23523 =  ( n97 ) & ( n22166 )  ;
assign n23524 =  ( n97 ) & ( n22168 )  ;
assign n23525 =  ( n97 ) & ( n22170 )  ;
assign n23526 =  ( n98 ) & ( n22140 )  ;
assign n23527 =  ( n98 ) & ( n22142 )  ;
assign n23528 =  ( n98 ) & ( n22144 )  ;
assign n23529 =  ( n98 ) & ( n22146 )  ;
assign n23530 =  ( n98 ) & ( n22148 )  ;
assign n23531 =  ( n98 ) & ( n22150 )  ;
assign n23532 =  ( n98 ) & ( n22152 )  ;
assign n23533 =  ( n98 ) & ( n22154 )  ;
assign n23534 =  ( n98 ) & ( n22156 )  ;
assign n23535 =  ( n98 ) & ( n22158 )  ;
assign n23536 =  ( n98 ) & ( n22160 )  ;
assign n23537 =  ( n98 ) & ( n22162 )  ;
assign n23538 =  ( n98 ) & ( n22164 )  ;
assign n23539 =  ( n98 ) & ( n22166 )  ;
assign n23540 =  ( n98 ) & ( n22168 )  ;
assign n23541 =  ( n98 ) & ( n22170 )  ;
assign n23542 =  ( n99 ) & ( n22140 )  ;
assign n23543 =  ( n99 ) & ( n22142 )  ;
assign n23544 =  ( n99 ) & ( n22144 )  ;
assign n23545 =  ( n99 ) & ( n22146 )  ;
assign n23546 =  ( n99 ) & ( n22148 )  ;
assign n23547 =  ( n99 ) & ( n22150 )  ;
assign n23548 =  ( n99 ) & ( n22152 )  ;
assign n23549 =  ( n99 ) & ( n22154 )  ;
assign n23550 =  ( n99 ) & ( n22156 )  ;
assign n23551 =  ( n99 ) & ( n22158 )  ;
assign n23552 =  ( n99 ) & ( n22160 )  ;
assign n23553 =  ( n99 ) & ( n22162 )  ;
assign n23554 =  ( n99 ) & ( n22164 )  ;
assign n23555 =  ( n99 ) & ( n22166 )  ;
assign n23556 =  ( n99 ) & ( n22168 )  ;
assign n23557 =  ( n99 ) & ( n22170 )  ;
assign n23558 =  ( n100 ) & ( n22140 )  ;
assign n23559 =  ( n100 ) & ( n22142 )  ;
assign n23560 =  ( n100 ) & ( n22144 )  ;
assign n23561 =  ( n100 ) & ( n22146 )  ;
assign n23562 =  ( n100 ) & ( n22148 )  ;
assign n23563 =  ( n100 ) & ( n22150 )  ;
assign n23564 =  ( n100 ) & ( n22152 )  ;
assign n23565 =  ( n100 ) & ( n22154 )  ;
assign n23566 =  ( n100 ) & ( n22156 )  ;
assign n23567 =  ( n100 ) & ( n22158 )  ;
assign n23568 =  ( n100 ) & ( n22160 )  ;
assign n23569 =  ( n100 ) & ( n22162 )  ;
assign n23570 =  ( n100 ) & ( n22164 )  ;
assign n23571 =  ( n100 ) & ( n22166 )  ;
assign n23572 =  ( n100 ) & ( n22168 )  ;
assign n23573 =  ( n100 ) & ( n22170 )  ;
assign n23574 =  ( n101 ) & ( n22140 )  ;
assign n23575 =  ( n101 ) & ( n22142 )  ;
assign n23576 =  ( n101 ) & ( n22144 )  ;
assign n23577 =  ( n101 ) & ( n22146 )  ;
assign n23578 =  ( n101 ) & ( n22148 )  ;
assign n23579 =  ( n101 ) & ( n22150 )  ;
assign n23580 =  ( n101 ) & ( n22152 )  ;
assign n23581 =  ( n101 ) & ( n22154 )  ;
assign n23582 =  ( n101 ) & ( n22156 )  ;
assign n23583 =  ( n101 ) & ( n22158 )  ;
assign n23584 =  ( n101 ) & ( n22160 )  ;
assign n23585 =  ( n101 ) & ( n22162 )  ;
assign n23586 =  ( n101 ) & ( n22164 )  ;
assign n23587 =  ( n101 ) & ( n22166 )  ;
assign n23588 =  ( n101 ) & ( n22168 )  ;
assign n23589 =  ( n101 ) & ( n22170 )  ;
assign n23590 =  ( n102 ) & ( n22140 )  ;
assign n23591 =  ( n102 ) & ( n22142 )  ;
assign n23592 =  ( n102 ) & ( n22144 )  ;
assign n23593 =  ( n102 ) & ( n22146 )  ;
assign n23594 =  ( n102 ) & ( n22148 )  ;
assign n23595 =  ( n102 ) & ( n22150 )  ;
assign n23596 =  ( n102 ) & ( n22152 )  ;
assign n23597 =  ( n102 ) & ( n22154 )  ;
assign n23598 =  ( n102 ) & ( n22156 )  ;
assign n23599 =  ( n102 ) & ( n22158 )  ;
assign n23600 =  ( n102 ) & ( n22160 )  ;
assign n23601 =  ( n102 ) & ( n22162 )  ;
assign n23602 =  ( n102 ) & ( n22164 )  ;
assign n23603 =  ( n102 ) & ( n22166 )  ;
assign n23604 =  ( n102 ) & ( n22168 )  ;
assign n23605 =  ( n102 ) & ( n22170 )  ;
assign n23606 =  ( n103 ) & ( n22140 )  ;
assign n23607 =  ( n103 ) & ( n22142 )  ;
assign n23608 =  ( n103 ) & ( n22144 )  ;
assign n23609 =  ( n103 ) & ( n22146 )  ;
assign n23610 =  ( n103 ) & ( n22148 )  ;
assign n23611 =  ( n103 ) & ( n22150 )  ;
assign n23612 =  ( n103 ) & ( n22152 )  ;
assign n23613 =  ( n103 ) & ( n22154 )  ;
assign n23614 =  ( n103 ) & ( n22156 )  ;
assign n23615 =  ( n103 ) & ( n22158 )  ;
assign n23616 =  ( n103 ) & ( n22160 )  ;
assign n23617 =  ( n103 ) & ( n22162 )  ;
assign n23618 =  ( n103 ) & ( n22164 )  ;
assign n23619 =  ( n103 ) & ( n22166 )  ;
assign n23620 =  ( n103 ) & ( n22168 )  ;
assign n23621 =  ( n103 ) & ( n22170 )  ;
assign n23622 =  ( n104 ) & ( n22140 )  ;
assign n23623 =  ( n104 ) & ( n22142 )  ;
assign n23624 =  ( n104 ) & ( n22144 )  ;
assign n23625 =  ( n104 ) & ( n22146 )  ;
assign n23626 =  ( n104 ) & ( n22148 )  ;
assign n23627 =  ( n104 ) & ( n22150 )  ;
assign n23628 =  ( n104 ) & ( n22152 )  ;
assign n23629 =  ( n104 ) & ( n22154 )  ;
assign n23630 =  ( n104 ) & ( n22156 )  ;
assign n23631 =  ( n104 ) & ( n22158 )  ;
assign n23632 =  ( n104 ) & ( n22160 )  ;
assign n23633 =  ( n104 ) & ( n22162 )  ;
assign n23634 =  ( n104 ) & ( n22164 )  ;
assign n23635 =  ( n104 ) & ( n22166 )  ;
assign n23636 =  ( n104 ) & ( n22168 )  ;
assign n23637 =  ( n104 ) & ( n22170 )  ;
assign n23638 =  ( n105 ) & ( n22140 )  ;
assign n23639 =  ( n105 ) & ( n22142 )  ;
assign n23640 =  ( n105 ) & ( n22144 )  ;
assign n23641 =  ( n105 ) & ( n22146 )  ;
assign n23642 =  ( n105 ) & ( n22148 )  ;
assign n23643 =  ( n105 ) & ( n22150 )  ;
assign n23644 =  ( n105 ) & ( n22152 )  ;
assign n23645 =  ( n105 ) & ( n22154 )  ;
assign n23646 =  ( n105 ) & ( n22156 )  ;
assign n23647 =  ( n105 ) & ( n22158 )  ;
assign n23648 =  ( n105 ) & ( n22160 )  ;
assign n23649 =  ( n105 ) & ( n22162 )  ;
assign n23650 =  ( n105 ) & ( n22164 )  ;
assign n23651 =  ( n105 ) & ( n22166 )  ;
assign n23652 =  ( n105 ) & ( n22168 )  ;
assign n23653 =  ( n105 ) & ( n22170 )  ;
assign n23654 =  ( n106 ) & ( n22140 )  ;
assign n23655 =  ( n106 ) & ( n22142 )  ;
assign n23656 =  ( n106 ) & ( n22144 )  ;
assign n23657 =  ( n106 ) & ( n22146 )  ;
assign n23658 =  ( n106 ) & ( n22148 )  ;
assign n23659 =  ( n106 ) & ( n22150 )  ;
assign n23660 =  ( n106 ) & ( n22152 )  ;
assign n23661 =  ( n106 ) & ( n22154 )  ;
assign n23662 =  ( n106 ) & ( n22156 )  ;
assign n23663 =  ( n106 ) & ( n22158 )  ;
assign n23664 =  ( n106 ) & ( n22160 )  ;
assign n23665 =  ( n106 ) & ( n22162 )  ;
assign n23666 =  ( n106 ) & ( n22164 )  ;
assign n23667 =  ( n106 ) & ( n22166 )  ;
assign n23668 =  ( n106 ) & ( n22168 )  ;
assign n23669 =  ( n106 ) & ( n22170 )  ;
assign n23670 =  ( n107 ) & ( n22140 )  ;
assign n23671 =  ( n107 ) & ( n22142 )  ;
assign n23672 =  ( n107 ) & ( n22144 )  ;
assign n23673 =  ( n107 ) & ( n22146 )  ;
assign n23674 =  ( n107 ) & ( n22148 )  ;
assign n23675 =  ( n107 ) & ( n22150 )  ;
assign n23676 =  ( n107 ) & ( n22152 )  ;
assign n23677 =  ( n107 ) & ( n22154 )  ;
assign n23678 =  ( n107 ) & ( n22156 )  ;
assign n23679 =  ( n107 ) & ( n22158 )  ;
assign n23680 =  ( n107 ) & ( n22160 )  ;
assign n23681 =  ( n107 ) & ( n22162 )  ;
assign n23682 =  ( n107 ) & ( n22164 )  ;
assign n23683 =  ( n107 ) & ( n22166 )  ;
assign n23684 =  ( n107 ) & ( n22168 )  ;
assign n23685 =  ( n107 ) & ( n22170 )  ;
assign n23686 =  ( n108 ) & ( n22140 )  ;
assign n23687 =  ( n108 ) & ( n22142 )  ;
assign n23688 =  ( n108 ) & ( n22144 )  ;
assign n23689 =  ( n108 ) & ( n22146 )  ;
assign n23690 =  ( n108 ) & ( n22148 )  ;
assign n23691 =  ( n108 ) & ( n22150 )  ;
assign n23692 =  ( n108 ) & ( n22152 )  ;
assign n23693 =  ( n108 ) & ( n22154 )  ;
assign n23694 =  ( n108 ) & ( n22156 )  ;
assign n23695 =  ( n108 ) & ( n22158 )  ;
assign n23696 =  ( n108 ) & ( n22160 )  ;
assign n23697 =  ( n108 ) & ( n22162 )  ;
assign n23698 =  ( n108 ) & ( n22164 )  ;
assign n23699 =  ( n108 ) & ( n22166 )  ;
assign n23700 =  ( n108 ) & ( n22168 )  ;
assign n23701 =  ( n108 ) & ( n22170 )  ;
assign n23702 =  ( n23701 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n23703 =  ( n23700 ) ? ( VREG_0_1 ) : ( n23702 ) ;
assign n23704 =  ( n23699 ) ? ( VREG_0_2 ) : ( n23703 ) ;
assign n23705 =  ( n23698 ) ? ( VREG_0_3 ) : ( n23704 ) ;
assign n23706 =  ( n23697 ) ? ( VREG_0_4 ) : ( n23705 ) ;
assign n23707 =  ( n23696 ) ? ( VREG_0_5 ) : ( n23706 ) ;
assign n23708 =  ( n23695 ) ? ( VREG_0_6 ) : ( n23707 ) ;
assign n23709 =  ( n23694 ) ? ( VREG_0_7 ) : ( n23708 ) ;
assign n23710 =  ( n23693 ) ? ( VREG_0_8 ) : ( n23709 ) ;
assign n23711 =  ( n23692 ) ? ( VREG_0_9 ) : ( n23710 ) ;
assign n23712 =  ( n23691 ) ? ( VREG_0_10 ) : ( n23711 ) ;
assign n23713 =  ( n23690 ) ? ( VREG_0_11 ) : ( n23712 ) ;
assign n23714 =  ( n23689 ) ? ( VREG_0_12 ) : ( n23713 ) ;
assign n23715 =  ( n23688 ) ? ( VREG_0_13 ) : ( n23714 ) ;
assign n23716 =  ( n23687 ) ? ( VREG_0_14 ) : ( n23715 ) ;
assign n23717 =  ( n23686 ) ? ( VREG_0_15 ) : ( n23716 ) ;
assign n23718 =  ( n23685 ) ? ( VREG_1_0 ) : ( n23717 ) ;
assign n23719 =  ( n23684 ) ? ( VREG_1_1 ) : ( n23718 ) ;
assign n23720 =  ( n23683 ) ? ( VREG_1_2 ) : ( n23719 ) ;
assign n23721 =  ( n23682 ) ? ( VREG_1_3 ) : ( n23720 ) ;
assign n23722 =  ( n23681 ) ? ( VREG_1_4 ) : ( n23721 ) ;
assign n23723 =  ( n23680 ) ? ( VREG_1_5 ) : ( n23722 ) ;
assign n23724 =  ( n23679 ) ? ( VREG_1_6 ) : ( n23723 ) ;
assign n23725 =  ( n23678 ) ? ( VREG_1_7 ) : ( n23724 ) ;
assign n23726 =  ( n23677 ) ? ( VREG_1_8 ) : ( n23725 ) ;
assign n23727 =  ( n23676 ) ? ( VREG_1_9 ) : ( n23726 ) ;
assign n23728 =  ( n23675 ) ? ( VREG_1_10 ) : ( n23727 ) ;
assign n23729 =  ( n23674 ) ? ( VREG_1_11 ) : ( n23728 ) ;
assign n23730 =  ( n23673 ) ? ( VREG_1_12 ) : ( n23729 ) ;
assign n23731 =  ( n23672 ) ? ( VREG_1_13 ) : ( n23730 ) ;
assign n23732 =  ( n23671 ) ? ( VREG_1_14 ) : ( n23731 ) ;
assign n23733 =  ( n23670 ) ? ( VREG_1_15 ) : ( n23732 ) ;
assign n23734 =  ( n23669 ) ? ( VREG_2_0 ) : ( n23733 ) ;
assign n23735 =  ( n23668 ) ? ( VREG_2_1 ) : ( n23734 ) ;
assign n23736 =  ( n23667 ) ? ( VREG_2_2 ) : ( n23735 ) ;
assign n23737 =  ( n23666 ) ? ( VREG_2_3 ) : ( n23736 ) ;
assign n23738 =  ( n23665 ) ? ( VREG_2_4 ) : ( n23737 ) ;
assign n23739 =  ( n23664 ) ? ( VREG_2_5 ) : ( n23738 ) ;
assign n23740 =  ( n23663 ) ? ( VREG_2_6 ) : ( n23739 ) ;
assign n23741 =  ( n23662 ) ? ( VREG_2_7 ) : ( n23740 ) ;
assign n23742 =  ( n23661 ) ? ( VREG_2_8 ) : ( n23741 ) ;
assign n23743 =  ( n23660 ) ? ( VREG_2_9 ) : ( n23742 ) ;
assign n23744 =  ( n23659 ) ? ( VREG_2_10 ) : ( n23743 ) ;
assign n23745 =  ( n23658 ) ? ( VREG_2_11 ) : ( n23744 ) ;
assign n23746 =  ( n23657 ) ? ( VREG_2_12 ) : ( n23745 ) ;
assign n23747 =  ( n23656 ) ? ( VREG_2_13 ) : ( n23746 ) ;
assign n23748 =  ( n23655 ) ? ( VREG_2_14 ) : ( n23747 ) ;
assign n23749 =  ( n23654 ) ? ( VREG_2_15 ) : ( n23748 ) ;
assign n23750 =  ( n23653 ) ? ( VREG_3_0 ) : ( n23749 ) ;
assign n23751 =  ( n23652 ) ? ( VREG_3_1 ) : ( n23750 ) ;
assign n23752 =  ( n23651 ) ? ( VREG_3_2 ) : ( n23751 ) ;
assign n23753 =  ( n23650 ) ? ( VREG_3_3 ) : ( n23752 ) ;
assign n23754 =  ( n23649 ) ? ( VREG_3_4 ) : ( n23753 ) ;
assign n23755 =  ( n23648 ) ? ( VREG_3_5 ) : ( n23754 ) ;
assign n23756 =  ( n23647 ) ? ( VREG_3_6 ) : ( n23755 ) ;
assign n23757 =  ( n23646 ) ? ( VREG_3_7 ) : ( n23756 ) ;
assign n23758 =  ( n23645 ) ? ( VREG_3_8 ) : ( n23757 ) ;
assign n23759 =  ( n23644 ) ? ( VREG_3_9 ) : ( n23758 ) ;
assign n23760 =  ( n23643 ) ? ( VREG_3_10 ) : ( n23759 ) ;
assign n23761 =  ( n23642 ) ? ( VREG_3_11 ) : ( n23760 ) ;
assign n23762 =  ( n23641 ) ? ( VREG_3_12 ) : ( n23761 ) ;
assign n23763 =  ( n23640 ) ? ( VREG_3_13 ) : ( n23762 ) ;
assign n23764 =  ( n23639 ) ? ( VREG_3_14 ) : ( n23763 ) ;
assign n23765 =  ( n23638 ) ? ( VREG_3_15 ) : ( n23764 ) ;
assign n23766 =  ( n23637 ) ? ( VREG_4_0 ) : ( n23765 ) ;
assign n23767 =  ( n23636 ) ? ( VREG_4_1 ) : ( n23766 ) ;
assign n23768 =  ( n23635 ) ? ( VREG_4_2 ) : ( n23767 ) ;
assign n23769 =  ( n23634 ) ? ( VREG_4_3 ) : ( n23768 ) ;
assign n23770 =  ( n23633 ) ? ( VREG_4_4 ) : ( n23769 ) ;
assign n23771 =  ( n23632 ) ? ( VREG_4_5 ) : ( n23770 ) ;
assign n23772 =  ( n23631 ) ? ( VREG_4_6 ) : ( n23771 ) ;
assign n23773 =  ( n23630 ) ? ( VREG_4_7 ) : ( n23772 ) ;
assign n23774 =  ( n23629 ) ? ( VREG_4_8 ) : ( n23773 ) ;
assign n23775 =  ( n23628 ) ? ( VREG_4_9 ) : ( n23774 ) ;
assign n23776 =  ( n23627 ) ? ( VREG_4_10 ) : ( n23775 ) ;
assign n23777 =  ( n23626 ) ? ( VREG_4_11 ) : ( n23776 ) ;
assign n23778 =  ( n23625 ) ? ( VREG_4_12 ) : ( n23777 ) ;
assign n23779 =  ( n23624 ) ? ( VREG_4_13 ) : ( n23778 ) ;
assign n23780 =  ( n23623 ) ? ( VREG_4_14 ) : ( n23779 ) ;
assign n23781 =  ( n23622 ) ? ( VREG_4_15 ) : ( n23780 ) ;
assign n23782 =  ( n23621 ) ? ( VREG_5_0 ) : ( n23781 ) ;
assign n23783 =  ( n23620 ) ? ( VREG_5_1 ) : ( n23782 ) ;
assign n23784 =  ( n23619 ) ? ( VREG_5_2 ) : ( n23783 ) ;
assign n23785 =  ( n23618 ) ? ( VREG_5_3 ) : ( n23784 ) ;
assign n23786 =  ( n23617 ) ? ( VREG_5_4 ) : ( n23785 ) ;
assign n23787 =  ( n23616 ) ? ( VREG_5_5 ) : ( n23786 ) ;
assign n23788 =  ( n23615 ) ? ( VREG_5_6 ) : ( n23787 ) ;
assign n23789 =  ( n23614 ) ? ( VREG_5_7 ) : ( n23788 ) ;
assign n23790 =  ( n23613 ) ? ( VREG_5_8 ) : ( n23789 ) ;
assign n23791 =  ( n23612 ) ? ( VREG_5_9 ) : ( n23790 ) ;
assign n23792 =  ( n23611 ) ? ( VREG_5_10 ) : ( n23791 ) ;
assign n23793 =  ( n23610 ) ? ( VREG_5_11 ) : ( n23792 ) ;
assign n23794 =  ( n23609 ) ? ( VREG_5_12 ) : ( n23793 ) ;
assign n23795 =  ( n23608 ) ? ( VREG_5_13 ) : ( n23794 ) ;
assign n23796 =  ( n23607 ) ? ( VREG_5_14 ) : ( n23795 ) ;
assign n23797 =  ( n23606 ) ? ( VREG_5_15 ) : ( n23796 ) ;
assign n23798 =  ( n23605 ) ? ( VREG_6_0 ) : ( n23797 ) ;
assign n23799 =  ( n23604 ) ? ( VREG_6_1 ) : ( n23798 ) ;
assign n23800 =  ( n23603 ) ? ( VREG_6_2 ) : ( n23799 ) ;
assign n23801 =  ( n23602 ) ? ( VREG_6_3 ) : ( n23800 ) ;
assign n23802 =  ( n23601 ) ? ( VREG_6_4 ) : ( n23801 ) ;
assign n23803 =  ( n23600 ) ? ( VREG_6_5 ) : ( n23802 ) ;
assign n23804 =  ( n23599 ) ? ( VREG_6_6 ) : ( n23803 ) ;
assign n23805 =  ( n23598 ) ? ( VREG_6_7 ) : ( n23804 ) ;
assign n23806 =  ( n23597 ) ? ( VREG_6_8 ) : ( n23805 ) ;
assign n23807 =  ( n23596 ) ? ( VREG_6_9 ) : ( n23806 ) ;
assign n23808 =  ( n23595 ) ? ( VREG_6_10 ) : ( n23807 ) ;
assign n23809 =  ( n23594 ) ? ( VREG_6_11 ) : ( n23808 ) ;
assign n23810 =  ( n23593 ) ? ( VREG_6_12 ) : ( n23809 ) ;
assign n23811 =  ( n23592 ) ? ( VREG_6_13 ) : ( n23810 ) ;
assign n23812 =  ( n23591 ) ? ( VREG_6_14 ) : ( n23811 ) ;
assign n23813 =  ( n23590 ) ? ( VREG_6_15 ) : ( n23812 ) ;
assign n23814 =  ( n23589 ) ? ( VREG_7_0 ) : ( n23813 ) ;
assign n23815 =  ( n23588 ) ? ( VREG_7_1 ) : ( n23814 ) ;
assign n23816 =  ( n23587 ) ? ( VREG_7_2 ) : ( n23815 ) ;
assign n23817 =  ( n23586 ) ? ( VREG_7_3 ) : ( n23816 ) ;
assign n23818 =  ( n23585 ) ? ( VREG_7_4 ) : ( n23817 ) ;
assign n23819 =  ( n23584 ) ? ( VREG_7_5 ) : ( n23818 ) ;
assign n23820 =  ( n23583 ) ? ( VREG_7_6 ) : ( n23819 ) ;
assign n23821 =  ( n23582 ) ? ( VREG_7_7 ) : ( n23820 ) ;
assign n23822 =  ( n23581 ) ? ( VREG_7_8 ) : ( n23821 ) ;
assign n23823 =  ( n23580 ) ? ( VREG_7_9 ) : ( n23822 ) ;
assign n23824 =  ( n23579 ) ? ( VREG_7_10 ) : ( n23823 ) ;
assign n23825 =  ( n23578 ) ? ( VREG_7_11 ) : ( n23824 ) ;
assign n23826 =  ( n23577 ) ? ( VREG_7_12 ) : ( n23825 ) ;
assign n23827 =  ( n23576 ) ? ( VREG_7_13 ) : ( n23826 ) ;
assign n23828 =  ( n23575 ) ? ( VREG_7_14 ) : ( n23827 ) ;
assign n23829 =  ( n23574 ) ? ( VREG_7_15 ) : ( n23828 ) ;
assign n23830 =  ( n23573 ) ? ( VREG_8_0 ) : ( n23829 ) ;
assign n23831 =  ( n23572 ) ? ( VREG_8_1 ) : ( n23830 ) ;
assign n23832 =  ( n23571 ) ? ( VREG_8_2 ) : ( n23831 ) ;
assign n23833 =  ( n23570 ) ? ( VREG_8_3 ) : ( n23832 ) ;
assign n23834 =  ( n23569 ) ? ( VREG_8_4 ) : ( n23833 ) ;
assign n23835 =  ( n23568 ) ? ( VREG_8_5 ) : ( n23834 ) ;
assign n23836 =  ( n23567 ) ? ( VREG_8_6 ) : ( n23835 ) ;
assign n23837 =  ( n23566 ) ? ( VREG_8_7 ) : ( n23836 ) ;
assign n23838 =  ( n23565 ) ? ( VREG_8_8 ) : ( n23837 ) ;
assign n23839 =  ( n23564 ) ? ( VREG_8_9 ) : ( n23838 ) ;
assign n23840 =  ( n23563 ) ? ( VREG_8_10 ) : ( n23839 ) ;
assign n23841 =  ( n23562 ) ? ( VREG_8_11 ) : ( n23840 ) ;
assign n23842 =  ( n23561 ) ? ( VREG_8_12 ) : ( n23841 ) ;
assign n23843 =  ( n23560 ) ? ( VREG_8_13 ) : ( n23842 ) ;
assign n23844 =  ( n23559 ) ? ( VREG_8_14 ) : ( n23843 ) ;
assign n23845 =  ( n23558 ) ? ( VREG_8_15 ) : ( n23844 ) ;
assign n23846 =  ( n23557 ) ? ( VREG_9_0 ) : ( n23845 ) ;
assign n23847 =  ( n23556 ) ? ( VREG_9_1 ) : ( n23846 ) ;
assign n23848 =  ( n23555 ) ? ( VREG_9_2 ) : ( n23847 ) ;
assign n23849 =  ( n23554 ) ? ( VREG_9_3 ) : ( n23848 ) ;
assign n23850 =  ( n23553 ) ? ( VREG_9_4 ) : ( n23849 ) ;
assign n23851 =  ( n23552 ) ? ( VREG_9_5 ) : ( n23850 ) ;
assign n23852 =  ( n23551 ) ? ( VREG_9_6 ) : ( n23851 ) ;
assign n23853 =  ( n23550 ) ? ( VREG_9_7 ) : ( n23852 ) ;
assign n23854 =  ( n23549 ) ? ( VREG_9_8 ) : ( n23853 ) ;
assign n23855 =  ( n23548 ) ? ( VREG_9_9 ) : ( n23854 ) ;
assign n23856 =  ( n23547 ) ? ( VREG_9_10 ) : ( n23855 ) ;
assign n23857 =  ( n23546 ) ? ( VREG_9_11 ) : ( n23856 ) ;
assign n23858 =  ( n23545 ) ? ( VREG_9_12 ) : ( n23857 ) ;
assign n23859 =  ( n23544 ) ? ( VREG_9_13 ) : ( n23858 ) ;
assign n23860 =  ( n23543 ) ? ( VREG_9_14 ) : ( n23859 ) ;
assign n23861 =  ( n23542 ) ? ( VREG_9_15 ) : ( n23860 ) ;
assign n23862 =  ( n23541 ) ? ( VREG_10_0 ) : ( n23861 ) ;
assign n23863 =  ( n23540 ) ? ( VREG_10_1 ) : ( n23862 ) ;
assign n23864 =  ( n23539 ) ? ( VREG_10_2 ) : ( n23863 ) ;
assign n23865 =  ( n23538 ) ? ( VREG_10_3 ) : ( n23864 ) ;
assign n23866 =  ( n23537 ) ? ( VREG_10_4 ) : ( n23865 ) ;
assign n23867 =  ( n23536 ) ? ( VREG_10_5 ) : ( n23866 ) ;
assign n23868 =  ( n23535 ) ? ( VREG_10_6 ) : ( n23867 ) ;
assign n23869 =  ( n23534 ) ? ( VREG_10_7 ) : ( n23868 ) ;
assign n23870 =  ( n23533 ) ? ( VREG_10_8 ) : ( n23869 ) ;
assign n23871 =  ( n23532 ) ? ( VREG_10_9 ) : ( n23870 ) ;
assign n23872 =  ( n23531 ) ? ( VREG_10_10 ) : ( n23871 ) ;
assign n23873 =  ( n23530 ) ? ( VREG_10_11 ) : ( n23872 ) ;
assign n23874 =  ( n23529 ) ? ( VREG_10_12 ) : ( n23873 ) ;
assign n23875 =  ( n23528 ) ? ( VREG_10_13 ) : ( n23874 ) ;
assign n23876 =  ( n23527 ) ? ( VREG_10_14 ) : ( n23875 ) ;
assign n23877 =  ( n23526 ) ? ( VREG_10_15 ) : ( n23876 ) ;
assign n23878 =  ( n23525 ) ? ( VREG_11_0 ) : ( n23877 ) ;
assign n23879 =  ( n23524 ) ? ( VREG_11_1 ) : ( n23878 ) ;
assign n23880 =  ( n23523 ) ? ( VREG_11_2 ) : ( n23879 ) ;
assign n23881 =  ( n23522 ) ? ( VREG_11_3 ) : ( n23880 ) ;
assign n23882 =  ( n23521 ) ? ( VREG_11_4 ) : ( n23881 ) ;
assign n23883 =  ( n23520 ) ? ( VREG_11_5 ) : ( n23882 ) ;
assign n23884 =  ( n23519 ) ? ( VREG_11_6 ) : ( n23883 ) ;
assign n23885 =  ( n23518 ) ? ( VREG_11_7 ) : ( n23884 ) ;
assign n23886 =  ( n23517 ) ? ( VREG_11_8 ) : ( n23885 ) ;
assign n23887 =  ( n23516 ) ? ( VREG_11_9 ) : ( n23886 ) ;
assign n23888 =  ( n23515 ) ? ( VREG_11_10 ) : ( n23887 ) ;
assign n23889 =  ( n23514 ) ? ( VREG_11_11 ) : ( n23888 ) ;
assign n23890 =  ( n23513 ) ? ( VREG_11_12 ) : ( n23889 ) ;
assign n23891 =  ( n23512 ) ? ( VREG_11_13 ) : ( n23890 ) ;
assign n23892 =  ( n23511 ) ? ( VREG_11_14 ) : ( n23891 ) ;
assign n23893 =  ( n23510 ) ? ( VREG_11_15 ) : ( n23892 ) ;
assign n23894 =  ( n23509 ) ? ( VREG_12_0 ) : ( n23893 ) ;
assign n23895 =  ( n23508 ) ? ( VREG_12_1 ) : ( n23894 ) ;
assign n23896 =  ( n23507 ) ? ( VREG_12_2 ) : ( n23895 ) ;
assign n23897 =  ( n23506 ) ? ( VREG_12_3 ) : ( n23896 ) ;
assign n23898 =  ( n23505 ) ? ( VREG_12_4 ) : ( n23897 ) ;
assign n23899 =  ( n23504 ) ? ( VREG_12_5 ) : ( n23898 ) ;
assign n23900 =  ( n23503 ) ? ( VREG_12_6 ) : ( n23899 ) ;
assign n23901 =  ( n23502 ) ? ( VREG_12_7 ) : ( n23900 ) ;
assign n23902 =  ( n23501 ) ? ( VREG_12_8 ) : ( n23901 ) ;
assign n23903 =  ( n23500 ) ? ( VREG_12_9 ) : ( n23902 ) ;
assign n23904 =  ( n23499 ) ? ( VREG_12_10 ) : ( n23903 ) ;
assign n23905 =  ( n23498 ) ? ( VREG_12_11 ) : ( n23904 ) ;
assign n23906 =  ( n23497 ) ? ( VREG_12_12 ) : ( n23905 ) ;
assign n23907 =  ( n23496 ) ? ( VREG_12_13 ) : ( n23906 ) ;
assign n23908 =  ( n23495 ) ? ( VREG_12_14 ) : ( n23907 ) ;
assign n23909 =  ( n23494 ) ? ( VREG_12_15 ) : ( n23908 ) ;
assign n23910 =  ( n23493 ) ? ( VREG_13_0 ) : ( n23909 ) ;
assign n23911 =  ( n23492 ) ? ( VREG_13_1 ) : ( n23910 ) ;
assign n23912 =  ( n23491 ) ? ( VREG_13_2 ) : ( n23911 ) ;
assign n23913 =  ( n23490 ) ? ( VREG_13_3 ) : ( n23912 ) ;
assign n23914 =  ( n23489 ) ? ( VREG_13_4 ) : ( n23913 ) ;
assign n23915 =  ( n23488 ) ? ( VREG_13_5 ) : ( n23914 ) ;
assign n23916 =  ( n23487 ) ? ( VREG_13_6 ) : ( n23915 ) ;
assign n23917 =  ( n23486 ) ? ( VREG_13_7 ) : ( n23916 ) ;
assign n23918 =  ( n23485 ) ? ( VREG_13_8 ) : ( n23917 ) ;
assign n23919 =  ( n23484 ) ? ( VREG_13_9 ) : ( n23918 ) ;
assign n23920 =  ( n23483 ) ? ( VREG_13_10 ) : ( n23919 ) ;
assign n23921 =  ( n23482 ) ? ( VREG_13_11 ) : ( n23920 ) ;
assign n23922 =  ( n23481 ) ? ( VREG_13_12 ) : ( n23921 ) ;
assign n23923 =  ( n23480 ) ? ( VREG_13_13 ) : ( n23922 ) ;
assign n23924 =  ( n23479 ) ? ( VREG_13_14 ) : ( n23923 ) ;
assign n23925 =  ( n23478 ) ? ( VREG_13_15 ) : ( n23924 ) ;
assign n23926 =  ( n23477 ) ? ( VREG_14_0 ) : ( n23925 ) ;
assign n23927 =  ( n23476 ) ? ( VREG_14_1 ) : ( n23926 ) ;
assign n23928 =  ( n23475 ) ? ( VREG_14_2 ) : ( n23927 ) ;
assign n23929 =  ( n23474 ) ? ( VREG_14_3 ) : ( n23928 ) ;
assign n23930 =  ( n23473 ) ? ( VREG_14_4 ) : ( n23929 ) ;
assign n23931 =  ( n23472 ) ? ( VREG_14_5 ) : ( n23930 ) ;
assign n23932 =  ( n23471 ) ? ( VREG_14_6 ) : ( n23931 ) ;
assign n23933 =  ( n23470 ) ? ( VREG_14_7 ) : ( n23932 ) ;
assign n23934 =  ( n23469 ) ? ( VREG_14_8 ) : ( n23933 ) ;
assign n23935 =  ( n23468 ) ? ( VREG_14_9 ) : ( n23934 ) ;
assign n23936 =  ( n23467 ) ? ( VREG_14_10 ) : ( n23935 ) ;
assign n23937 =  ( n23466 ) ? ( VREG_14_11 ) : ( n23936 ) ;
assign n23938 =  ( n23465 ) ? ( VREG_14_12 ) : ( n23937 ) ;
assign n23939 =  ( n23464 ) ? ( VREG_14_13 ) : ( n23938 ) ;
assign n23940 =  ( n23463 ) ? ( VREG_14_14 ) : ( n23939 ) ;
assign n23941 =  ( n23462 ) ? ( VREG_14_15 ) : ( n23940 ) ;
assign n23942 =  ( n23461 ) ? ( VREG_15_0 ) : ( n23941 ) ;
assign n23943 =  ( n23460 ) ? ( VREG_15_1 ) : ( n23942 ) ;
assign n23944 =  ( n23459 ) ? ( VREG_15_2 ) : ( n23943 ) ;
assign n23945 =  ( n23458 ) ? ( VREG_15_3 ) : ( n23944 ) ;
assign n23946 =  ( n23457 ) ? ( VREG_15_4 ) : ( n23945 ) ;
assign n23947 =  ( n23456 ) ? ( VREG_15_5 ) : ( n23946 ) ;
assign n23948 =  ( n23455 ) ? ( VREG_15_6 ) : ( n23947 ) ;
assign n23949 =  ( n23454 ) ? ( VREG_15_7 ) : ( n23948 ) ;
assign n23950 =  ( n23453 ) ? ( VREG_15_8 ) : ( n23949 ) ;
assign n23951 =  ( n23452 ) ? ( VREG_15_9 ) : ( n23950 ) ;
assign n23952 =  ( n23451 ) ? ( VREG_15_10 ) : ( n23951 ) ;
assign n23953 =  ( n23450 ) ? ( VREG_15_11 ) : ( n23952 ) ;
assign n23954 =  ( n23449 ) ? ( VREG_15_12 ) : ( n23953 ) ;
assign n23955 =  ( n23448 ) ? ( VREG_15_13 ) : ( n23954 ) ;
assign n23956 =  ( n23447 ) ? ( VREG_15_14 ) : ( n23955 ) ;
assign n23957 =  ( n23446 ) ? ( VREG_15_15 ) : ( n23956 ) ;
assign n23958 =  ( n23445 ) ? ( VREG_16_0 ) : ( n23957 ) ;
assign n23959 =  ( n23444 ) ? ( VREG_16_1 ) : ( n23958 ) ;
assign n23960 =  ( n23443 ) ? ( VREG_16_2 ) : ( n23959 ) ;
assign n23961 =  ( n23442 ) ? ( VREG_16_3 ) : ( n23960 ) ;
assign n23962 =  ( n23441 ) ? ( VREG_16_4 ) : ( n23961 ) ;
assign n23963 =  ( n23440 ) ? ( VREG_16_5 ) : ( n23962 ) ;
assign n23964 =  ( n23439 ) ? ( VREG_16_6 ) : ( n23963 ) ;
assign n23965 =  ( n23438 ) ? ( VREG_16_7 ) : ( n23964 ) ;
assign n23966 =  ( n23437 ) ? ( VREG_16_8 ) : ( n23965 ) ;
assign n23967 =  ( n23436 ) ? ( VREG_16_9 ) : ( n23966 ) ;
assign n23968 =  ( n23435 ) ? ( VREG_16_10 ) : ( n23967 ) ;
assign n23969 =  ( n23434 ) ? ( VREG_16_11 ) : ( n23968 ) ;
assign n23970 =  ( n23433 ) ? ( VREG_16_12 ) : ( n23969 ) ;
assign n23971 =  ( n23432 ) ? ( VREG_16_13 ) : ( n23970 ) ;
assign n23972 =  ( n23431 ) ? ( VREG_16_14 ) : ( n23971 ) ;
assign n23973 =  ( n23430 ) ? ( VREG_16_15 ) : ( n23972 ) ;
assign n23974 =  ( n23429 ) ? ( VREG_17_0 ) : ( n23973 ) ;
assign n23975 =  ( n23428 ) ? ( VREG_17_1 ) : ( n23974 ) ;
assign n23976 =  ( n23427 ) ? ( VREG_17_2 ) : ( n23975 ) ;
assign n23977 =  ( n23426 ) ? ( VREG_17_3 ) : ( n23976 ) ;
assign n23978 =  ( n23425 ) ? ( VREG_17_4 ) : ( n23977 ) ;
assign n23979 =  ( n23424 ) ? ( VREG_17_5 ) : ( n23978 ) ;
assign n23980 =  ( n23423 ) ? ( VREG_17_6 ) : ( n23979 ) ;
assign n23981 =  ( n23422 ) ? ( VREG_17_7 ) : ( n23980 ) ;
assign n23982 =  ( n23421 ) ? ( VREG_17_8 ) : ( n23981 ) ;
assign n23983 =  ( n23420 ) ? ( VREG_17_9 ) : ( n23982 ) ;
assign n23984 =  ( n23419 ) ? ( VREG_17_10 ) : ( n23983 ) ;
assign n23985 =  ( n23418 ) ? ( VREG_17_11 ) : ( n23984 ) ;
assign n23986 =  ( n23417 ) ? ( VREG_17_12 ) : ( n23985 ) ;
assign n23987 =  ( n23416 ) ? ( VREG_17_13 ) : ( n23986 ) ;
assign n23988 =  ( n23415 ) ? ( VREG_17_14 ) : ( n23987 ) ;
assign n23989 =  ( n23414 ) ? ( VREG_17_15 ) : ( n23988 ) ;
assign n23990 =  ( n23413 ) ? ( VREG_18_0 ) : ( n23989 ) ;
assign n23991 =  ( n23412 ) ? ( VREG_18_1 ) : ( n23990 ) ;
assign n23992 =  ( n23411 ) ? ( VREG_18_2 ) : ( n23991 ) ;
assign n23993 =  ( n23410 ) ? ( VREG_18_3 ) : ( n23992 ) ;
assign n23994 =  ( n23409 ) ? ( VREG_18_4 ) : ( n23993 ) ;
assign n23995 =  ( n23408 ) ? ( VREG_18_5 ) : ( n23994 ) ;
assign n23996 =  ( n23407 ) ? ( VREG_18_6 ) : ( n23995 ) ;
assign n23997 =  ( n23406 ) ? ( VREG_18_7 ) : ( n23996 ) ;
assign n23998 =  ( n23405 ) ? ( VREG_18_8 ) : ( n23997 ) ;
assign n23999 =  ( n23404 ) ? ( VREG_18_9 ) : ( n23998 ) ;
assign n24000 =  ( n23403 ) ? ( VREG_18_10 ) : ( n23999 ) ;
assign n24001 =  ( n23402 ) ? ( VREG_18_11 ) : ( n24000 ) ;
assign n24002 =  ( n23401 ) ? ( VREG_18_12 ) : ( n24001 ) ;
assign n24003 =  ( n23400 ) ? ( VREG_18_13 ) : ( n24002 ) ;
assign n24004 =  ( n23399 ) ? ( VREG_18_14 ) : ( n24003 ) ;
assign n24005 =  ( n23398 ) ? ( VREG_18_15 ) : ( n24004 ) ;
assign n24006 =  ( n23397 ) ? ( VREG_19_0 ) : ( n24005 ) ;
assign n24007 =  ( n23396 ) ? ( VREG_19_1 ) : ( n24006 ) ;
assign n24008 =  ( n23395 ) ? ( VREG_19_2 ) : ( n24007 ) ;
assign n24009 =  ( n23394 ) ? ( VREG_19_3 ) : ( n24008 ) ;
assign n24010 =  ( n23393 ) ? ( VREG_19_4 ) : ( n24009 ) ;
assign n24011 =  ( n23392 ) ? ( VREG_19_5 ) : ( n24010 ) ;
assign n24012 =  ( n23391 ) ? ( VREG_19_6 ) : ( n24011 ) ;
assign n24013 =  ( n23390 ) ? ( VREG_19_7 ) : ( n24012 ) ;
assign n24014 =  ( n23389 ) ? ( VREG_19_8 ) : ( n24013 ) ;
assign n24015 =  ( n23388 ) ? ( VREG_19_9 ) : ( n24014 ) ;
assign n24016 =  ( n23387 ) ? ( VREG_19_10 ) : ( n24015 ) ;
assign n24017 =  ( n23386 ) ? ( VREG_19_11 ) : ( n24016 ) ;
assign n24018 =  ( n23385 ) ? ( VREG_19_12 ) : ( n24017 ) ;
assign n24019 =  ( n23384 ) ? ( VREG_19_13 ) : ( n24018 ) ;
assign n24020 =  ( n23383 ) ? ( VREG_19_14 ) : ( n24019 ) ;
assign n24021 =  ( n23382 ) ? ( VREG_19_15 ) : ( n24020 ) ;
assign n24022 =  ( n23381 ) ? ( VREG_20_0 ) : ( n24021 ) ;
assign n24023 =  ( n23380 ) ? ( VREG_20_1 ) : ( n24022 ) ;
assign n24024 =  ( n23379 ) ? ( VREG_20_2 ) : ( n24023 ) ;
assign n24025 =  ( n23378 ) ? ( VREG_20_3 ) : ( n24024 ) ;
assign n24026 =  ( n23377 ) ? ( VREG_20_4 ) : ( n24025 ) ;
assign n24027 =  ( n23376 ) ? ( VREG_20_5 ) : ( n24026 ) ;
assign n24028 =  ( n23375 ) ? ( VREG_20_6 ) : ( n24027 ) ;
assign n24029 =  ( n23374 ) ? ( VREG_20_7 ) : ( n24028 ) ;
assign n24030 =  ( n23373 ) ? ( VREG_20_8 ) : ( n24029 ) ;
assign n24031 =  ( n23372 ) ? ( VREG_20_9 ) : ( n24030 ) ;
assign n24032 =  ( n23371 ) ? ( VREG_20_10 ) : ( n24031 ) ;
assign n24033 =  ( n23370 ) ? ( VREG_20_11 ) : ( n24032 ) ;
assign n24034 =  ( n23369 ) ? ( VREG_20_12 ) : ( n24033 ) ;
assign n24035 =  ( n23368 ) ? ( VREG_20_13 ) : ( n24034 ) ;
assign n24036 =  ( n23367 ) ? ( VREG_20_14 ) : ( n24035 ) ;
assign n24037 =  ( n23366 ) ? ( VREG_20_15 ) : ( n24036 ) ;
assign n24038 =  ( n23365 ) ? ( VREG_21_0 ) : ( n24037 ) ;
assign n24039 =  ( n23364 ) ? ( VREG_21_1 ) : ( n24038 ) ;
assign n24040 =  ( n23363 ) ? ( VREG_21_2 ) : ( n24039 ) ;
assign n24041 =  ( n23362 ) ? ( VREG_21_3 ) : ( n24040 ) ;
assign n24042 =  ( n23361 ) ? ( VREG_21_4 ) : ( n24041 ) ;
assign n24043 =  ( n23360 ) ? ( VREG_21_5 ) : ( n24042 ) ;
assign n24044 =  ( n23359 ) ? ( VREG_21_6 ) : ( n24043 ) ;
assign n24045 =  ( n23358 ) ? ( VREG_21_7 ) : ( n24044 ) ;
assign n24046 =  ( n23357 ) ? ( VREG_21_8 ) : ( n24045 ) ;
assign n24047 =  ( n23356 ) ? ( VREG_21_9 ) : ( n24046 ) ;
assign n24048 =  ( n23355 ) ? ( VREG_21_10 ) : ( n24047 ) ;
assign n24049 =  ( n23354 ) ? ( VREG_21_11 ) : ( n24048 ) ;
assign n24050 =  ( n23353 ) ? ( VREG_21_12 ) : ( n24049 ) ;
assign n24051 =  ( n23352 ) ? ( VREG_21_13 ) : ( n24050 ) ;
assign n24052 =  ( n23351 ) ? ( VREG_21_14 ) : ( n24051 ) ;
assign n24053 =  ( n23350 ) ? ( VREG_21_15 ) : ( n24052 ) ;
assign n24054 =  ( n23349 ) ? ( VREG_22_0 ) : ( n24053 ) ;
assign n24055 =  ( n23348 ) ? ( VREG_22_1 ) : ( n24054 ) ;
assign n24056 =  ( n23347 ) ? ( VREG_22_2 ) : ( n24055 ) ;
assign n24057 =  ( n23346 ) ? ( VREG_22_3 ) : ( n24056 ) ;
assign n24058 =  ( n23345 ) ? ( VREG_22_4 ) : ( n24057 ) ;
assign n24059 =  ( n23344 ) ? ( VREG_22_5 ) : ( n24058 ) ;
assign n24060 =  ( n23343 ) ? ( VREG_22_6 ) : ( n24059 ) ;
assign n24061 =  ( n23342 ) ? ( VREG_22_7 ) : ( n24060 ) ;
assign n24062 =  ( n23341 ) ? ( VREG_22_8 ) : ( n24061 ) ;
assign n24063 =  ( n23340 ) ? ( VREG_22_9 ) : ( n24062 ) ;
assign n24064 =  ( n23339 ) ? ( VREG_22_10 ) : ( n24063 ) ;
assign n24065 =  ( n23338 ) ? ( VREG_22_11 ) : ( n24064 ) ;
assign n24066 =  ( n23337 ) ? ( VREG_22_12 ) : ( n24065 ) ;
assign n24067 =  ( n23336 ) ? ( VREG_22_13 ) : ( n24066 ) ;
assign n24068 =  ( n23335 ) ? ( VREG_22_14 ) : ( n24067 ) ;
assign n24069 =  ( n23334 ) ? ( VREG_22_15 ) : ( n24068 ) ;
assign n24070 =  ( n23333 ) ? ( VREG_23_0 ) : ( n24069 ) ;
assign n24071 =  ( n23332 ) ? ( VREG_23_1 ) : ( n24070 ) ;
assign n24072 =  ( n23331 ) ? ( VREG_23_2 ) : ( n24071 ) ;
assign n24073 =  ( n23330 ) ? ( VREG_23_3 ) : ( n24072 ) ;
assign n24074 =  ( n23329 ) ? ( VREG_23_4 ) : ( n24073 ) ;
assign n24075 =  ( n23328 ) ? ( VREG_23_5 ) : ( n24074 ) ;
assign n24076 =  ( n23327 ) ? ( VREG_23_6 ) : ( n24075 ) ;
assign n24077 =  ( n23326 ) ? ( VREG_23_7 ) : ( n24076 ) ;
assign n24078 =  ( n23325 ) ? ( VREG_23_8 ) : ( n24077 ) ;
assign n24079 =  ( n23324 ) ? ( VREG_23_9 ) : ( n24078 ) ;
assign n24080 =  ( n23323 ) ? ( VREG_23_10 ) : ( n24079 ) ;
assign n24081 =  ( n23322 ) ? ( VREG_23_11 ) : ( n24080 ) ;
assign n24082 =  ( n23321 ) ? ( VREG_23_12 ) : ( n24081 ) ;
assign n24083 =  ( n23320 ) ? ( VREG_23_13 ) : ( n24082 ) ;
assign n24084 =  ( n23319 ) ? ( VREG_23_14 ) : ( n24083 ) ;
assign n24085 =  ( n23318 ) ? ( VREG_23_15 ) : ( n24084 ) ;
assign n24086 =  ( n23317 ) ? ( VREG_24_0 ) : ( n24085 ) ;
assign n24087 =  ( n23316 ) ? ( VREG_24_1 ) : ( n24086 ) ;
assign n24088 =  ( n23315 ) ? ( VREG_24_2 ) : ( n24087 ) ;
assign n24089 =  ( n23314 ) ? ( VREG_24_3 ) : ( n24088 ) ;
assign n24090 =  ( n23313 ) ? ( VREG_24_4 ) : ( n24089 ) ;
assign n24091 =  ( n23312 ) ? ( VREG_24_5 ) : ( n24090 ) ;
assign n24092 =  ( n23311 ) ? ( VREG_24_6 ) : ( n24091 ) ;
assign n24093 =  ( n23310 ) ? ( VREG_24_7 ) : ( n24092 ) ;
assign n24094 =  ( n23309 ) ? ( VREG_24_8 ) : ( n24093 ) ;
assign n24095 =  ( n23308 ) ? ( VREG_24_9 ) : ( n24094 ) ;
assign n24096 =  ( n23307 ) ? ( VREG_24_10 ) : ( n24095 ) ;
assign n24097 =  ( n23306 ) ? ( VREG_24_11 ) : ( n24096 ) ;
assign n24098 =  ( n23305 ) ? ( VREG_24_12 ) : ( n24097 ) ;
assign n24099 =  ( n23304 ) ? ( VREG_24_13 ) : ( n24098 ) ;
assign n24100 =  ( n23303 ) ? ( VREG_24_14 ) : ( n24099 ) ;
assign n24101 =  ( n23302 ) ? ( VREG_24_15 ) : ( n24100 ) ;
assign n24102 =  ( n23301 ) ? ( VREG_25_0 ) : ( n24101 ) ;
assign n24103 =  ( n23300 ) ? ( VREG_25_1 ) : ( n24102 ) ;
assign n24104 =  ( n23299 ) ? ( VREG_25_2 ) : ( n24103 ) ;
assign n24105 =  ( n23298 ) ? ( VREG_25_3 ) : ( n24104 ) ;
assign n24106 =  ( n23297 ) ? ( VREG_25_4 ) : ( n24105 ) ;
assign n24107 =  ( n23296 ) ? ( VREG_25_5 ) : ( n24106 ) ;
assign n24108 =  ( n23295 ) ? ( VREG_25_6 ) : ( n24107 ) ;
assign n24109 =  ( n23294 ) ? ( VREG_25_7 ) : ( n24108 ) ;
assign n24110 =  ( n23293 ) ? ( VREG_25_8 ) : ( n24109 ) ;
assign n24111 =  ( n23292 ) ? ( VREG_25_9 ) : ( n24110 ) ;
assign n24112 =  ( n23291 ) ? ( VREG_25_10 ) : ( n24111 ) ;
assign n24113 =  ( n23290 ) ? ( VREG_25_11 ) : ( n24112 ) ;
assign n24114 =  ( n23289 ) ? ( VREG_25_12 ) : ( n24113 ) ;
assign n24115 =  ( n23288 ) ? ( VREG_25_13 ) : ( n24114 ) ;
assign n24116 =  ( n23287 ) ? ( VREG_25_14 ) : ( n24115 ) ;
assign n24117 =  ( n23286 ) ? ( VREG_25_15 ) : ( n24116 ) ;
assign n24118 =  ( n23285 ) ? ( VREG_26_0 ) : ( n24117 ) ;
assign n24119 =  ( n23284 ) ? ( VREG_26_1 ) : ( n24118 ) ;
assign n24120 =  ( n23283 ) ? ( VREG_26_2 ) : ( n24119 ) ;
assign n24121 =  ( n23282 ) ? ( VREG_26_3 ) : ( n24120 ) ;
assign n24122 =  ( n23281 ) ? ( VREG_26_4 ) : ( n24121 ) ;
assign n24123 =  ( n23280 ) ? ( VREG_26_5 ) : ( n24122 ) ;
assign n24124 =  ( n23279 ) ? ( VREG_26_6 ) : ( n24123 ) ;
assign n24125 =  ( n23278 ) ? ( VREG_26_7 ) : ( n24124 ) ;
assign n24126 =  ( n23277 ) ? ( VREG_26_8 ) : ( n24125 ) ;
assign n24127 =  ( n23276 ) ? ( VREG_26_9 ) : ( n24126 ) ;
assign n24128 =  ( n23275 ) ? ( VREG_26_10 ) : ( n24127 ) ;
assign n24129 =  ( n23274 ) ? ( VREG_26_11 ) : ( n24128 ) ;
assign n24130 =  ( n23273 ) ? ( VREG_26_12 ) : ( n24129 ) ;
assign n24131 =  ( n23272 ) ? ( VREG_26_13 ) : ( n24130 ) ;
assign n24132 =  ( n23271 ) ? ( VREG_26_14 ) : ( n24131 ) ;
assign n24133 =  ( n23270 ) ? ( VREG_26_15 ) : ( n24132 ) ;
assign n24134 =  ( n23269 ) ? ( VREG_27_0 ) : ( n24133 ) ;
assign n24135 =  ( n23268 ) ? ( VREG_27_1 ) : ( n24134 ) ;
assign n24136 =  ( n23267 ) ? ( VREG_27_2 ) : ( n24135 ) ;
assign n24137 =  ( n23266 ) ? ( VREG_27_3 ) : ( n24136 ) ;
assign n24138 =  ( n23265 ) ? ( VREG_27_4 ) : ( n24137 ) ;
assign n24139 =  ( n23264 ) ? ( VREG_27_5 ) : ( n24138 ) ;
assign n24140 =  ( n23263 ) ? ( VREG_27_6 ) : ( n24139 ) ;
assign n24141 =  ( n23262 ) ? ( VREG_27_7 ) : ( n24140 ) ;
assign n24142 =  ( n23261 ) ? ( VREG_27_8 ) : ( n24141 ) ;
assign n24143 =  ( n23260 ) ? ( VREG_27_9 ) : ( n24142 ) ;
assign n24144 =  ( n23259 ) ? ( VREG_27_10 ) : ( n24143 ) ;
assign n24145 =  ( n23258 ) ? ( VREG_27_11 ) : ( n24144 ) ;
assign n24146 =  ( n23257 ) ? ( VREG_27_12 ) : ( n24145 ) ;
assign n24147 =  ( n23256 ) ? ( VREG_27_13 ) : ( n24146 ) ;
assign n24148 =  ( n23255 ) ? ( VREG_27_14 ) : ( n24147 ) ;
assign n24149 =  ( n23254 ) ? ( VREG_27_15 ) : ( n24148 ) ;
assign n24150 =  ( n23253 ) ? ( VREG_28_0 ) : ( n24149 ) ;
assign n24151 =  ( n23252 ) ? ( VREG_28_1 ) : ( n24150 ) ;
assign n24152 =  ( n23251 ) ? ( VREG_28_2 ) : ( n24151 ) ;
assign n24153 =  ( n23250 ) ? ( VREG_28_3 ) : ( n24152 ) ;
assign n24154 =  ( n23249 ) ? ( VREG_28_4 ) : ( n24153 ) ;
assign n24155 =  ( n23248 ) ? ( VREG_28_5 ) : ( n24154 ) ;
assign n24156 =  ( n23247 ) ? ( VREG_28_6 ) : ( n24155 ) ;
assign n24157 =  ( n23246 ) ? ( VREG_28_7 ) : ( n24156 ) ;
assign n24158 =  ( n23245 ) ? ( VREG_28_8 ) : ( n24157 ) ;
assign n24159 =  ( n23244 ) ? ( VREG_28_9 ) : ( n24158 ) ;
assign n24160 =  ( n23243 ) ? ( VREG_28_10 ) : ( n24159 ) ;
assign n24161 =  ( n23242 ) ? ( VREG_28_11 ) : ( n24160 ) ;
assign n24162 =  ( n23241 ) ? ( VREG_28_12 ) : ( n24161 ) ;
assign n24163 =  ( n23240 ) ? ( VREG_28_13 ) : ( n24162 ) ;
assign n24164 =  ( n23239 ) ? ( VREG_28_14 ) : ( n24163 ) ;
assign n24165 =  ( n23238 ) ? ( VREG_28_15 ) : ( n24164 ) ;
assign n24166 =  ( n23237 ) ? ( VREG_29_0 ) : ( n24165 ) ;
assign n24167 =  ( n23236 ) ? ( VREG_29_1 ) : ( n24166 ) ;
assign n24168 =  ( n23235 ) ? ( VREG_29_2 ) : ( n24167 ) ;
assign n24169 =  ( n23234 ) ? ( VREG_29_3 ) : ( n24168 ) ;
assign n24170 =  ( n23233 ) ? ( VREG_29_4 ) : ( n24169 ) ;
assign n24171 =  ( n23232 ) ? ( VREG_29_5 ) : ( n24170 ) ;
assign n24172 =  ( n23231 ) ? ( VREG_29_6 ) : ( n24171 ) ;
assign n24173 =  ( n23230 ) ? ( VREG_29_7 ) : ( n24172 ) ;
assign n24174 =  ( n23229 ) ? ( VREG_29_8 ) : ( n24173 ) ;
assign n24175 =  ( n23228 ) ? ( VREG_29_9 ) : ( n24174 ) ;
assign n24176 =  ( n23227 ) ? ( VREG_29_10 ) : ( n24175 ) ;
assign n24177 =  ( n23226 ) ? ( VREG_29_11 ) : ( n24176 ) ;
assign n24178 =  ( n23225 ) ? ( VREG_29_12 ) : ( n24177 ) ;
assign n24179 =  ( n23224 ) ? ( VREG_29_13 ) : ( n24178 ) ;
assign n24180 =  ( n23223 ) ? ( VREG_29_14 ) : ( n24179 ) ;
assign n24181 =  ( n23222 ) ? ( VREG_29_15 ) : ( n24180 ) ;
assign n24182 =  ( n23221 ) ? ( VREG_30_0 ) : ( n24181 ) ;
assign n24183 =  ( n23220 ) ? ( VREG_30_1 ) : ( n24182 ) ;
assign n24184 =  ( n23219 ) ? ( VREG_30_2 ) : ( n24183 ) ;
assign n24185 =  ( n23218 ) ? ( VREG_30_3 ) : ( n24184 ) ;
assign n24186 =  ( n23217 ) ? ( VREG_30_4 ) : ( n24185 ) ;
assign n24187 =  ( n23216 ) ? ( VREG_30_5 ) : ( n24186 ) ;
assign n24188 =  ( n23215 ) ? ( VREG_30_6 ) : ( n24187 ) ;
assign n24189 =  ( n23214 ) ? ( VREG_30_7 ) : ( n24188 ) ;
assign n24190 =  ( n23213 ) ? ( VREG_30_8 ) : ( n24189 ) ;
assign n24191 =  ( n23212 ) ? ( VREG_30_9 ) : ( n24190 ) ;
assign n24192 =  ( n23211 ) ? ( VREG_30_10 ) : ( n24191 ) ;
assign n24193 =  ( n23210 ) ? ( VREG_30_11 ) : ( n24192 ) ;
assign n24194 =  ( n23209 ) ? ( VREG_30_12 ) : ( n24193 ) ;
assign n24195 =  ( n23208 ) ? ( VREG_30_13 ) : ( n24194 ) ;
assign n24196 =  ( n23207 ) ? ( VREG_30_14 ) : ( n24195 ) ;
assign n24197 =  ( n23206 ) ? ( VREG_30_15 ) : ( n24196 ) ;
assign n24198 =  ( n23205 ) ? ( VREG_31_0 ) : ( n24197 ) ;
assign n24199 =  ( n23204 ) ? ( VREG_31_1 ) : ( n24198 ) ;
assign n24200 =  ( n23203 ) ? ( VREG_31_2 ) : ( n24199 ) ;
assign n24201 =  ( n23202 ) ? ( VREG_31_3 ) : ( n24200 ) ;
assign n24202 =  ( n23201 ) ? ( VREG_31_4 ) : ( n24201 ) ;
assign n24203 =  ( n23200 ) ? ( VREG_31_5 ) : ( n24202 ) ;
assign n24204 =  ( n23199 ) ? ( VREG_31_6 ) : ( n24203 ) ;
assign n24205 =  ( n23198 ) ? ( VREG_31_7 ) : ( n24204 ) ;
assign n24206 =  ( n23197 ) ? ( VREG_31_8 ) : ( n24205 ) ;
assign n24207 =  ( n23196 ) ? ( VREG_31_9 ) : ( n24206 ) ;
assign n24208 =  ( n23195 ) ? ( VREG_31_10 ) : ( n24207 ) ;
assign n24209 =  ( n23194 ) ? ( VREG_31_11 ) : ( n24208 ) ;
assign n24210 =  ( n23193 ) ? ( VREG_31_12 ) : ( n24209 ) ;
assign n24211 =  ( n23192 ) ? ( VREG_31_13 ) : ( n24210 ) ;
assign n24212 =  ( n23191 ) ? ( VREG_31_14 ) : ( n24211 ) ;
assign n24213 =  ( n23190 ) ? ( VREG_31_15 ) : ( n24212 ) ;
assign n24214 =  ( n23179 ) + ( n24213 )  ;
assign n24215 =  ( n23179 ) - ( n24213 )  ;
assign n24216 =  ( n23179 ) & ( n24213 )  ;
assign n24217 =  ( n23179 ) | ( n24213 )  ;
assign n24218 =  ( ( n23179 ) * ( n24213 ))  ;
assign n24219 =  ( n148 ) ? ( n24218 ) : ( VREG_0_4 ) ;
assign n24220 =  ( n146 ) ? ( n24217 ) : ( n24219 ) ;
assign n24221 =  ( n144 ) ? ( n24216 ) : ( n24220 ) ;
assign n24222 =  ( n142 ) ? ( n24215 ) : ( n24221 ) ;
assign n24223 =  ( n10 ) ? ( n24214 ) : ( n24222 ) ;
assign n24224 = n3030[4:4] ;
assign n24225 =  ( n24224 ) == ( 1'd0 )  ;
assign n24226 =  ( n24225 ) ? ( VREG_0_4 ) : ( n23189 ) ;
assign n24227 =  ( n24225 ) ? ( VREG_0_4 ) : ( n24223 ) ;
assign n24228 =  ( n3034 ) ? ( n24227 ) : ( VREG_0_4 ) ;
assign n24229 =  ( n2965 ) ? ( n24226 ) : ( n24228 ) ;
assign n24230 =  ( n1930 ) ? ( n24223 ) : ( n24229 ) ;
assign n24231 =  ( n879 ) ? ( n23189 ) : ( n24230 ) ;
assign n24232 =  ( n23179 ) + ( n164 )  ;
assign n24233 =  ( n23179 ) - ( n164 )  ;
assign n24234 =  ( n23179 ) & ( n164 )  ;
assign n24235 =  ( n23179 ) | ( n164 )  ;
assign n24236 =  ( ( n23179 ) * ( n164 ))  ;
assign n24237 =  ( n172 ) ? ( n24236 ) : ( VREG_0_4 ) ;
assign n24238 =  ( n170 ) ? ( n24235 ) : ( n24237 ) ;
assign n24239 =  ( n168 ) ? ( n24234 ) : ( n24238 ) ;
assign n24240 =  ( n166 ) ? ( n24233 ) : ( n24239 ) ;
assign n24241 =  ( n162 ) ? ( n24232 ) : ( n24240 ) ;
assign n24242 =  ( n23179 ) + ( n180 )  ;
assign n24243 =  ( n23179 ) - ( n180 )  ;
assign n24244 =  ( n23179 ) & ( n180 )  ;
assign n24245 =  ( n23179 ) | ( n180 )  ;
assign n24246 =  ( ( n23179 ) * ( n180 ))  ;
assign n24247 =  ( n172 ) ? ( n24246 ) : ( VREG_0_4 ) ;
assign n24248 =  ( n170 ) ? ( n24245 ) : ( n24247 ) ;
assign n24249 =  ( n168 ) ? ( n24244 ) : ( n24248 ) ;
assign n24250 =  ( n166 ) ? ( n24243 ) : ( n24249 ) ;
assign n24251 =  ( n162 ) ? ( n24242 ) : ( n24250 ) ;
assign n24252 =  ( n24225 ) ? ( VREG_0_4 ) : ( n24251 ) ;
assign n24253 =  ( n3051 ) ? ( n24252 ) : ( VREG_0_4 ) ;
assign n24254 =  ( n3040 ) ? ( n24241 ) : ( n24253 ) ;
assign n24255 =  ( n192 ) ? ( VREG_0_4 ) : ( VREG_0_4 ) ;
assign n24256 =  ( n157 ) ? ( n24254 ) : ( n24255 ) ;
assign n24257 =  ( n6 ) ? ( n24231 ) : ( n24256 ) ;
assign n24258 =  ( n4 ) ? ( n24257 ) : ( VREG_0_4 ) ;
assign n24259 =  ( 32'd5 ) == ( 32'd15 )  ;
assign n24260 =  ( n12 ) & ( n24259 )  ;
assign n24261 =  ( 32'd5 ) == ( 32'd14 )  ;
assign n24262 =  ( n12 ) & ( n24261 )  ;
assign n24263 =  ( 32'd5 ) == ( 32'd13 )  ;
assign n24264 =  ( n12 ) & ( n24263 )  ;
assign n24265 =  ( 32'd5 ) == ( 32'd12 )  ;
assign n24266 =  ( n12 ) & ( n24265 )  ;
assign n24267 =  ( 32'd5 ) == ( 32'd11 )  ;
assign n24268 =  ( n12 ) & ( n24267 )  ;
assign n24269 =  ( 32'd5 ) == ( 32'd10 )  ;
assign n24270 =  ( n12 ) & ( n24269 )  ;
assign n24271 =  ( 32'd5 ) == ( 32'd9 )  ;
assign n24272 =  ( n12 ) & ( n24271 )  ;
assign n24273 =  ( 32'd5 ) == ( 32'd8 )  ;
assign n24274 =  ( n12 ) & ( n24273 )  ;
assign n24275 =  ( 32'd5 ) == ( 32'd7 )  ;
assign n24276 =  ( n12 ) & ( n24275 )  ;
assign n24277 =  ( 32'd5 ) == ( 32'd6 )  ;
assign n24278 =  ( n12 ) & ( n24277 )  ;
assign n24279 =  ( 32'd5 ) == ( 32'd5 )  ;
assign n24280 =  ( n12 ) & ( n24279 )  ;
assign n24281 =  ( 32'd5 ) == ( 32'd4 )  ;
assign n24282 =  ( n12 ) & ( n24281 )  ;
assign n24283 =  ( 32'd5 ) == ( 32'd3 )  ;
assign n24284 =  ( n12 ) & ( n24283 )  ;
assign n24285 =  ( 32'd5 ) == ( 32'd2 )  ;
assign n24286 =  ( n12 ) & ( n24285 )  ;
assign n24287 =  ( 32'd5 ) == ( 32'd1 )  ;
assign n24288 =  ( n12 ) & ( n24287 )  ;
assign n24289 =  ( 32'd5 ) == ( 32'd0 )  ;
assign n24290 =  ( n12 ) & ( n24289 )  ;
assign n24291 =  ( n13 ) & ( n24259 )  ;
assign n24292 =  ( n13 ) & ( n24261 )  ;
assign n24293 =  ( n13 ) & ( n24263 )  ;
assign n24294 =  ( n13 ) & ( n24265 )  ;
assign n24295 =  ( n13 ) & ( n24267 )  ;
assign n24296 =  ( n13 ) & ( n24269 )  ;
assign n24297 =  ( n13 ) & ( n24271 )  ;
assign n24298 =  ( n13 ) & ( n24273 )  ;
assign n24299 =  ( n13 ) & ( n24275 )  ;
assign n24300 =  ( n13 ) & ( n24277 )  ;
assign n24301 =  ( n13 ) & ( n24279 )  ;
assign n24302 =  ( n13 ) & ( n24281 )  ;
assign n24303 =  ( n13 ) & ( n24283 )  ;
assign n24304 =  ( n13 ) & ( n24285 )  ;
assign n24305 =  ( n13 ) & ( n24287 )  ;
assign n24306 =  ( n13 ) & ( n24289 )  ;
assign n24307 =  ( n14 ) & ( n24259 )  ;
assign n24308 =  ( n14 ) & ( n24261 )  ;
assign n24309 =  ( n14 ) & ( n24263 )  ;
assign n24310 =  ( n14 ) & ( n24265 )  ;
assign n24311 =  ( n14 ) & ( n24267 )  ;
assign n24312 =  ( n14 ) & ( n24269 )  ;
assign n24313 =  ( n14 ) & ( n24271 )  ;
assign n24314 =  ( n14 ) & ( n24273 )  ;
assign n24315 =  ( n14 ) & ( n24275 )  ;
assign n24316 =  ( n14 ) & ( n24277 )  ;
assign n24317 =  ( n14 ) & ( n24279 )  ;
assign n24318 =  ( n14 ) & ( n24281 )  ;
assign n24319 =  ( n14 ) & ( n24283 )  ;
assign n24320 =  ( n14 ) & ( n24285 )  ;
assign n24321 =  ( n14 ) & ( n24287 )  ;
assign n24322 =  ( n14 ) & ( n24289 )  ;
assign n24323 =  ( n15 ) & ( n24259 )  ;
assign n24324 =  ( n15 ) & ( n24261 )  ;
assign n24325 =  ( n15 ) & ( n24263 )  ;
assign n24326 =  ( n15 ) & ( n24265 )  ;
assign n24327 =  ( n15 ) & ( n24267 )  ;
assign n24328 =  ( n15 ) & ( n24269 )  ;
assign n24329 =  ( n15 ) & ( n24271 )  ;
assign n24330 =  ( n15 ) & ( n24273 )  ;
assign n24331 =  ( n15 ) & ( n24275 )  ;
assign n24332 =  ( n15 ) & ( n24277 )  ;
assign n24333 =  ( n15 ) & ( n24279 )  ;
assign n24334 =  ( n15 ) & ( n24281 )  ;
assign n24335 =  ( n15 ) & ( n24283 )  ;
assign n24336 =  ( n15 ) & ( n24285 )  ;
assign n24337 =  ( n15 ) & ( n24287 )  ;
assign n24338 =  ( n15 ) & ( n24289 )  ;
assign n24339 =  ( n16 ) & ( n24259 )  ;
assign n24340 =  ( n16 ) & ( n24261 )  ;
assign n24341 =  ( n16 ) & ( n24263 )  ;
assign n24342 =  ( n16 ) & ( n24265 )  ;
assign n24343 =  ( n16 ) & ( n24267 )  ;
assign n24344 =  ( n16 ) & ( n24269 )  ;
assign n24345 =  ( n16 ) & ( n24271 )  ;
assign n24346 =  ( n16 ) & ( n24273 )  ;
assign n24347 =  ( n16 ) & ( n24275 )  ;
assign n24348 =  ( n16 ) & ( n24277 )  ;
assign n24349 =  ( n16 ) & ( n24279 )  ;
assign n24350 =  ( n16 ) & ( n24281 )  ;
assign n24351 =  ( n16 ) & ( n24283 )  ;
assign n24352 =  ( n16 ) & ( n24285 )  ;
assign n24353 =  ( n16 ) & ( n24287 )  ;
assign n24354 =  ( n16 ) & ( n24289 )  ;
assign n24355 =  ( n17 ) & ( n24259 )  ;
assign n24356 =  ( n17 ) & ( n24261 )  ;
assign n24357 =  ( n17 ) & ( n24263 )  ;
assign n24358 =  ( n17 ) & ( n24265 )  ;
assign n24359 =  ( n17 ) & ( n24267 )  ;
assign n24360 =  ( n17 ) & ( n24269 )  ;
assign n24361 =  ( n17 ) & ( n24271 )  ;
assign n24362 =  ( n17 ) & ( n24273 )  ;
assign n24363 =  ( n17 ) & ( n24275 )  ;
assign n24364 =  ( n17 ) & ( n24277 )  ;
assign n24365 =  ( n17 ) & ( n24279 )  ;
assign n24366 =  ( n17 ) & ( n24281 )  ;
assign n24367 =  ( n17 ) & ( n24283 )  ;
assign n24368 =  ( n17 ) & ( n24285 )  ;
assign n24369 =  ( n17 ) & ( n24287 )  ;
assign n24370 =  ( n17 ) & ( n24289 )  ;
assign n24371 =  ( n18 ) & ( n24259 )  ;
assign n24372 =  ( n18 ) & ( n24261 )  ;
assign n24373 =  ( n18 ) & ( n24263 )  ;
assign n24374 =  ( n18 ) & ( n24265 )  ;
assign n24375 =  ( n18 ) & ( n24267 )  ;
assign n24376 =  ( n18 ) & ( n24269 )  ;
assign n24377 =  ( n18 ) & ( n24271 )  ;
assign n24378 =  ( n18 ) & ( n24273 )  ;
assign n24379 =  ( n18 ) & ( n24275 )  ;
assign n24380 =  ( n18 ) & ( n24277 )  ;
assign n24381 =  ( n18 ) & ( n24279 )  ;
assign n24382 =  ( n18 ) & ( n24281 )  ;
assign n24383 =  ( n18 ) & ( n24283 )  ;
assign n24384 =  ( n18 ) & ( n24285 )  ;
assign n24385 =  ( n18 ) & ( n24287 )  ;
assign n24386 =  ( n18 ) & ( n24289 )  ;
assign n24387 =  ( n19 ) & ( n24259 )  ;
assign n24388 =  ( n19 ) & ( n24261 )  ;
assign n24389 =  ( n19 ) & ( n24263 )  ;
assign n24390 =  ( n19 ) & ( n24265 )  ;
assign n24391 =  ( n19 ) & ( n24267 )  ;
assign n24392 =  ( n19 ) & ( n24269 )  ;
assign n24393 =  ( n19 ) & ( n24271 )  ;
assign n24394 =  ( n19 ) & ( n24273 )  ;
assign n24395 =  ( n19 ) & ( n24275 )  ;
assign n24396 =  ( n19 ) & ( n24277 )  ;
assign n24397 =  ( n19 ) & ( n24279 )  ;
assign n24398 =  ( n19 ) & ( n24281 )  ;
assign n24399 =  ( n19 ) & ( n24283 )  ;
assign n24400 =  ( n19 ) & ( n24285 )  ;
assign n24401 =  ( n19 ) & ( n24287 )  ;
assign n24402 =  ( n19 ) & ( n24289 )  ;
assign n24403 =  ( n20 ) & ( n24259 )  ;
assign n24404 =  ( n20 ) & ( n24261 )  ;
assign n24405 =  ( n20 ) & ( n24263 )  ;
assign n24406 =  ( n20 ) & ( n24265 )  ;
assign n24407 =  ( n20 ) & ( n24267 )  ;
assign n24408 =  ( n20 ) & ( n24269 )  ;
assign n24409 =  ( n20 ) & ( n24271 )  ;
assign n24410 =  ( n20 ) & ( n24273 )  ;
assign n24411 =  ( n20 ) & ( n24275 )  ;
assign n24412 =  ( n20 ) & ( n24277 )  ;
assign n24413 =  ( n20 ) & ( n24279 )  ;
assign n24414 =  ( n20 ) & ( n24281 )  ;
assign n24415 =  ( n20 ) & ( n24283 )  ;
assign n24416 =  ( n20 ) & ( n24285 )  ;
assign n24417 =  ( n20 ) & ( n24287 )  ;
assign n24418 =  ( n20 ) & ( n24289 )  ;
assign n24419 =  ( n21 ) & ( n24259 )  ;
assign n24420 =  ( n21 ) & ( n24261 )  ;
assign n24421 =  ( n21 ) & ( n24263 )  ;
assign n24422 =  ( n21 ) & ( n24265 )  ;
assign n24423 =  ( n21 ) & ( n24267 )  ;
assign n24424 =  ( n21 ) & ( n24269 )  ;
assign n24425 =  ( n21 ) & ( n24271 )  ;
assign n24426 =  ( n21 ) & ( n24273 )  ;
assign n24427 =  ( n21 ) & ( n24275 )  ;
assign n24428 =  ( n21 ) & ( n24277 )  ;
assign n24429 =  ( n21 ) & ( n24279 )  ;
assign n24430 =  ( n21 ) & ( n24281 )  ;
assign n24431 =  ( n21 ) & ( n24283 )  ;
assign n24432 =  ( n21 ) & ( n24285 )  ;
assign n24433 =  ( n21 ) & ( n24287 )  ;
assign n24434 =  ( n21 ) & ( n24289 )  ;
assign n24435 =  ( n22 ) & ( n24259 )  ;
assign n24436 =  ( n22 ) & ( n24261 )  ;
assign n24437 =  ( n22 ) & ( n24263 )  ;
assign n24438 =  ( n22 ) & ( n24265 )  ;
assign n24439 =  ( n22 ) & ( n24267 )  ;
assign n24440 =  ( n22 ) & ( n24269 )  ;
assign n24441 =  ( n22 ) & ( n24271 )  ;
assign n24442 =  ( n22 ) & ( n24273 )  ;
assign n24443 =  ( n22 ) & ( n24275 )  ;
assign n24444 =  ( n22 ) & ( n24277 )  ;
assign n24445 =  ( n22 ) & ( n24279 )  ;
assign n24446 =  ( n22 ) & ( n24281 )  ;
assign n24447 =  ( n22 ) & ( n24283 )  ;
assign n24448 =  ( n22 ) & ( n24285 )  ;
assign n24449 =  ( n22 ) & ( n24287 )  ;
assign n24450 =  ( n22 ) & ( n24289 )  ;
assign n24451 =  ( n23 ) & ( n24259 )  ;
assign n24452 =  ( n23 ) & ( n24261 )  ;
assign n24453 =  ( n23 ) & ( n24263 )  ;
assign n24454 =  ( n23 ) & ( n24265 )  ;
assign n24455 =  ( n23 ) & ( n24267 )  ;
assign n24456 =  ( n23 ) & ( n24269 )  ;
assign n24457 =  ( n23 ) & ( n24271 )  ;
assign n24458 =  ( n23 ) & ( n24273 )  ;
assign n24459 =  ( n23 ) & ( n24275 )  ;
assign n24460 =  ( n23 ) & ( n24277 )  ;
assign n24461 =  ( n23 ) & ( n24279 )  ;
assign n24462 =  ( n23 ) & ( n24281 )  ;
assign n24463 =  ( n23 ) & ( n24283 )  ;
assign n24464 =  ( n23 ) & ( n24285 )  ;
assign n24465 =  ( n23 ) & ( n24287 )  ;
assign n24466 =  ( n23 ) & ( n24289 )  ;
assign n24467 =  ( n24 ) & ( n24259 )  ;
assign n24468 =  ( n24 ) & ( n24261 )  ;
assign n24469 =  ( n24 ) & ( n24263 )  ;
assign n24470 =  ( n24 ) & ( n24265 )  ;
assign n24471 =  ( n24 ) & ( n24267 )  ;
assign n24472 =  ( n24 ) & ( n24269 )  ;
assign n24473 =  ( n24 ) & ( n24271 )  ;
assign n24474 =  ( n24 ) & ( n24273 )  ;
assign n24475 =  ( n24 ) & ( n24275 )  ;
assign n24476 =  ( n24 ) & ( n24277 )  ;
assign n24477 =  ( n24 ) & ( n24279 )  ;
assign n24478 =  ( n24 ) & ( n24281 )  ;
assign n24479 =  ( n24 ) & ( n24283 )  ;
assign n24480 =  ( n24 ) & ( n24285 )  ;
assign n24481 =  ( n24 ) & ( n24287 )  ;
assign n24482 =  ( n24 ) & ( n24289 )  ;
assign n24483 =  ( n25 ) & ( n24259 )  ;
assign n24484 =  ( n25 ) & ( n24261 )  ;
assign n24485 =  ( n25 ) & ( n24263 )  ;
assign n24486 =  ( n25 ) & ( n24265 )  ;
assign n24487 =  ( n25 ) & ( n24267 )  ;
assign n24488 =  ( n25 ) & ( n24269 )  ;
assign n24489 =  ( n25 ) & ( n24271 )  ;
assign n24490 =  ( n25 ) & ( n24273 )  ;
assign n24491 =  ( n25 ) & ( n24275 )  ;
assign n24492 =  ( n25 ) & ( n24277 )  ;
assign n24493 =  ( n25 ) & ( n24279 )  ;
assign n24494 =  ( n25 ) & ( n24281 )  ;
assign n24495 =  ( n25 ) & ( n24283 )  ;
assign n24496 =  ( n25 ) & ( n24285 )  ;
assign n24497 =  ( n25 ) & ( n24287 )  ;
assign n24498 =  ( n25 ) & ( n24289 )  ;
assign n24499 =  ( n26 ) & ( n24259 )  ;
assign n24500 =  ( n26 ) & ( n24261 )  ;
assign n24501 =  ( n26 ) & ( n24263 )  ;
assign n24502 =  ( n26 ) & ( n24265 )  ;
assign n24503 =  ( n26 ) & ( n24267 )  ;
assign n24504 =  ( n26 ) & ( n24269 )  ;
assign n24505 =  ( n26 ) & ( n24271 )  ;
assign n24506 =  ( n26 ) & ( n24273 )  ;
assign n24507 =  ( n26 ) & ( n24275 )  ;
assign n24508 =  ( n26 ) & ( n24277 )  ;
assign n24509 =  ( n26 ) & ( n24279 )  ;
assign n24510 =  ( n26 ) & ( n24281 )  ;
assign n24511 =  ( n26 ) & ( n24283 )  ;
assign n24512 =  ( n26 ) & ( n24285 )  ;
assign n24513 =  ( n26 ) & ( n24287 )  ;
assign n24514 =  ( n26 ) & ( n24289 )  ;
assign n24515 =  ( n27 ) & ( n24259 )  ;
assign n24516 =  ( n27 ) & ( n24261 )  ;
assign n24517 =  ( n27 ) & ( n24263 )  ;
assign n24518 =  ( n27 ) & ( n24265 )  ;
assign n24519 =  ( n27 ) & ( n24267 )  ;
assign n24520 =  ( n27 ) & ( n24269 )  ;
assign n24521 =  ( n27 ) & ( n24271 )  ;
assign n24522 =  ( n27 ) & ( n24273 )  ;
assign n24523 =  ( n27 ) & ( n24275 )  ;
assign n24524 =  ( n27 ) & ( n24277 )  ;
assign n24525 =  ( n27 ) & ( n24279 )  ;
assign n24526 =  ( n27 ) & ( n24281 )  ;
assign n24527 =  ( n27 ) & ( n24283 )  ;
assign n24528 =  ( n27 ) & ( n24285 )  ;
assign n24529 =  ( n27 ) & ( n24287 )  ;
assign n24530 =  ( n27 ) & ( n24289 )  ;
assign n24531 =  ( n28 ) & ( n24259 )  ;
assign n24532 =  ( n28 ) & ( n24261 )  ;
assign n24533 =  ( n28 ) & ( n24263 )  ;
assign n24534 =  ( n28 ) & ( n24265 )  ;
assign n24535 =  ( n28 ) & ( n24267 )  ;
assign n24536 =  ( n28 ) & ( n24269 )  ;
assign n24537 =  ( n28 ) & ( n24271 )  ;
assign n24538 =  ( n28 ) & ( n24273 )  ;
assign n24539 =  ( n28 ) & ( n24275 )  ;
assign n24540 =  ( n28 ) & ( n24277 )  ;
assign n24541 =  ( n28 ) & ( n24279 )  ;
assign n24542 =  ( n28 ) & ( n24281 )  ;
assign n24543 =  ( n28 ) & ( n24283 )  ;
assign n24544 =  ( n28 ) & ( n24285 )  ;
assign n24545 =  ( n28 ) & ( n24287 )  ;
assign n24546 =  ( n28 ) & ( n24289 )  ;
assign n24547 =  ( n29 ) & ( n24259 )  ;
assign n24548 =  ( n29 ) & ( n24261 )  ;
assign n24549 =  ( n29 ) & ( n24263 )  ;
assign n24550 =  ( n29 ) & ( n24265 )  ;
assign n24551 =  ( n29 ) & ( n24267 )  ;
assign n24552 =  ( n29 ) & ( n24269 )  ;
assign n24553 =  ( n29 ) & ( n24271 )  ;
assign n24554 =  ( n29 ) & ( n24273 )  ;
assign n24555 =  ( n29 ) & ( n24275 )  ;
assign n24556 =  ( n29 ) & ( n24277 )  ;
assign n24557 =  ( n29 ) & ( n24279 )  ;
assign n24558 =  ( n29 ) & ( n24281 )  ;
assign n24559 =  ( n29 ) & ( n24283 )  ;
assign n24560 =  ( n29 ) & ( n24285 )  ;
assign n24561 =  ( n29 ) & ( n24287 )  ;
assign n24562 =  ( n29 ) & ( n24289 )  ;
assign n24563 =  ( n30 ) & ( n24259 )  ;
assign n24564 =  ( n30 ) & ( n24261 )  ;
assign n24565 =  ( n30 ) & ( n24263 )  ;
assign n24566 =  ( n30 ) & ( n24265 )  ;
assign n24567 =  ( n30 ) & ( n24267 )  ;
assign n24568 =  ( n30 ) & ( n24269 )  ;
assign n24569 =  ( n30 ) & ( n24271 )  ;
assign n24570 =  ( n30 ) & ( n24273 )  ;
assign n24571 =  ( n30 ) & ( n24275 )  ;
assign n24572 =  ( n30 ) & ( n24277 )  ;
assign n24573 =  ( n30 ) & ( n24279 )  ;
assign n24574 =  ( n30 ) & ( n24281 )  ;
assign n24575 =  ( n30 ) & ( n24283 )  ;
assign n24576 =  ( n30 ) & ( n24285 )  ;
assign n24577 =  ( n30 ) & ( n24287 )  ;
assign n24578 =  ( n30 ) & ( n24289 )  ;
assign n24579 =  ( n31 ) & ( n24259 )  ;
assign n24580 =  ( n31 ) & ( n24261 )  ;
assign n24581 =  ( n31 ) & ( n24263 )  ;
assign n24582 =  ( n31 ) & ( n24265 )  ;
assign n24583 =  ( n31 ) & ( n24267 )  ;
assign n24584 =  ( n31 ) & ( n24269 )  ;
assign n24585 =  ( n31 ) & ( n24271 )  ;
assign n24586 =  ( n31 ) & ( n24273 )  ;
assign n24587 =  ( n31 ) & ( n24275 )  ;
assign n24588 =  ( n31 ) & ( n24277 )  ;
assign n24589 =  ( n31 ) & ( n24279 )  ;
assign n24590 =  ( n31 ) & ( n24281 )  ;
assign n24591 =  ( n31 ) & ( n24283 )  ;
assign n24592 =  ( n31 ) & ( n24285 )  ;
assign n24593 =  ( n31 ) & ( n24287 )  ;
assign n24594 =  ( n31 ) & ( n24289 )  ;
assign n24595 =  ( n32 ) & ( n24259 )  ;
assign n24596 =  ( n32 ) & ( n24261 )  ;
assign n24597 =  ( n32 ) & ( n24263 )  ;
assign n24598 =  ( n32 ) & ( n24265 )  ;
assign n24599 =  ( n32 ) & ( n24267 )  ;
assign n24600 =  ( n32 ) & ( n24269 )  ;
assign n24601 =  ( n32 ) & ( n24271 )  ;
assign n24602 =  ( n32 ) & ( n24273 )  ;
assign n24603 =  ( n32 ) & ( n24275 )  ;
assign n24604 =  ( n32 ) & ( n24277 )  ;
assign n24605 =  ( n32 ) & ( n24279 )  ;
assign n24606 =  ( n32 ) & ( n24281 )  ;
assign n24607 =  ( n32 ) & ( n24283 )  ;
assign n24608 =  ( n32 ) & ( n24285 )  ;
assign n24609 =  ( n32 ) & ( n24287 )  ;
assign n24610 =  ( n32 ) & ( n24289 )  ;
assign n24611 =  ( n33 ) & ( n24259 )  ;
assign n24612 =  ( n33 ) & ( n24261 )  ;
assign n24613 =  ( n33 ) & ( n24263 )  ;
assign n24614 =  ( n33 ) & ( n24265 )  ;
assign n24615 =  ( n33 ) & ( n24267 )  ;
assign n24616 =  ( n33 ) & ( n24269 )  ;
assign n24617 =  ( n33 ) & ( n24271 )  ;
assign n24618 =  ( n33 ) & ( n24273 )  ;
assign n24619 =  ( n33 ) & ( n24275 )  ;
assign n24620 =  ( n33 ) & ( n24277 )  ;
assign n24621 =  ( n33 ) & ( n24279 )  ;
assign n24622 =  ( n33 ) & ( n24281 )  ;
assign n24623 =  ( n33 ) & ( n24283 )  ;
assign n24624 =  ( n33 ) & ( n24285 )  ;
assign n24625 =  ( n33 ) & ( n24287 )  ;
assign n24626 =  ( n33 ) & ( n24289 )  ;
assign n24627 =  ( n34 ) & ( n24259 )  ;
assign n24628 =  ( n34 ) & ( n24261 )  ;
assign n24629 =  ( n34 ) & ( n24263 )  ;
assign n24630 =  ( n34 ) & ( n24265 )  ;
assign n24631 =  ( n34 ) & ( n24267 )  ;
assign n24632 =  ( n34 ) & ( n24269 )  ;
assign n24633 =  ( n34 ) & ( n24271 )  ;
assign n24634 =  ( n34 ) & ( n24273 )  ;
assign n24635 =  ( n34 ) & ( n24275 )  ;
assign n24636 =  ( n34 ) & ( n24277 )  ;
assign n24637 =  ( n34 ) & ( n24279 )  ;
assign n24638 =  ( n34 ) & ( n24281 )  ;
assign n24639 =  ( n34 ) & ( n24283 )  ;
assign n24640 =  ( n34 ) & ( n24285 )  ;
assign n24641 =  ( n34 ) & ( n24287 )  ;
assign n24642 =  ( n34 ) & ( n24289 )  ;
assign n24643 =  ( n35 ) & ( n24259 )  ;
assign n24644 =  ( n35 ) & ( n24261 )  ;
assign n24645 =  ( n35 ) & ( n24263 )  ;
assign n24646 =  ( n35 ) & ( n24265 )  ;
assign n24647 =  ( n35 ) & ( n24267 )  ;
assign n24648 =  ( n35 ) & ( n24269 )  ;
assign n24649 =  ( n35 ) & ( n24271 )  ;
assign n24650 =  ( n35 ) & ( n24273 )  ;
assign n24651 =  ( n35 ) & ( n24275 )  ;
assign n24652 =  ( n35 ) & ( n24277 )  ;
assign n24653 =  ( n35 ) & ( n24279 )  ;
assign n24654 =  ( n35 ) & ( n24281 )  ;
assign n24655 =  ( n35 ) & ( n24283 )  ;
assign n24656 =  ( n35 ) & ( n24285 )  ;
assign n24657 =  ( n35 ) & ( n24287 )  ;
assign n24658 =  ( n35 ) & ( n24289 )  ;
assign n24659 =  ( n36 ) & ( n24259 )  ;
assign n24660 =  ( n36 ) & ( n24261 )  ;
assign n24661 =  ( n36 ) & ( n24263 )  ;
assign n24662 =  ( n36 ) & ( n24265 )  ;
assign n24663 =  ( n36 ) & ( n24267 )  ;
assign n24664 =  ( n36 ) & ( n24269 )  ;
assign n24665 =  ( n36 ) & ( n24271 )  ;
assign n24666 =  ( n36 ) & ( n24273 )  ;
assign n24667 =  ( n36 ) & ( n24275 )  ;
assign n24668 =  ( n36 ) & ( n24277 )  ;
assign n24669 =  ( n36 ) & ( n24279 )  ;
assign n24670 =  ( n36 ) & ( n24281 )  ;
assign n24671 =  ( n36 ) & ( n24283 )  ;
assign n24672 =  ( n36 ) & ( n24285 )  ;
assign n24673 =  ( n36 ) & ( n24287 )  ;
assign n24674 =  ( n36 ) & ( n24289 )  ;
assign n24675 =  ( n37 ) & ( n24259 )  ;
assign n24676 =  ( n37 ) & ( n24261 )  ;
assign n24677 =  ( n37 ) & ( n24263 )  ;
assign n24678 =  ( n37 ) & ( n24265 )  ;
assign n24679 =  ( n37 ) & ( n24267 )  ;
assign n24680 =  ( n37 ) & ( n24269 )  ;
assign n24681 =  ( n37 ) & ( n24271 )  ;
assign n24682 =  ( n37 ) & ( n24273 )  ;
assign n24683 =  ( n37 ) & ( n24275 )  ;
assign n24684 =  ( n37 ) & ( n24277 )  ;
assign n24685 =  ( n37 ) & ( n24279 )  ;
assign n24686 =  ( n37 ) & ( n24281 )  ;
assign n24687 =  ( n37 ) & ( n24283 )  ;
assign n24688 =  ( n37 ) & ( n24285 )  ;
assign n24689 =  ( n37 ) & ( n24287 )  ;
assign n24690 =  ( n37 ) & ( n24289 )  ;
assign n24691 =  ( n38 ) & ( n24259 )  ;
assign n24692 =  ( n38 ) & ( n24261 )  ;
assign n24693 =  ( n38 ) & ( n24263 )  ;
assign n24694 =  ( n38 ) & ( n24265 )  ;
assign n24695 =  ( n38 ) & ( n24267 )  ;
assign n24696 =  ( n38 ) & ( n24269 )  ;
assign n24697 =  ( n38 ) & ( n24271 )  ;
assign n24698 =  ( n38 ) & ( n24273 )  ;
assign n24699 =  ( n38 ) & ( n24275 )  ;
assign n24700 =  ( n38 ) & ( n24277 )  ;
assign n24701 =  ( n38 ) & ( n24279 )  ;
assign n24702 =  ( n38 ) & ( n24281 )  ;
assign n24703 =  ( n38 ) & ( n24283 )  ;
assign n24704 =  ( n38 ) & ( n24285 )  ;
assign n24705 =  ( n38 ) & ( n24287 )  ;
assign n24706 =  ( n38 ) & ( n24289 )  ;
assign n24707 =  ( n39 ) & ( n24259 )  ;
assign n24708 =  ( n39 ) & ( n24261 )  ;
assign n24709 =  ( n39 ) & ( n24263 )  ;
assign n24710 =  ( n39 ) & ( n24265 )  ;
assign n24711 =  ( n39 ) & ( n24267 )  ;
assign n24712 =  ( n39 ) & ( n24269 )  ;
assign n24713 =  ( n39 ) & ( n24271 )  ;
assign n24714 =  ( n39 ) & ( n24273 )  ;
assign n24715 =  ( n39 ) & ( n24275 )  ;
assign n24716 =  ( n39 ) & ( n24277 )  ;
assign n24717 =  ( n39 ) & ( n24279 )  ;
assign n24718 =  ( n39 ) & ( n24281 )  ;
assign n24719 =  ( n39 ) & ( n24283 )  ;
assign n24720 =  ( n39 ) & ( n24285 )  ;
assign n24721 =  ( n39 ) & ( n24287 )  ;
assign n24722 =  ( n39 ) & ( n24289 )  ;
assign n24723 =  ( n40 ) & ( n24259 )  ;
assign n24724 =  ( n40 ) & ( n24261 )  ;
assign n24725 =  ( n40 ) & ( n24263 )  ;
assign n24726 =  ( n40 ) & ( n24265 )  ;
assign n24727 =  ( n40 ) & ( n24267 )  ;
assign n24728 =  ( n40 ) & ( n24269 )  ;
assign n24729 =  ( n40 ) & ( n24271 )  ;
assign n24730 =  ( n40 ) & ( n24273 )  ;
assign n24731 =  ( n40 ) & ( n24275 )  ;
assign n24732 =  ( n40 ) & ( n24277 )  ;
assign n24733 =  ( n40 ) & ( n24279 )  ;
assign n24734 =  ( n40 ) & ( n24281 )  ;
assign n24735 =  ( n40 ) & ( n24283 )  ;
assign n24736 =  ( n40 ) & ( n24285 )  ;
assign n24737 =  ( n40 ) & ( n24287 )  ;
assign n24738 =  ( n40 ) & ( n24289 )  ;
assign n24739 =  ( n41 ) & ( n24259 )  ;
assign n24740 =  ( n41 ) & ( n24261 )  ;
assign n24741 =  ( n41 ) & ( n24263 )  ;
assign n24742 =  ( n41 ) & ( n24265 )  ;
assign n24743 =  ( n41 ) & ( n24267 )  ;
assign n24744 =  ( n41 ) & ( n24269 )  ;
assign n24745 =  ( n41 ) & ( n24271 )  ;
assign n24746 =  ( n41 ) & ( n24273 )  ;
assign n24747 =  ( n41 ) & ( n24275 )  ;
assign n24748 =  ( n41 ) & ( n24277 )  ;
assign n24749 =  ( n41 ) & ( n24279 )  ;
assign n24750 =  ( n41 ) & ( n24281 )  ;
assign n24751 =  ( n41 ) & ( n24283 )  ;
assign n24752 =  ( n41 ) & ( n24285 )  ;
assign n24753 =  ( n41 ) & ( n24287 )  ;
assign n24754 =  ( n41 ) & ( n24289 )  ;
assign n24755 =  ( n42 ) & ( n24259 )  ;
assign n24756 =  ( n42 ) & ( n24261 )  ;
assign n24757 =  ( n42 ) & ( n24263 )  ;
assign n24758 =  ( n42 ) & ( n24265 )  ;
assign n24759 =  ( n42 ) & ( n24267 )  ;
assign n24760 =  ( n42 ) & ( n24269 )  ;
assign n24761 =  ( n42 ) & ( n24271 )  ;
assign n24762 =  ( n42 ) & ( n24273 )  ;
assign n24763 =  ( n42 ) & ( n24275 )  ;
assign n24764 =  ( n42 ) & ( n24277 )  ;
assign n24765 =  ( n42 ) & ( n24279 )  ;
assign n24766 =  ( n42 ) & ( n24281 )  ;
assign n24767 =  ( n42 ) & ( n24283 )  ;
assign n24768 =  ( n42 ) & ( n24285 )  ;
assign n24769 =  ( n42 ) & ( n24287 )  ;
assign n24770 =  ( n42 ) & ( n24289 )  ;
assign n24771 =  ( n43 ) & ( n24259 )  ;
assign n24772 =  ( n43 ) & ( n24261 )  ;
assign n24773 =  ( n43 ) & ( n24263 )  ;
assign n24774 =  ( n43 ) & ( n24265 )  ;
assign n24775 =  ( n43 ) & ( n24267 )  ;
assign n24776 =  ( n43 ) & ( n24269 )  ;
assign n24777 =  ( n43 ) & ( n24271 )  ;
assign n24778 =  ( n43 ) & ( n24273 )  ;
assign n24779 =  ( n43 ) & ( n24275 )  ;
assign n24780 =  ( n43 ) & ( n24277 )  ;
assign n24781 =  ( n43 ) & ( n24279 )  ;
assign n24782 =  ( n43 ) & ( n24281 )  ;
assign n24783 =  ( n43 ) & ( n24283 )  ;
assign n24784 =  ( n43 ) & ( n24285 )  ;
assign n24785 =  ( n43 ) & ( n24287 )  ;
assign n24786 =  ( n43 ) & ( n24289 )  ;
assign n24787 =  ( n24786 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n24788 =  ( n24785 ) ? ( VREG_0_1 ) : ( n24787 ) ;
assign n24789 =  ( n24784 ) ? ( VREG_0_2 ) : ( n24788 ) ;
assign n24790 =  ( n24783 ) ? ( VREG_0_3 ) : ( n24789 ) ;
assign n24791 =  ( n24782 ) ? ( VREG_0_4 ) : ( n24790 ) ;
assign n24792 =  ( n24781 ) ? ( VREG_0_5 ) : ( n24791 ) ;
assign n24793 =  ( n24780 ) ? ( VREG_0_6 ) : ( n24792 ) ;
assign n24794 =  ( n24779 ) ? ( VREG_0_7 ) : ( n24793 ) ;
assign n24795 =  ( n24778 ) ? ( VREG_0_8 ) : ( n24794 ) ;
assign n24796 =  ( n24777 ) ? ( VREG_0_9 ) : ( n24795 ) ;
assign n24797 =  ( n24776 ) ? ( VREG_0_10 ) : ( n24796 ) ;
assign n24798 =  ( n24775 ) ? ( VREG_0_11 ) : ( n24797 ) ;
assign n24799 =  ( n24774 ) ? ( VREG_0_12 ) : ( n24798 ) ;
assign n24800 =  ( n24773 ) ? ( VREG_0_13 ) : ( n24799 ) ;
assign n24801 =  ( n24772 ) ? ( VREG_0_14 ) : ( n24800 ) ;
assign n24802 =  ( n24771 ) ? ( VREG_0_15 ) : ( n24801 ) ;
assign n24803 =  ( n24770 ) ? ( VREG_1_0 ) : ( n24802 ) ;
assign n24804 =  ( n24769 ) ? ( VREG_1_1 ) : ( n24803 ) ;
assign n24805 =  ( n24768 ) ? ( VREG_1_2 ) : ( n24804 ) ;
assign n24806 =  ( n24767 ) ? ( VREG_1_3 ) : ( n24805 ) ;
assign n24807 =  ( n24766 ) ? ( VREG_1_4 ) : ( n24806 ) ;
assign n24808 =  ( n24765 ) ? ( VREG_1_5 ) : ( n24807 ) ;
assign n24809 =  ( n24764 ) ? ( VREG_1_6 ) : ( n24808 ) ;
assign n24810 =  ( n24763 ) ? ( VREG_1_7 ) : ( n24809 ) ;
assign n24811 =  ( n24762 ) ? ( VREG_1_8 ) : ( n24810 ) ;
assign n24812 =  ( n24761 ) ? ( VREG_1_9 ) : ( n24811 ) ;
assign n24813 =  ( n24760 ) ? ( VREG_1_10 ) : ( n24812 ) ;
assign n24814 =  ( n24759 ) ? ( VREG_1_11 ) : ( n24813 ) ;
assign n24815 =  ( n24758 ) ? ( VREG_1_12 ) : ( n24814 ) ;
assign n24816 =  ( n24757 ) ? ( VREG_1_13 ) : ( n24815 ) ;
assign n24817 =  ( n24756 ) ? ( VREG_1_14 ) : ( n24816 ) ;
assign n24818 =  ( n24755 ) ? ( VREG_1_15 ) : ( n24817 ) ;
assign n24819 =  ( n24754 ) ? ( VREG_2_0 ) : ( n24818 ) ;
assign n24820 =  ( n24753 ) ? ( VREG_2_1 ) : ( n24819 ) ;
assign n24821 =  ( n24752 ) ? ( VREG_2_2 ) : ( n24820 ) ;
assign n24822 =  ( n24751 ) ? ( VREG_2_3 ) : ( n24821 ) ;
assign n24823 =  ( n24750 ) ? ( VREG_2_4 ) : ( n24822 ) ;
assign n24824 =  ( n24749 ) ? ( VREG_2_5 ) : ( n24823 ) ;
assign n24825 =  ( n24748 ) ? ( VREG_2_6 ) : ( n24824 ) ;
assign n24826 =  ( n24747 ) ? ( VREG_2_7 ) : ( n24825 ) ;
assign n24827 =  ( n24746 ) ? ( VREG_2_8 ) : ( n24826 ) ;
assign n24828 =  ( n24745 ) ? ( VREG_2_9 ) : ( n24827 ) ;
assign n24829 =  ( n24744 ) ? ( VREG_2_10 ) : ( n24828 ) ;
assign n24830 =  ( n24743 ) ? ( VREG_2_11 ) : ( n24829 ) ;
assign n24831 =  ( n24742 ) ? ( VREG_2_12 ) : ( n24830 ) ;
assign n24832 =  ( n24741 ) ? ( VREG_2_13 ) : ( n24831 ) ;
assign n24833 =  ( n24740 ) ? ( VREG_2_14 ) : ( n24832 ) ;
assign n24834 =  ( n24739 ) ? ( VREG_2_15 ) : ( n24833 ) ;
assign n24835 =  ( n24738 ) ? ( VREG_3_0 ) : ( n24834 ) ;
assign n24836 =  ( n24737 ) ? ( VREG_3_1 ) : ( n24835 ) ;
assign n24837 =  ( n24736 ) ? ( VREG_3_2 ) : ( n24836 ) ;
assign n24838 =  ( n24735 ) ? ( VREG_3_3 ) : ( n24837 ) ;
assign n24839 =  ( n24734 ) ? ( VREG_3_4 ) : ( n24838 ) ;
assign n24840 =  ( n24733 ) ? ( VREG_3_5 ) : ( n24839 ) ;
assign n24841 =  ( n24732 ) ? ( VREG_3_6 ) : ( n24840 ) ;
assign n24842 =  ( n24731 ) ? ( VREG_3_7 ) : ( n24841 ) ;
assign n24843 =  ( n24730 ) ? ( VREG_3_8 ) : ( n24842 ) ;
assign n24844 =  ( n24729 ) ? ( VREG_3_9 ) : ( n24843 ) ;
assign n24845 =  ( n24728 ) ? ( VREG_3_10 ) : ( n24844 ) ;
assign n24846 =  ( n24727 ) ? ( VREG_3_11 ) : ( n24845 ) ;
assign n24847 =  ( n24726 ) ? ( VREG_3_12 ) : ( n24846 ) ;
assign n24848 =  ( n24725 ) ? ( VREG_3_13 ) : ( n24847 ) ;
assign n24849 =  ( n24724 ) ? ( VREG_3_14 ) : ( n24848 ) ;
assign n24850 =  ( n24723 ) ? ( VREG_3_15 ) : ( n24849 ) ;
assign n24851 =  ( n24722 ) ? ( VREG_4_0 ) : ( n24850 ) ;
assign n24852 =  ( n24721 ) ? ( VREG_4_1 ) : ( n24851 ) ;
assign n24853 =  ( n24720 ) ? ( VREG_4_2 ) : ( n24852 ) ;
assign n24854 =  ( n24719 ) ? ( VREG_4_3 ) : ( n24853 ) ;
assign n24855 =  ( n24718 ) ? ( VREG_4_4 ) : ( n24854 ) ;
assign n24856 =  ( n24717 ) ? ( VREG_4_5 ) : ( n24855 ) ;
assign n24857 =  ( n24716 ) ? ( VREG_4_6 ) : ( n24856 ) ;
assign n24858 =  ( n24715 ) ? ( VREG_4_7 ) : ( n24857 ) ;
assign n24859 =  ( n24714 ) ? ( VREG_4_8 ) : ( n24858 ) ;
assign n24860 =  ( n24713 ) ? ( VREG_4_9 ) : ( n24859 ) ;
assign n24861 =  ( n24712 ) ? ( VREG_4_10 ) : ( n24860 ) ;
assign n24862 =  ( n24711 ) ? ( VREG_4_11 ) : ( n24861 ) ;
assign n24863 =  ( n24710 ) ? ( VREG_4_12 ) : ( n24862 ) ;
assign n24864 =  ( n24709 ) ? ( VREG_4_13 ) : ( n24863 ) ;
assign n24865 =  ( n24708 ) ? ( VREG_4_14 ) : ( n24864 ) ;
assign n24866 =  ( n24707 ) ? ( VREG_4_15 ) : ( n24865 ) ;
assign n24867 =  ( n24706 ) ? ( VREG_5_0 ) : ( n24866 ) ;
assign n24868 =  ( n24705 ) ? ( VREG_5_1 ) : ( n24867 ) ;
assign n24869 =  ( n24704 ) ? ( VREG_5_2 ) : ( n24868 ) ;
assign n24870 =  ( n24703 ) ? ( VREG_5_3 ) : ( n24869 ) ;
assign n24871 =  ( n24702 ) ? ( VREG_5_4 ) : ( n24870 ) ;
assign n24872 =  ( n24701 ) ? ( VREG_5_5 ) : ( n24871 ) ;
assign n24873 =  ( n24700 ) ? ( VREG_5_6 ) : ( n24872 ) ;
assign n24874 =  ( n24699 ) ? ( VREG_5_7 ) : ( n24873 ) ;
assign n24875 =  ( n24698 ) ? ( VREG_5_8 ) : ( n24874 ) ;
assign n24876 =  ( n24697 ) ? ( VREG_5_9 ) : ( n24875 ) ;
assign n24877 =  ( n24696 ) ? ( VREG_5_10 ) : ( n24876 ) ;
assign n24878 =  ( n24695 ) ? ( VREG_5_11 ) : ( n24877 ) ;
assign n24879 =  ( n24694 ) ? ( VREG_5_12 ) : ( n24878 ) ;
assign n24880 =  ( n24693 ) ? ( VREG_5_13 ) : ( n24879 ) ;
assign n24881 =  ( n24692 ) ? ( VREG_5_14 ) : ( n24880 ) ;
assign n24882 =  ( n24691 ) ? ( VREG_5_15 ) : ( n24881 ) ;
assign n24883 =  ( n24690 ) ? ( VREG_6_0 ) : ( n24882 ) ;
assign n24884 =  ( n24689 ) ? ( VREG_6_1 ) : ( n24883 ) ;
assign n24885 =  ( n24688 ) ? ( VREG_6_2 ) : ( n24884 ) ;
assign n24886 =  ( n24687 ) ? ( VREG_6_3 ) : ( n24885 ) ;
assign n24887 =  ( n24686 ) ? ( VREG_6_4 ) : ( n24886 ) ;
assign n24888 =  ( n24685 ) ? ( VREG_6_5 ) : ( n24887 ) ;
assign n24889 =  ( n24684 ) ? ( VREG_6_6 ) : ( n24888 ) ;
assign n24890 =  ( n24683 ) ? ( VREG_6_7 ) : ( n24889 ) ;
assign n24891 =  ( n24682 ) ? ( VREG_6_8 ) : ( n24890 ) ;
assign n24892 =  ( n24681 ) ? ( VREG_6_9 ) : ( n24891 ) ;
assign n24893 =  ( n24680 ) ? ( VREG_6_10 ) : ( n24892 ) ;
assign n24894 =  ( n24679 ) ? ( VREG_6_11 ) : ( n24893 ) ;
assign n24895 =  ( n24678 ) ? ( VREG_6_12 ) : ( n24894 ) ;
assign n24896 =  ( n24677 ) ? ( VREG_6_13 ) : ( n24895 ) ;
assign n24897 =  ( n24676 ) ? ( VREG_6_14 ) : ( n24896 ) ;
assign n24898 =  ( n24675 ) ? ( VREG_6_15 ) : ( n24897 ) ;
assign n24899 =  ( n24674 ) ? ( VREG_7_0 ) : ( n24898 ) ;
assign n24900 =  ( n24673 ) ? ( VREG_7_1 ) : ( n24899 ) ;
assign n24901 =  ( n24672 ) ? ( VREG_7_2 ) : ( n24900 ) ;
assign n24902 =  ( n24671 ) ? ( VREG_7_3 ) : ( n24901 ) ;
assign n24903 =  ( n24670 ) ? ( VREG_7_4 ) : ( n24902 ) ;
assign n24904 =  ( n24669 ) ? ( VREG_7_5 ) : ( n24903 ) ;
assign n24905 =  ( n24668 ) ? ( VREG_7_6 ) : ( n24904 ) ;
assign n24906 =  ( n24667 ) ? ( VREG_7_7 ) : ( n24905 ) ;
assign n24907 =  ( n24666 ) ? ( VREG_7_8 ) : ( n24906 ) ;
assign n24908 =  ( n24665 ) ? ( VREG_7_9 ) : ( n24907 ) ;
assign n24909 =  ( n24664 ) ? ( VREG_7_10 ) : ( n24908 ) ;
assign n24910 =  ( n24663 ) ? ( VREG_7_11 ) : ( n24909 ) ;
assign n24911 =  ( n24662 ) ? ( VREG_7_12 ) : ( n24910 ) ;
assign n24912 =  ( n24661 ) ? ( VREG_7_13 ) : ( n24911 ) ;
assign n24913 =  ( n24660 ) ? ( VREG_7_14 ) : ( n24912 ) ;
assign n24914 =  ( n24659 ) ? ( VREG_7_15 ) : ( n24913 ) ;
assign n24915 =  ( n24658 ) ? ( VREG_8_0 ) : ( n24914 ) ;
assign n24916 =  ( n24657 ) ? ( VREG_8_1 ) : ( n24915 ) ;
assign n24917 =  ( n24656 ) ? ( VREG_8_2 ) : ( n24916 ) ;
assign n24918 =  ( n24655 ) ? ( VREG_8_3 ) : ( n24917 ) ;
assign n24919 =  ( n24654 ) ? ( VREG_8_4 ) : ( n24918 ) ;
assign n24920 =  ( n24653 ) ? ( VREG_8_5 ) : ( n24919 ) ;
assign n24921 =  ( n24652 ) ? ( VREG_8_6 ) : ( n24920 ) ;
assign n24922 =  ( n24651 ) ? ( VREG_8_7 ) : ( n24921 ) ;
assign n24923 =  ( n24650 ) ? ( VREG_8_8 ) : ( n24922 ) ;
assign n24924 =  ( n24649 ) ? ( VREG_8_9 ) : ( n24923 ) ;
assign n24925 =  ( n24648 ) ? ( VREG_8_10 ) : ( n24924 ) ;
assign n24926 =  ( n24647 ) ? ( VREG_8_11 ) : ( n24925 ) ;
assign n24927 =  ( n24646 ) ? ( VREG_8_12 ) : ( n24926 ) ;
assign n24928 =  ( n24645 ) ? ( VREG_8_13 ) : ( n24927 ) ;
assign n24929 =  ( n24644 ) ? ( VREG_8_14 ) : ( n24928 ) ;
assign n24930 =  ( n24643 ) ? ( VREG_8_15 ) : ( n24929 ) ;
assign n24931 =  ( n24642 ) ? ( VREG_9_0 ) : ( n24930 ) ;
assign n24932 =  ( n24641 ) ? ( VREG_9_1 ) : ( n24931 ) ;
assign n24933 =  ( n24640 ) ? ( VREG_9_2 ) : ( n24932 ) ;
assign n24934 =  ( n24639 ) ? ( VREG_9_3 ) : ( n24933 ) ;
assign n24935 =  ( n24638 ) ? ( VREG_9_4 ) : ( n24934 ) ;
assign n24936 =  ( n24637 ) ? ( VREG_9_5 ) : ( n24935 ) ;
assign n24937 =  ( n24636 ) ? ( VREG_9_6 ) : ( n24936 ) ;
assign n24938 =  ( n24635 ) ? ( VREG_9_7 ) : ( n24937 ) ;
assign n24939 =  ( n24634 ) ? ( VREG_9_8 ) : ( n24938 ) ;
assign n24940 =  ( n24633 ) ? ( VREG_9_9 ) : ( n24939 ) ;
assign n24941 =  ( n24632 ) ? ( VREG_9_10 ) : ( n24940 ) ;
assign n24942 =  ( n24631 ) ? ( VREG_9_11 ) : ( n24941 ) ;
assign n24943 =  ( n24630 ) ? ( VREG_9_12 ) : ( n24942 ) ;
assign n24944 =  ( n24629 ) ? ( VREG_9_13 ) : ( n24943 ) ;
assign n24945 =  ( n24628 ) ? ( VREG_9_14 ) : ( n24944 ) ;
assign n24946 =  ( n24627 ) ? ( VREG_9_15 ) : ( n24945 ) ;
assign n24947 =  ( n24626 ) ? ( VREG_10_0 ) : ( n24946 ) ;
assign n24948 =  ( n24625 ) ? ( VREG_10_1 ) : ( n24947 ) ;
assign n24949 =  ( n24624 ) ? ( VREG_10_2 ) : ( n24948 ) ;
assign n24950 =  ( n24623 ) ? ( VREG_10_3 ) : ( n24949 ) ;
assign n24951 =  ( n24622 ) ? ( VREG_10_4 ) : ( n24950 ) ;
assign n24952 =  ( n24621 ) ? ( VREG_10_5 ) : ( n24951 ) ;
assign n24953 =  ( n24620 ) ? ( VREG_10_6 ) : ( n24952 ) ;
assign n24954 =  ( n24619 ) ? ( VREG_10_7 ) : ( n24953 ) ;
assign n24955 =  ( n24618 ) ? ( VREG_10_8 ) : ( n24954 ) ;
assign n24956 =  ( n24617 ) ? ( VREG_10_9 ) : ( n24955 ) ;
assign n24957 =  ( n24616 ) ? ( VREG_10_10 ) : ( n24956 ) ;
assign n24958 =  ( n24615 ) ? ( VREG_10_11 ) : ( n24957 ) ;
assign n24959 =  ( n24614 ) ? ( VREG_10_12 ) : ( n24958 ) ;
assign n24960 =  ( n24613 ) ? ( VREG_10_13 ) : ( n24959 ) ;
assign n24961 =  ( n24612 ) ? ( VREG_10_14 ) : ( n24960 ) ;
assign n24962 =  ( n24611 ) ? ( VREG_10_15 ) : ( n24961 ) ;
assign n24963 =  ( n24610 ) ? ( VREG_11_0 ) : ( n24962 ) ;
assign n24964 =  ( n24609 ) ? ( VREG_11_1 ) : ( n24963 ) ;
assign n24965 =  ( n24608 ) ? ( VREG_11_2 ) : ( n24964 ) ;
assign n24966 =  ( n24607 ) ? ( VREG_11_3 ) : ( n24965 ) ;
assign n24967 =  ( n24606 ) ? ( VREG_11_4 ) : ( n24966 ) ;
assign n24968 =  ( n24605 ) ? ( VREG_11_5 ) : ( n24967 ) ;
assign n24969 =  ( n24604 ) ? ( VREG_11_6 ) : ( n24968 ) ;
assign n24970 =  ( n24603 ) ? ( VREG_11_7 ) : ( n24969 ) ;
assign n24971 =  ( n24602 ) ? ( VREG_11_8 ) : ( n24970 ) ;
assign n24972 =  ( n24601 ) ? ( VREG_11_9 ) : ( n24971 ) ;
assign n24973 =  ( n24600 ) ? ( VREG_11_10 ) : ( n24972 ) ;
assign n24974 =  ( n24599 ) ? ( VREG_11_11 ) : ( n24973 ) ;
assign n24975 =  ( n24598 ) ? ( VREG_11_12 ) : ( n24974 ) ;
assign n24976 =  ( n24597 ) ? ( VREG_11_13 ) : ( n24975 ) ;
assign n24977 =  ( n24596 ) ? ( VREG_11_14 ) : ( n24976 ) ;
assign n24978 =  ( n24595 ) ? ( VREG_11_15 ) : ( n24977 ) ;
assign n24979 =  ( n24594 ) ? ( VREG_12_0 ) : ( n24978 ) ;
assign n24980 =  ( n24593 ) ? ( VREG_12_1 ) : ( n24979 ) ;
assign n24981 =  ( n24592 ) ? ( VREG_12_2 ) : ( n24980 ) ;
assign n24982 =  ( n24591 ) ? ( VREG_12_3 ) : ( n24981 ) ;
assign n24983 =  ( n24590 ) ? ( VREG_12_4 ) : ( n24982 ) ;
assign n24984 =  ( n24589 ) ? ( VREG_12_5 ) : ( n24983 ) ;
assign n24985 =  ( n24588 ) ? ( VREG_12_6 ) : ( n24984 ) ;
assign n24986 =  ( n24587 ) ? ( VREG_12_7 ) : ( n24985 ) ;
assign n24987 =  ( n24586 ) ? ( VREG_12_8 ) : ( n24986 ) ;
assign n24988 =  ( n24585 ) ? ( VREG_12_9 ) : ( n24987 ) ;
assign n24989 =  ( n24584 ) ? ( VREG_12_10 ) : ( n24988 ) ;
assign n24990 =  ( n24583 ) ? ( VREG_12_11 ) : ( n24989 ) ;
assign n24991 =  ( n24582 ) ? ( VREG_12_12 ) : ( n24990 ) ;
assign n24992 =  ( n24581 ) ? ( VREG_12_13 ) : ( n24991 ) ;
assign n24993 =  ( n24580 ) ? ( VREG_12_14 ) : ( n24992 ) ;
assign n24994 =  ( n24579 ) ? ( VREG_12_15 ) : ( n24993 ) ;
assign n24995 =  ( n24578 ) ? ( VREG_13_0 ) : ( n24994 ) ;
assign n24996 =  ( n24577 ) ? ( VREG_13_1 ) : ( n24995 ) ;
assign n24997 =  ( n24576 ) ? ( VREG_13_2 ) : ( n24996 ) ;
assign n24998 =  ( n24575 ) ? ( VREG_13_3 ) : ( n24997 ) ;
assign n24999 =  ( n24574 ) ? ( VREG_13_4 ) : ( n24998 ) ;
assign n25000 =  ( n24573 ) ? ( VREG_13_5 ) : ( n24999 ) ;
assign n25001 =  ( n24572 ) ? ( VREG_13_6 ) : ( n25000 ) ;
assign n25002 =  ( n24571 ) ? ( VREG_13_7 ) : ( n25001 ) ;
assign n25003 =  ( n24570 ) ? ( VREG_13_8 ) : ( n25002 ) ;
assign n25004 =  ( n24569 ) ? ( VREG_13_9 ) : ( n25003 ) ;
assign n25005 =  ( n24568 ) ? ( VREG_13_10 ) : ( n25004 ) ;
assign n25006 =  ( n24567 ) ? ( VREG_13_11 ) : ( n25005 ) ;
assign n25007 =  ( n24566 ) ? ( VREG_13_12 ) : ( n25006 ) ;
assign n25008 =  ( n24565 ) ? ( VREG_13_13 ) : ( n25007 ) ;
assign n25009 =  ( n24564 ) ? ( VREG_13_14 ) : ( n25008 ) ;
assign n25010 =  ( n24563 ) ? ( VREG_13_15 ) : ( n25009 ) ;
assign n25011 =  ( n24562 ) ? ( VREG_14_0 ) : ( n25010 ) ;
assign n25012 =  ( n24561 ) ? ( VREG_14_1 ) : ( n25011 ) ;
assign n25013 =  ( n24560 ) ? ( VREG_14_2 ) : ( n25012 ) ;
assign n25014 =  ( n24559 ) ? ( VREG_14_3 ) : ( n25013 ) ;
assign n25015 =  ( n24558 ) ? ( VREG_14_4 ) : ( n25014 ) ;
assign n25016 =  ( n24557 ) ? ( VREG_14_5 ) : ( n25015 ) ;
assign n25017 =  ( n24556 ) ? ( VREG_14_6 ) : ( n25016 ) ;
assign n25018 =  ( n24555 ) ? ( VREG_14_7 ) : ( n25017 ) ;
assign n25019 =  ( n24554 ) ? ( VREG_14_8 ) : ( n25018 ) ;
assign n25020 =  ( n24553 ) ? ( VREG_14_9 ) : ( n25019 ) ;
assign n25021 =  ( n24552 ) ? ( VREG_14_10 ) : ( n25020 ) ;
assign n25022 =  ( n24551 ) ? ( VREG_14_11 ) : ( n25021 ) ;
assign n25023 =  ( n24550 ) ? ( VREG_14_12 ) : ( n25022 ) ;
assign n25024 =  ( n24549 ) ? ( VREG_14_13 ) : ( n25023 ) ;
assign n25025 =  ( n24548 ) ? ( VREG_14_14 ) : ( n25024 ) ;
assign n25026 =  ( n24547 ) ? ( VREG_14_15 ) : ( n25025 ) ;
assign n25027 =  ( n24546 ) ? ( VREG_15_0 ) : ( n25026 ) ;
assign n25028 =  ( n24545 ) ? ( VREG_15_1 ) : ( n25027 ) ;
assign n25029 =  ( n24544 ) ? ( VREG_15_2 ) : ( n25028 ) ;
assign n25030 =  ( n24543 ) ? ( VREG_15_3 ) : ( n25029 ) ;
assign n25031 =  ( n24542 ) ? ( VREG_15_4 ) : ( n25030 ) ;
assign n25032 =  ( n24541 ) ? ( VREG_15_5 ) : ( n25031 ) ;
assign n25033 =  ( n24540 ) ? ( VREG_15_6 ) : ( n25032 ) ;
assign n25034 =  ( n24539 ) ? ( VREG_15_7 ) : ( n25033 ) ;
assign n25035 =  ( n24538 ) ? ( VREG_15_8 ) : ( n25034 ) ;
assign n25036 =  ( n24537 ) ? ( VREG_15_9 ) : ( n25035 ) ;
assign n25037 =  ( n24536 ) ? ( VREG_15_10 ) : ( n25036 ) ;
assign n25038 =  ( n24535 ) ? ( VREG_15_11 ) : ( n25037 ) ;
assign n25039 =  ( n24534 ) ? ( VREG_15_12 ) : ( n25038 ) ;
assign n25040 =  ( n24533 ) ? ( VREG_15_13 ) : ( n25039 ) ;
assign n25041 =  ( n24532 ) ? ( VREG_15_14 ) : ( n25040 ) ;
assign n25042 =  ( n24531 ) ? ( VREG_15_15 ) : ( n25041 ) ;
assign n25043 =  ( n24530 ) ? ( VREG_16_0 ) : ( n25042 ) ;
assign n25044 =  ( n24529 ) ? ( VREG_16_1 ) : ( n25043 ) ;
assign n25045 =  ( n24528 ) ? ( VREG_16_2 ) : ( n25044 ) ;
assign n25046 =  ( n24527 ) ? ( VREG_16_3 ) : ( n25045 ) ;
assign n25047 =  ( n24526 ) ? ( VREG_16_4 ) : ( n25046 ) ;
assign n25048 =  ( n24525 ) ? ( VREG_16_5 ) : ( n25047 ) ;
assign n25049 =  ( n24524 ) ? ( VREG_16_6 ) : ( n25048 ) ;
assign n25050 =  ( n24523 ) ? ( VREG_16_7 ) : ( n25049 ) ;
assign n25051 =  ( n24522 ) ? ( VREG_16_8 ) : ( n25050 ) ;
assign n25052 =  ( n24521 ) ? ( VREG_16_9 ) : ( n25051 ) ;
assign n25053 =  ( n24520 ) ? ( VREG_16_10 ) : ( n25052 ) ;
assign n25054 =  ( n24519 ) ? ( VREG_16_11 ) : ( n25053 ) ;
assign n25055 =  ( n24518 ) ? ( VREG_16_12 ) : ( n25054 ) ;
assign n25056 =  ( n24517 ) ? ( VREG_16_13 ) : ( n25055 ) ;
assign n25057 =  ( n24516 ) ? ( VREG_16_14 ) : ( n25056 ) ;
assign n25058 =  ( n24515 ) ? ( VREG_16_15 ) : ( n25057 ) ;
assign n25059 =  ( n24514 ) ? ( VREG_17_0 ) : ( n25058 ) ;
assign n25060 =  ( n24513 ) ? ( VREG_17_1 ) : ( n25059 ) ;
assign n25061 =  ( n24512 ) ? ( VREG_17_2 ) : ( n25060 ) ;
assign n25062 =  ( n24511 ) ? ( VREG_17_3 ) : ( n25061 ) ;
assign n25063 =  ( n24510 ) ? ( VREG_17_4 ) : ( n25062 ) ;
assign n25064 =  ( n24509 ) ? ( VREG_17_5 ) : ( n25063 ) ;
assign n25065 =  ( n24508 ) ? ( VREG_17_6 ) : ( n25064 ) ;
assign n25066 =  ( n24507 ) ? ( VREG_17_7 ) : ( n25065 ) ;
assign n25067 =  ( n24506 ) ? ( VREG_17_8 ) : ( n25066 ) ;
assign n25068 =  ( n24505 ) ? ( VREG_17_9 ) : ( n25067 ) ;
assign n25069 =  ( n24504 ) ? ( VREG_17_10 ) : ( n25068 ) ;
assign n25070 =  ( n24503 ) ? ( VREG_17_11 ) : ( n25069 ) ;
assign n25071 =  ( n24502 ) ? ( VREG_17_12 ) : ( n25070 ) ;
assign n25072 =  ( n24501 ) ? ( VREG_17_13 ) : ( n25071 ) ;
assign n25073 =  ( n24500 ) ? ( VREG_17_14 ) : ( n25072 ) ;
assign n25074 =  ( n24499 ) ? ( VREG_17_15 ) : ( n25073 ) ;
assign n25075 =  ( n24498 ) ? ( VREG_18_0 ) : ( n25074 ) ;
assign n25076 =  ( n24497 ) ? ( VREG_18_1 ) : ( n25075 ) ;
assign n25077 =  ( n24496 ) ? ( VREG_18_2 ) : ( n25076 ) ;
assign n25078 =  ( n24495 ) ? ( VREG_18_3 ) : ( n25077 ) ;
assign n25079 =  ( n24494 ) ? ( VREG_18_4 ) : ( n25078 ) ;
assign n25080 =  ( n24493 ) ? ( VREG_18_5 ) : ( n25079 ) ;
assign n25081 =  ( n24492 ) ? ( VREG_18_6 ) : ( n25080 ) ;
assign n25082 =  ( n24491 ) ? ( VREG_18_7 ) : ( n25081 ) ;
assign n25083 =  ( n24490 ) ? ( VREG_18_8 ) : ( n25082 ) ;
assign n25084 =  ( n24489 ) ? ( VREG_18_9 ) : ( n25083 ) ;
assign n25085 =  ( n24488 ) ? ( VREG_18_10 ) : ( n25084 ) ;
assign n25086 =  ( n24487 ) ? ( VREG_18_11 ) : ( n25085 ) ;
assign n25087 =  ( n24486 ) ? ( VREG_18_12 ) : ( n25086 ) ;
assign n25088 =  ( n24485 ) ? ( VREG_18_13 ) : ( n25087 ) ;
assign n25089 =  ( n24484 ) ? ( VREG_18_14 ) : ( n25088 ) ;
assign n25090 =  ( n24483 ) ? ( VREG_18_15 ) : ( n25089 ) ;
assign n25091 =  ( n24482 ) ? ( VREG_19_0 ) : ( n25090 ) ;
assign n25092 =  ( n24481 ) ? ( VREG_19_1 ) : ( n25091 ) ;
assign n25093 =  ( n24480 ) ? ( VREG_19_2 ) : ( n25092 ) ;
assign n25094 =  ( n24479 ) ? ( VREG_19_3 ) : ( n25093 ) ;
assign n25095 =  ( n24478 ) ? ( VREG_19_4 ) : ( n25094 ) ;
assign n25096 =  ( n24477 ) ? ( VREG_19_5 ) : ( n25095 ) ;
assign n25097 =  ( n24476 ) ? ( VREG_19_6 ) : ( n25096 ) ;
assign n25098 =  ( n24475 ) ? ( VREG_19_7 ) : ( n25097 ) ;
assign n25099 =  ( n24474 ) ? ( VREG_19_8 ) : ( n25098 ) ;
assign n25100 =  ( n24473 ) ? ( VREG_19_9 ) : ( n25099 ) ;
assign n25101 =  ( n24472 ) ? ( VREG_19_10 ) : ( n25100 ) ;
assign n25102 =  ( n24471 ) ? ( VREG_19_11 ) : ( n25101 ) ;
assign n25103 =  ( n24470 ) ? ( VREG_19_12 ) : ( n25102 ) ;
assign n25104 =  ( n24469 ) ? ( VREG_19_13 ) : ( n25103 ) ;
assign n25105 =  ( n24468 ) ? ( VREG_19_14 ) : ( n25104 ) ;
assign n25106 =  ( n24467 ) ? ( VREG_19_15 ) : ( n25105 ) ;
assign n25107 =  ( n24466 ) ? ( VREG_20_0 ) : ( n25106 ) ;
assign n25108 =  ( n24465 ) ? ( VREG_20_1 ) : ( n25107 ) ;
assign n25109 =  ( n24464 ) ? ( VREG_20_2 ) : ( n25108 ) ;
assign n25110 =  ( n24463 ) ? ( VREG_20_3 ) : ( n25109 ) ;
assign n25111 =  ( n24462 ) ? ( VREG_20_4 ) : ( n25110 ) ;
assign n25112 =  ( n24461 ) ? ( VREG_20_5 ) : ( n25111 ) ;
assign n25113 =  ( n24460 ) ? ( VREG_20_6 ) : ( n25112 ) ;
assign n25114 =  ( n24459 ) ? ( VREG_20_7 ) : ( n25113 ) ;
assign n25115 =  ( n24458 ) ? ( VREG_20_8 ) : ( n25114 ) ;
assign n25116 =  ( n24457 ) ? ( VREG_20_9 ) : ( n25115 ) ;
assign n25117 =  ( n24456 ) ? ( VREG_20_10 ) : ( n25116 ) ;
assign n25118 =  ( n24455 ) ? ( VREG_20_11 ) : ( n25117 ) ;
assign n25119 =  ( n24454 ) ? ( VREG_20_12 ) : ( n25118 ) ;
assign n25120 =  ( n24453 ) ? ( VREG_20_13 ) : ( n25119 ) ;
assign n25121 =  ( n24452 ) ? ( VREG_20_14 ) : ( n25120 ) ;
assign n25122 =  ( n24451 ) ? ( VREG_20_15 ) : ( n25121 ) ;
assign n25123 =  ( n24450 ) ? ( VREG_21_0 ) : ( n25122 ) ;
assign n25124 =  ( n24449 ) ? ( VREG_21_1 ) : ( n25123 ) ;
assign n25125 =  ( n24448 ) ? ( VREG_21_2 ) : ( n25124 ) ;
assign n25126 =  ( n24447 ) ? ( VREG_21_3 ) : ( n25125 ) ;
assign n25127 =  ( n24446 ) ? ( VREG_21_4 ) : ( n25126 ) ;
assign n25128 =  ( n24445 ) ? ( VREG_21_5 ) : ( n25127 ) ;
assign n25129 =  ( n24444 ) ? ( VREG_21_6 ) : ( n25128 ) ;
assign n25130 =  ( n24443 ) ? ( VREG_21_7 ) : ( n25129 ) ;
assign n25131 =  ( n24442 ) ? ( VREG_21_8 ) : ( n25130 ) ;
assign n25132 =  ( n24441 ) ? ( VREG_21_9 ) : ( n25131 ) ;
assign n25133 =  ( n24440 ) ? ( VREG_21_10 ) : ( n25132 ) ;
assign n25134 =  ( n24439 ) ? ( VREG_21_11 ) : ( n25133 ) ;
assign n25135 =  ( n24438 ) ? ( VREG_21_12 ) : ( n25134 ) ;
assign n25136 =  ( n24437 ) ? ( VREG_21_13 ) : ( n25135 ) ;
assign n25137 =  ( n24436 ) ? ( VREG_21_14 ) : ( n25136 ) ;
assign n25138 =  ( n24435 ) ? ( VREG_21_15 ) : ( n25137 ) ;
assign n25139 =  ( n24434 ) ? ( VREG_22_0 ) : ( n25138 ) ;
assign n25140 =  ( n24433 ) ? ( VREG_22_1 ) : ( n25139 ) ;
assign n25141 =  ( n24432 ) ? ( VREG_22_2 ) : ( n25140 ) ;
assign n25142 =  ( n24431 ) ? ( VREG_22_3 ) : ( n25141 ) ;
assign n25143 =  ( n24430 ) ? ( VREG_22_4 ) : ( n25142 ) ;
assign n25144 =  ( n24429 ) ? ( VREG_22_5 ) : ( n25143 ) ;
assign n25145 =  ( n24428 ) ? ( VREG_22_6 ) : ( n25144 ) ;
assign n25146 =  ( n24427 ) ? ( VREG_22_7 ) : ( n25145 ) ;
assign n25147 =  ( n24426 ) ? ( VREG_22_8 ) : ( n25146 ) ;
assign n25148 =  ( n24425 ) ? ( VREG_22_9 ) : ( n25147 ) ;
assign n25149 =  ( n24424 ) ? ( VREG_22_10 ) : ( n25148 ) ;
assign n25150 =  ( n24423 ) ? ( VREG_22_11 ) : ( n25149 ) ;
assign n25151 =  ( n24422 ) ? ( VREG_22_12 ) : ( n25150 ) ;
assign n25152 =  ( n24421 ) ? ( VREG_22_13 ) : ( n25151 ) ;
assign n25153 =  ( n24420 ) ? ( VREG_22_14 ) : ( n25152 ) ;
assign n25154 =  ( n24419 ) ? ( VREG_22_15 ) : ( n25153 ) ;
assign n25155 =  ( n24418 ) ? ( VREG_23_0 ) : ( n25154 ) ;
assign n25156 =  ( n24417 ) ? ( VREG_23_1 ) : ( n25155 ) ;
assign n25157 =  ( n24416 ) ? ( VREG_23_2 ) : ( n25156 ) ;
assign n25158 =  ( n24415 ) ? ( VREG_23_3 ) : ( n25157 ) ;
assign n25159 =  ( n24414 ) ? ( VREG_23_4 ) : ( n25158 ) ;
assign n25160 =  ( n24413 ) ? ( VREG_23_5 ) : ( n25159 ) ;
assign n25161 =  ( n24412 ) ? ( VREG_23_6 ) : ( n25160 ) ;
assign n25162 =  ( n24411 ) ? ( VREG_23_7 ) : ( n25161 ) ;
assign n25163 =  ( n24410 ) ? ( VREG_23_8 ) : ( n25162 ) ;
assign n25164 =  ( n24409 ) ? ( VREG_23_9 ) : ( n25163 ) ;
assign n25165 =  ( n24408 ) ? ( VREG_23_10 ) : ( n25164 ) ;
assign n25166 =  ( n24407 ) ? ( VREG_23_11 ) : ( n25165 ) ;
assign n25167 =  ( n24406 ) ? ( VREG_23_12 ) : ( n25166 ) ;
assign n25168 =  ( n24405 ) ? ( VREG_23_13 ) : ( n25167 ) ;
assign n25169 =  ( n24404 ) ? ( VREG_23_14 ) : ( n25168 ) ;
assign n25170 =  ( n24403 ) ? ( VREG_23_15 ) : ( n25169 ) ;
assign n25171 =  ( n24402 ) ? ( VREG_24_0 ) : ( n25170 ) ;
assign n25172 =  ( n24401 ) ? ( VREG_24_1 ) : ( n25171 ) ;
assign n25173 =  ( n24400 ) ? ( VREG_24_2 ) : ( n25172 ) ;
assign n25174 =  ( n24399 ) ? ( VREG_24_3 ) : ( n25173 ) ;
assign n25175 =  ( n24398 ) ? ( VREG_24_4 ) : ( n25174 ) ;
assign n25176 =  ( n24397 ) ? ( VREG_24_5 ) : ( n25175 ) ;
assign n25177 =  ( n24396 ) ? ( VREG_24_6 ) : ( n25176 ) ;
assign n25178 =  ( n24395 ) ? ( VREG_24_7 ) : ( n25177 ) ;
assign n25179 =  ( n24394 ) ? ( VREG_24_8 ) : ( n25178 ) ;
assign n25180 =  ( n24393 ) ? ( VREG_24_9 ) : ( n25179 ) ;
assign n25181 =  ( n24392 ) ? ( VREG_24_10 ) : ( n25180 ) ;
assign n25182 =  ( n24391 ) ? ( VREG_24_11 ) : ( n25181 ) ;
assign n25183 =  ( n24390 ) ? ( VREG_24_12 ) : ( n25182 ) ;
assign n25184 =  ( n24389 ) ? ( VREG_24_13 ) : ( n25183 ) ;
assign n25185 =  ( n24388 ) ? ( VREG_24_14 ) : ( n25184 ) ;
assign n25186 =  ( n24387 ) ? ( VREG_24_15 ) : ( n25185 ) ;
assign n25187 =  ( n24386 ) ? ( VREG_25_0 ) : ( n25186 ) ;
assign n25188 =  ( n24385 ) ? ( VREG_25_1 ) : ( n25187 ) ;
assign n25189 =  ( n24384 ) ? ( VREG_25_2 ) : ( n25188 ) ;
assign n25190 =  ( n24383 ) ? ( VREG_25_3 ) : ( n25189 ) ;
assign n25191 =  ( n24382 ) ? ( VREG_25_4 ) : ( n25190 ) ;
assign n25192 =  ( n24381 ) ? ( VREG_25_5 ) : ( n25191 ) ;
assign n25193 =  ( n24380 ) ? ( VREG_25_6 ) : ( n25192 ) ;
assign n25194 =  ( n24379 ) ? ( VREG_25_7 ) : ( n25193 ) ;
assign n25195 =  ( n24378 ) ? ( VREG_25_8 ) : ( n25194 ) ;
assign n25196 =  ( n24377 ) ? ( VREG_25_9 ) : ( n25195 ) ;
assign n25197 =  ( n24376 ) ? ( VREG_25_10 ) : ( n25196 ) ;
assign n25198 =  ( n24375 ) ? ( VREG_25_11 ) : ( n25197 ) ;
assign n25199 =  ( n24374 ) ? ( VREG_25_12 ) : ( n25198 ) ;
assign n25200 =  ( n24373 ) ? ( VREG_25_13 ) : ( n25199 ) ;
assign n25201 =  ( n24372 ) ? ( VREG_25_14 ) : ( n25200 ) ;
assign n25202 =  ( n24371 ) ? ( VREG_25_15 ) : ( n25201 ) ;
assign n25203 =  ( n24370 ) ? ( VREG_26_0 ) : ( n25202 ) ;
assign n25204 =  ( n24369 ) ? ( VREG_26_1 ) : ( n25203 ) ;
assign n25205 =  ( n24368 ) ? ( VREG_26_2 ) : ( n25204 ) ;
assign n25206 =  ( n24367 ) ? ( VREG_26_3 ) : ( n25205 ) ;
assign n25207 =  ( n24366 ) ? ( VREG_26_4 ) : ( n25206 ) ;
assign n25208 =  ( n24365 ) ? ( VREG_26_5 ) : ( n25207 ) ;
assign n25209 =  ( n24364 ) ? ( VREG_26_6 ) : ( n25208 ) ;
assign n25210 =  ( n24363 ) ? ( VREG_26_7 ) : ( n25209 ) ;
assign n25211 =  ( n24362 ) ? ( VREG_26_8 ) : ( n25210 ) ;
assign n25212 =  ( n24361 ) ? ( VREG_26_9 ) : ( n25211 ) ;
assign n25213 =  ( n24360 ) ? ( VREG_26_10 ) : ( n25212 ) ;
assign n25214 =  ( n24359 ) ? ( VREG_26_11 ) : ( n25213 ) ;
assign n25215 =  ( n24358 ) ? ( VREG_26_12 ) : ( n25214 ) ;
assign n25216 =  ( n24357 ) ? ( VREG_26_13 ) : ( n25215 ) ;
assign n25217 =  ( n24356 ) ? ( VREG_26_14 ) : ( n25216 ) ;
assign n25218 =  ( n24355 ) ? ( VREG_26_15 ) : ( n25217 ) ;
assign n25219 =  ( n24354 ) ? ( VREG_27_0 ) : ( n25218 ) ;
assign n25220 =  ( n24353 ) ? ( VREG_27_1 ) : ( n25219 ) ;
assign n25221 =  ( n24352 ) ? ( VREG_27_2 ) : ( n25220 ) ;
assign n25222 =  ( n24351 ) ? ( VREG_27_3 ) : ( n25221 ) ;
assign n25223 =  ( n24350 ) ? ( VREG_27_4 ) : ( n25222 ) ;
assign n25224 =  ( n24349 ) ? ( VREG_27_5 ) : ( n25223 ) ;
assign n25225 =  ( n24348 ) ? ( VREG_27_6 ) : ( n25224 ) ;
assign n25226 =  ( n24347 ) ? ( VREG_27_7 ) : ( n25225 ) ;
assign n25227 =  ( n24346 ) ? ( VREG_27_8 ) : ( n25226 ) ;
assign n25228 =  ( n24345 ) ? ( VREG_27_9 ) : ( n25227 ) ;
assign n25229 =  ( n24344 ) ? ( VREG_27_10 ) : ( n25228 ) ;
assign n25230 =  ( n24343 ) ? ( VREG_27_11 ) : ( n25229 ) ;
assign n25231 =  ( n24342 ) ? ( VREG_27_12 ) : ( n25230 ) ;
assign n25232 =  ( n24341 ) ? ( VREG_27_13 ) : ( n25231 ) ;
assign n25233 =  ( n24340 ) ? ( VREG_27_14 ) : ( n25232 ) ;
assign n25234 =  ( n24339 ) ? ( VREG_27_15 ) : ( n25233 ) ;
assign n25235 =  ( n24338 ) ? ( VREG_28_0 ) : ( n25234 ) ;
assign n25236 =  ( n24337 ) ? ( VREG_28_1 ) : ( n25235 ) ;
assign n25237 =  ( n24336 ) ? ( VREG_28_2 ) : ( n25236 ) ;
assign n25238 =  ( n24335 ) ? ( VREG_28_3 ) : ( n25237 ) ;
assign n25239 =  ( n24334 ) ? ( VREG_28_4 ) : ( n25238 ) ;
assign n25240 =  ( n24333 ) ? ( VREG_28_5 ) : ( n25239 ) ;
assign n25241 =  ( n24332 ) ? ( VREG_28_6 ) : ( n25240 ) ;
assign n25242 =  ( n24331 ) ? ( VREG_28_7 ) : ( n25241 ) ;
assign n25243 =  ( n24330 ) ? ( VREG_28_8 ) : ( n25242 ) ;
assign n25244 =  ( n24329 ) ? ( VREG_28_9 ) : ( n25243 ) ;
assign n25245 =  ( n24328 ) ? ( VREG_28_10 ) : ( n25244 ) ;
assign n25246 =  ( n24327 ) ? ( VREG_28_11 ) : ( n25245 ) ;
assign n25247 =  ( n24326 ) ? ( VREG_28_12 ) : ( n25246 ) ;
assign n25248 =  ( n24325 ) ? ( VREG_28_13 ) : ( n25247 ) ;
assign n25249 =  ( n24324 ) ? ( VREG_28_14 ) : ( n25248 ) ;
assign n25250 =  ( n24323 ) ? ( VREG_28_15 ) : ( n25249 ) ;
assign n25251 =  ( n24322 ) ? ( VREG_29_0 ) : ( n25250 ) ;
assign n25252 =  ( n24321 ) ? ( VREG_29_1 ) : ( n25251 ) ;
assign n25253 =  ( n24320 ) ? ( VREG_29_2 ) : ( n25252 ) ;
assign n25254 =  ( n24319 ) ? ( VREG_29_3 ) : ( n25253 ) ;
assign n25255 =  ( n24318 ) ? ( VREG_29_4 ) : ( n25254 ) ;
assign n25256 =  ( n24317 ) ? ( VREG_29_5 ) : ( n25255 ) ;
assign n25257 =  ( n24316 ) ? ( VREG_29_6 ) : ( n25256 ) ;
assign n25258 =  ( n24315 ) ? ( VREG_29_7 ) : ( n25257 ) ;
assign n25259 =  ( n24314 ) ? ( VREG_29_8 ) : ( n25258 ) ;
assign n25260 =  ( n24313 ) ? ( VREG_29_9 ) : ( n25259 ) ;
assign n25261 =  ( n24312 ) ? ( VREG_29_10 ) : ( n25260 ) ;
assign n25262 =  ( n24311 ) ? ( VREG_29_11 ) : ( n25261 ) ;
assign n25263 =  ( n24310 ) ? ( VREG_29_12 ) : ( n25262 ) ;
assign n25264 =  ( n24309 ) ? ( VREG_29_13 ) : ( n25263 ) ;
assign n25265 =  ( n24308 ) ? ( VREG_29_14 ) : ( n25264 ) ;
assign n25266 =  ( n24307 ) ? ( VREG_29_15 ) : ( n25265 ) ;
assign n25267 =  ( n24306 ) ? ( VREG_30_0 ) : ( n25266 ) ;
assign n25268 =  ( n24305 ) ? ( VREG_30_1 ) : ( n25267 ) ;
assign n25269 =  ( n24304 ) ? ( VREG_30_2 ) : ( n25268 ) ;
assign n25270 =  ( n24303 ) ? ( VREG_30_3 ) : ( n25269 ) ;
assign n25271 =  ( n24302 ) ? ( VREG_30_4 ) : ( n25270 ) ;
assign n25272 =  ( n24301 ) ? ( VREG_30_5 ) : ( n25271 ) ;
assign n25273 =  ( n24300 ) ? ( VREG_30_6 ) : ( n25272 ) ;
assign n25274 =  ( n24299 ) ? ( VREG_30_7 ) : ( n25273 ) ;
assign n25275 =  ( n24298 ) ? ( VREG_30_8 ) : ( n25274 ) ;
assign n25276 =  ( n24297 ) ? ( VREG_30_9 ) : ( n25275 ) ;
assign n25277 =  ( n24296 ) ? ( VREG_30_10 ) : ( n25276 ) ;
assign n25278 =  ( n24295 ) ? ( VREG_30_11 ) : ( n25277 ) ;
assign n25279 =  ( n24294 ) ? ( VREG_30_12 ) : ( n25278 ) ;
assign n25280 =  ( n24293 ) ? ( VREG_30_13 ) : ( n25279 ) ;
assign n25281 =  ( n24292 ) ? ( VREG_30_14 ) : ( n25280 ) ;
assign n25282 =  ( n24291 ) ? ( VREG_30_15 ) : ( n25281 ) ;
assign n25283 =  ( n24290 ) ? ( VREG_31_0 ) : ( n25282 ) ;
assign n25284 =  ( n24288 ) ? ( VREG_31_1 ) : ( n25283 ) ;
assign n25285 =  ( n24286 ) ? ( VREG_31_2 ) : ( n25284 ) ;
assign n25286 =  ( n24284 ) ? ( VREG_31_3 ) : ( n25285 ) ;
assign n25287 =  ( n24282 ) ? ( VREG_31_4 ) : ( n25286 ) ;
assign n25288 =  ( n24280 ) ? ( VREG_31_5 ) : ( n25287 ) ;
assign n25289 =  ( n24278 ) ? ( VREG_31_6 ) : ( n25288 ) ;
assign n25290 =  ( n24276 ) ? ( VREG_31_7 ) : ( n25289 ) ;
assign n25291 =  ( n24274 ) ? ( VREG_31_8 ) : ( n25290 ) ;
assign n25292 =  ( n24272 ) ? ( VREG_31_9 ) : ( n25291 ) ;
assign n25293 =  ( n24270 ) ? ( VREG_31_10 ) : ( n25292 ) ;
assign n25294 =  ( n24268 ) ? ( VREG_31_11 ) : ( n25293 ) ;
assign n25295 =  ( n24266 ) ? ( VREG_31_12 ) : ( n25294 ) ;
assign n25296 =  ( n24264 ) ? ( VREG_31_13 ) : ( n25295 ) ;
assign n25297 =  ( n24262 ) ? ( VREG_31_14 ) : ( n25296 ) ;
assign n25298 =  ( n24260 ) ? ( VREG_31_15 ) : ( n25297 ) ;
assign n25299 =  ( n25298 ) + ( n140 )  ;
assign n25300 =  ( n25298 ) - ( n140 )  ;
assign n25301 =  ( n25298 ) & ( n140 )  ;
assign n25302 =  ( n25298 ) | ( n140 )  ;
assign n25303 =  ( ( n25298 ) * ( n140 ))  ;
assign n25304 =  ( n148 ) ? ( n25303 ) : ( VREG_0_5 ) ;
assign n25305 =  ( n146 ) ? ( n25302 ) : ( n25304 ) ;
assign n25306 =  ( n144 ) ? ( n25301 ) : ( n25305 ) ;
assign n25307 =  ( n142 ) ? ( n25300 ) : ( n25306 ) ;
assign n25308 =  ( n10 ) ? ( n25299 ) : ( n25307 ) ;
assign n25309 =  ( n77 ) & ( n24259 )  ;
assign n25310 =  ( n77 ) & ( n24261 )  ;
assign n25311 =  ( n77 ) & ( n24263 )  ;
assign n25312 =  ( n77 ) & ( n24265 )  ;
assign n25313 =  ( n77 ) & ( n24267 )  ;
assign n25314 =  ( n77 ) & ( n24269 )  ;
assign n25315 =  ( n77 ) & ( n24271 )  ;
assign n25316 =  ( n77 ) & ( n24273 )  ;
assign n25317 =  ( n77 ) & ( n24275 )  ;
assign n25318 =  ( n77 ) & ( n24277 )  ;
assign n25319 =  ( n77 ) & ( n24279 )  ;
assign n25320 =  ( n77 ) & ( n24281 )  ;
assign n25321 =  ( n77 ) & ( n24283 )  ;
assign n25322 =  ( n77 ) & ( n24285 )  ;
assign n25323 =  ( n77 ) & ( n24287 )  ;
assign n25324 =  ( n77 ) & ( n24289 )  ;
assign n25325 =  ( n78 ) & ( n24259 )  ;
assign n25326 =  ( n78 ) & ( n24261 )  ;
assign n25327 =  ( n78 ) & ( n24263 )  ;
assign n25328 =  ( n78 ) & ( n24265 )  ;
assign n25329 =  ( n78 ) & ( n24267 )  ;
assign n25330 =  ( n78 ) & ( n24269 )  ;
assign n25331 =  ( n78 ) & ( n24271 )  ;
assign n25332 =  ( n78 ) & ( n24273 )  ;
assign n25333 =  ( n78 ) & ( n24275 )  ;
assign n25334 =  ( n78 ) & ( n24277 )  ;
assign n25335 =  ( n78 ) & ( n24279 )  ;
assign n25336 =  ( n78 ) & ( n24281 )  ;
assign n25337 =  ( n78 ) & ( n24283 )  ;
assign n25338 =  ( n78 ) & ( n24285 )  ;
assign n25339 =  ( n78 ) & ( n24287 )  ;
assign n25340 =  ( n78 ) & ( n24289 )  ;
assign n25341 =  ( n79 ) & ( n24259 )  ;
assign n25342 =  ( n79 ) & ( n24261 )  ;
assign n25343 =  ( n79 ) & ( n24263 )  ;
assign n25344 =  ( n79 ) & ( n24265 )  ;
assign n25345 =  ( n79 ) & ( n24267 )  ;
assign n25346 =  ( n79 ) & ( n24269 )  ;
assign n25347 =  ( n79 ) & ( n24271 )  ;
assign n25348 =  ( n79 ) & ( n24273 )  ;
assign n25349 =  ( n79 ) & ( n24275 )  ;
assign n25350 =  ( n79 ) & ( n24277 )  ;
assign n25351 =  ( n79 ) & ( n24279 )  ;
assign n25352 =  ( n79 ) & ( n24281 )  ;
assign n25353 =  ( n79 ) & ( n24283 )  ;
assign n25354 =  ( n79 ) & ( n24285 )  ;
assign n25355 =  ( n79 ) & ( n24287 )  ;
assign n25356 =  ( n79 ) & ( n24289 )  ;
assign n25357 =  ( n80 ) & ( n24259 )  ;
assign n25358 =  ( n80 ) & ( n24261 )  ;
assign n25359 =  ( n80 ) & ( n24263 )  ;
assign n25360 =  ( n80 ) & ( n24265 )  ;
assign n25361 =  ( n80 ) & ( n24267 )  ;
assign n25362 =  ( n80 ) & ( n24269 )  ;
assign n25363 =  ( n80 ) & ( n24271 )  ;
assign n25364 =  ( n80 ) & ( n24273 )  ;
assign n25365 =  ( n80 ) & ( n24275 )  ;
assign n25366 =  ( n80 ) & ( n24277 )  ;
assign n25367 =  ( n80 ) & ( n24279 )  ;
assign n25368 =  ( n80 ) & ( n24281 )  ;
assign n25369 =  ( n80 ) & ( n24283 )  ;
assign n25370 =  ( n80 ) & ( n24285 )  ;
assign n25371 =  ( n80 ) & ( n24287 )  ;
assign n25372 =  ( n80 ) & ( n24289 )  ;
assign n25373 =  ( n81 ) & ( n24259 )  ;
assign n25374 =  ( n81 ) & ( n24261 )  ;
assign n25375 =  ( n81 ) & ( n24263 )  ;
assign n25376 =  ( n81 ) & ( n24265 )  ;
assign n25377 =  ( n81 ) & ( n24267 )  ;
assign n25378 =  ( n81 ) & ( n24269 )  ;
assign n25379 =  ( n81 ) & ( n24271 )  ;
assign n25380 =  ( n81 ) & ( n24273 )  ;
assign n25381 =  ( n81 ) & ( n24275 )  ;
assign n25382 =  ( n81 ) & ( n24277 )  ;
assign n25383 =  ( n81 ) & ( n24279 )  ;
assign n25384 =  ( n81 ) & ( n24281 )  ;
assign n25385 =  ( n81 ) & ( n24283 )  ;
assign n25386 =  ( n81 ) & ( n24285 )  ;
assign n25387 =  ( n81 ) & ( n24287 )  ;
assign n25388 =  ( n81 ) & ( n24289 )  ;
assign n25389 =  ( n82 ) & ( n24259 )  ;
assign n25390 =  ( n82 ) & ( n24261 )  ;
assign n25391 =  ( n82 ) & ( n24263 )  ;
assign n25392 =  ( n82 ) & ( n24265 )  ;
assign n25393 =  ( n82 ) & ( n24267 )  ;
assign n25394 =  ( n82 ) & ( n24269 )  ;
assign n25395 =  ( n82 ) & ( n24271 )  ;
assign n25396 =  ( n82 ) & ( n24273 )  ;
assign n25397 =  ( n82 ) & ( n24275 )  ;
assign n25398 =  ( n82 ) & ( n24277 )  ;
assign n25399 =  ( n82 ) & ( n24279 )  ;
assign n25400 =  ( n82 ) & ( n24281 )  ;
assign n25401 =  ( n82 ) & ( n24283 )  ;
assign n25402 =  ( n82 ) & ( n24285 )  ;
assign n25403 =  ( n82 ) & ( n24287 )  ;
assign n25404 =  ( n82 ) & ( n24289 )  ;
assign n25405 =  ( n83 ) & ( n24259 )  ;
assign n25406 =  ( n83 ) & ( n24261 )  ;
assign n25407 =  ( n83 ) & ( n24263 )  ;
assign n25408 =  ( n83 ) & ( n24265 )  ;
assign n25409 =  ( n83 ) & ( n24267 )  ;
assign n25410 =  ( n83 ) & ( n24269 )  ;
assign n25411 =  ( n83 ) & ( n24271 )  ;
assign n25412 =  ( n83 ) & ( n24273 )  ;
assign n25413 =  ( n83 ) & ( n24275 )  ;
assign n25414 =  ( n83 ) & ( n24277 )  ;
assign n25415 =  ( n83 ) & ( n24279 )  ;
assign n25416 =  ( n83 ) & ( n24281 )  ;
assign n25417 =  ( n83 ) & ( n24283 )  ;
assign n25418 =  ( n83 ) & ( n24285 )  ;
assign n25419 =  ( n83 ) & ( n24287 )  ;
assign n25420 =  ( n83 ) & ( n24289 )  ;
assign n25421 =  ( n84 ) & ( n24259 )  ;
assign n25422 =  ( n84 ) & ( n24261 )  ;
assign n25423 =  ( n84 ) & ( n24263 )  ;
assign n25424 =  ( n84 ) & ( n24265 )  ;
assign n25425 =  ( n84 ) & ( n24267 )  ;
assign n25426 =  ( n84 ) & ( n24269 )  ;
assign n25427 =  ( n84 ) & ( n24271 )  ;
assign n25428 =  ( n84 ) & ( n24273 )  ;
assign n25429 =  ( n84 ) & ( n24275 )  ;
assign n25430 =  ( n84 ) & ( n24277 )  ;
assign n25431 =  ( n84 ) & ( n24279 )  ;
assign n25432 =  ( n84 ) & ( n24281 )  ;
assign n25433 =  ( n84 ) & ( n24283 )  ;
assign n25434 =  ( n84 ) & ( n24285 )  ;
assign n25435 =  ( n84 ) & ( n24287 )  ;
assign n25436 =  ( n84 ) & ( n24289 )  ;
assign n25437 =  ( n85 ) & ( n24259 )  ;
assign n25438 =  ( n85 ) & ( n24261 )  ;
assign n25439 =  ( n85 ) & ( n24263 )  ;
assign n25440 =  ( n85 ) & ( n24265 )  ;
assign n25441 =  ( n85 ) & ( n24267 )  ;
assign n25442 =  ( n85 ) & ( n24269 )  ;
assign n25443 =  ( n85 ) & ( n24271 )  ;
assign n25444 =  ( n85 ) & ( n24273 )  ;
assign n25445 =  ( n85 ) & ( n24275 )  ;
assign n25446 =  ( n85 ) & ( n24277 )  ;
assign n25447 =  ( n85 ) & ( n24279 )  ;
assign n25448 =  ( n85 ) & ( n24281 )  ;
assign n25449 =  ( n85 ) & ( n24283 )  ;
assign n25450 =  ( n85 ) & ( n24285 )  ;
assign n25451 =  ( n85 ) & ( n24287 )  ;
assign n25452 =  ( n85 ) & ( n24289 )  ;
assign n25453 =  ( n86 ) & ( n24259 )  ;
assign n25454 =  ( n86 ) & ( n24261 )  ;
assign n25455 =  ( n86 ) & ( n24263 )  ;
assign n25456 =  ( n86 ) & ( n24265 )  ;
assign n25457 =  ( n86 ) & ( n24267 )  ;
assign n25458 =  ( n86 ) & ( n24269 )  ;
assign n25459 =  ( n86 ) & ( n24271 )  ;
assign n25460 =  ( n86 ) & ( n24273 )  ;
assign n25461 =  ( n86 ) & ( n24275 )  ;
assign n25462 =  ( n86 ) & ( n24277 )  ;
assign n25463 =  ( n86 ) & ( n24279 )  ;
assign n25464 =  ( n86 ) & ( n24281 )  ;
assign n25465 =  ( n86 ) & ( n24283 )  ;
assign n25466 =  ( n86 ) & ( n24285 )  ;
assign n25467 =  ( n86 ) & ( n24287 )  ;
assign n25468 =  ( n86 ) & ( n24289 )  ;
assign n25469 =  ( n87 ) & ( n24259 )  ;
assign n25470 =  ( n87 ) & ( n24261 )  ;
assign n25471 =  ( n87 ) & ( n24263 )  ;
assign n25472 =  ( n87 ) & ( n24265 )  ;
assign n25473 =  ( n87 ) & ( n24267 )  ;
assign n25474 =  ( n87 ) & ( n24269 )  ;
assign n25475 =  ( n87 ) & ( n24271 )  ;
assign n25476 =  ( n87 ) & ( n24273 )  ;
assign n25477 =  ( n87 ) & ( n24275 )  ;
assign n25478 =  ( n87 ) & ( n24277 )  ;
assign n25479 =  ( n87 ) & ( n24279 )  ;
assign n25480 =  ( n87 ) & ( n24281 )  ;
assign n25481 =  ( n87 ) & ( n24283 )  ;
assign n25482 =  ( n87 ) & ( n24285 )  ;
assign n25483 =  ( n87 ) & ( n24287 )  ;
assign n25484 =  ( n87 ) & ( n24289 )  ;
assign n25485 =  ( n88 ) & ( n24259 )  ;
assign n25486 =  ( n88 ) & ( n24261 )  ;
assign n25487 =  ( n88 ) & ( n24263 )  ;
assign n25488 =  ( n88 ) & ( n24265 )  ;
assign n25489 =  ( n88 ) & ( n24267 )  ;
assign n25490 =  ( n88 ) & ( n24269 )  ;
assign n25491 =  ( n88 ) & ( n24271 )  ;
assign n25492 =  ( n88 ) & ( n24273 )  ;
assign n25493 =  ( n88 ) & ( n24275 )  ;
assign n25494 =  ( n88 ) & ( n24277 )  ;
assign n25495 =  ( n88 ) & ( n24279 )  ;
assign n25496 =  ( n88 ) & ( n24281 )  ;
assign n25497 =  ( n88 ) & ( n24283 )  ;
assign n25498 =  ( n88 ) & ( n24285 )  ;
assign n25499 =  ( n88 ) & ( n24287 )  ;
assign n25500 =  ( n88 ) & ( n24289 )  ;
assign n25501 =  ( n89 ) & ( n24259 )  ;
assign n25502 =  ( n89 ) & ( n24261 )  ;
assign n25503 =  ( n89 ) & ( n24263 )  ;
assign n25504 =  ( n89 ) & ( n24265 )  ;
assign n25505 =  ( n89 ) & ( n24267 )  ;
assign n25506 =  ( n89 ) & ( n24269 )  ;
assign n25507 =  ( n89 ) & ( n24271 )  ;
assign n25508 =  ( n89 ) & ( n24273 )  ;
assign n25509 =  ( n89 ) & ( n24275 )  ;
assign n25510 =  ( n89 ) & ( n24277 )  ;
assign n25511 =  ( n89 ) & ( n24279 )  ;
assign n25512 =  ( n89 ) & ( n24281 )  ;
assign n25513 =  ( n89 ) & ( n24283 )  ;
assign n25514 =  ( n89 ) & ( n24285 )  ;
assign n25515 =  ( n89 ) & ( n24287 )  ;
assign n25516 =  ( n89 ) & ( n24289 )  ;
assign n25517 =  ( n90 ) & ( n24259 )  ;
assign n25518 =  ( n90 ) & ( n24261 )  ;
assign n25519 =  ( n90 ) & ( n24263 )  ;
assign n25520 =  ( n90 ) & ( n24265 )  ;
assign n25521 =  ( n90 ) & ( n24267 )  ;
assign n25522 =  ( n90 ) & ( n24269 )  ;
assign n25523 =  ( n90 ) & ( n24271 )  ;
assign n25524 =  ( n90 ) & ( n24273 )  ;
assign n25525 =  ( n90 ) & ( n24275 )  ;
assign n25526 =  ( n90 ) & ( n24277 )  ;
assign n25527 =  ( n90 ) & ( n24279 )  ;
assign n25528 =  ( n90 ) & ( n24281 )  ;
assign n25529 =  ( n90 ) & ( n24283 )  ;
assign n25530 =  ( n90 ) & ( n24285 )  ;
assign n25531 =  ( n90 ) & ( n24287 )  ;
assign n25532 =  ( n90 ) & ( n24289 )  ;
assign n25533 =  ( n91 ) & ( n24259 )  ;
assign n25534 =  ( n91 ) & ( n24261 )  ;
assign n25535 =  ( n91 ) & ( n24263 )  ;
assign n25536 =  ( n91 ) & ( n24265 )  ;
assign n25537 =  ( n91 ) & ( n24267 )  ;
assign n25538 =  ( n91 ) & ( n24269 )  ;
assign n25539 =  ( n91 ) & ( n24271 )  ;
assign n25540 =  ( n91 ) & ( n24273 )  ;
assign n25541 =  ( n91 ) & ( n24275 )  ;
assign n25542 =  ( n91 ) & ( n24277 )  ;
assign n25543 =  ( n91 ) & ( n24279 )  ;
assign n25544 =  ( n91 ) & ( n24281 )  ;
assign n25545 =  ( n91 ) & ( n24283 )  ;
assign n25546 =  ( n91 ) & ( n24285 )  ;
assign n25547 =  ( n91 ) & ( n24287 )  ;
assign n25548 =  ( n91 ) & ( n24289 )  ;
assign n25549 =  ( n92 ) & ( n24259 )  ;
assign n25550 =  ( n92 ) & ( n24261 )  ;
assign n25551 =  ( n92 ) & ( n24263 )  ;
assign n25552 =  ( n92 ) & ( n24265 )  ;
assign n25553 =  ( n92 ) & ( n24267 )  ;
assign n25554 =  ( n92 ) & ( n24269 )  ;
assign n25555 =  ( n92 ) & ( n24271 )  ;
assign n25556 =  ( n92 ) & ( n24273 )  ;
assign n25557 =  ( n92 ) & ( n24275 )  ;
assign n25558 =  ( n92 ) & ( n24277 )  ;
assign n25559 =  ( n92 ) & ( n24279 )  ;
assign n25560 =  ( n92 ) & ( n24281 )  ;
assign n25561 =  ( n92 ) & ( n24283 )  ;
assign n25562 =  ( n92 ) & ( n24285 )  ;
assign n25563 =  ( n92 ) & ( n24287 )  ;
assign n25564 =  ( n92 ) & ( n24289 )  ;
assign n25565 =  ( n93 ) & ( n24259 )  ;
assign n25566 =  ( n93 ) & ( n24261 )  ;
assign n25567 =  ( n93 ) & ( n24263 )  ;
assign n25568 =  ( n93 ) & ( n24265 )  ;
assign n25569 =  ( n93 ) & ( n24267 )  ;
assign n25570 =  ( n93 ) & ( n24269 )  ;
assign n25571 =  ( n93 ) & ( n24271 )  ;
assign n25572 =  ( n93 ) & ( n24273 )  ;
assign n25573 =  ( n93 ) & ( n24275 )  ;
assign n25574 =  ( n93 ) & ( n24277 )  ;
assign n25575 =  ( n93 ) & ( n24279 )  ;
assign n25576 =  ( n93 ) & ( n24281 )  ;
assign n25577 =  ( n93 ) & ( n24283 )  ;
assign n25578 =  ( n93 ) & ( n24285 )  ;
assign n25579 =  ( n93 ) & ( n24287 )  ;
assign n25580 =  ( n93 ) & ( n24289 )  ;
assign n25581 =  ( n94 ) & ( n24259 )  ;
assign n25582 =  ( n94 ) & ( n24261 )  ;
assign n25583 =  ( n94 ) & ( n24263 )  ;
assign n25584 =  ( n94 ) & ( n24265 )  ;
assign n25585 =  ( n94 ) & ( n24267 )  ;
assign n25586 =  ( n94 ) & ( n24269 )  ;
assign n25587 =  ( n94 ) & ( n24271 )  ;
assign n25588 =  ( n94 ) & ( n24273 )  ;
assign n25589 =  ( n94 ) & ( n24275 )  ;
assign n25590 =  ( n94 ) & ( n24277 )  ;
assign n25591 =  ( n94 ) & ( n24279 )  ;
assign n25592 =  ( n94 ) & ( n24281 )  ;
assign n25593 =  ( n94 ) & ( n24283 )  ;
assign n25594 =  ( n94 ) & ( n24285 )  ;
assign n25595 =  ( n94 ) & ( n24287 )  ;
assign n25596 =  ( n94 ) & ( n24289 )  ;
assign n25597 =  ( n95 ) & ( n24259 )  ;
assign n25598 =  ( n95 ) & ( n24261 )  ;
assign n25599 =  ( n95 ) & ( n24263 )  ;
assign n25600 =  ( n95 ) & ( n24265 )  ;
assign n25601 =  ( n95 ) & ( n24267 )  ;
assign n25602 =  ( n95 ) & ( n24269 )  ;
assign n25603 =  ( n95 ) & ( n24271 )  ;
assign n25604 =  ( n95 ) & ( n24273 )  ;
assign n25605 =  ( n95 ) & ( n24275 )  ;
assign n25606 =  ( n95 ) & ( n24277 )  ;
assign n25607 =  ( n95 ) & ( n24279 )  ;
assign n25608 =  ( n95 ) & ( n24281 )  ;
assign n25609 =  ( n95 ) & ( n24283 )  ;
assign n25610 =  ( n95 ) & ( n24285 )  ;
assign n25611 =  ( n95 ) & ( n24287 )  ;
assign n25612 =  ( n95 ) & ( n24289 )  ;
assign n25613 =  ( n96 ) & ( n24259 )  ;
assign n25614 =  ( n96 ) & ( n24261 )  ;
assign n25615 =  ( n96 ) & ( n24263 )  ;
assign n25616 =  ( n96 ) & ( n24265 )  ;
assign n25617 =  ( n96 ) & ( n24267 )  ;
assign n25618 =  ( n96 ) & ( n24269 )  ;
assign n25619 =  ( n96 ) & ( n24271 )  ;
assign n25620 =  ( n96 ) & ( n24273 )  ;
assign n25621 =  ( n96 ) & ( n24275 )  ;
assign n25622 =  ( n96 ) & ( n24277 )  ;
assign n25623 =  ( n96 ) & ( n24279 )  ;
assign n25624 =  ( n96 ) & ( n24281 )  ;
assign n25625 =  ( n96 ) & ( n24283 )  ;
assign n25626 =  ( n96 ) & ( n24285 )  ;
assign n25627 =  ( n96 ) & ( n24287 )  ;
assign n25628 =  ( n96 ) & ( n24289 )  ;
assign n25629 =  ( n97 ) & ( n24259 )  ;
assign n25630 =  ( n97 ) & ( n24261 )  ;
assign n25631 =  ( n97 ) & ( n24263 )  ;
assign n25632 =  ( n97 ) & ( n24265 )  ;
assign n25633 =  ( n97 ) & ( n24267 )  ;
assign n25634 =  ( n97 ) & ( n24269 )  ;
assign n25635 =  ( n97 ) & ( n24271 )  ;
assign n25636 =  ( n97 ) & ( n24273 )  ;
assign n25637 =  ( n97 ) & ( n24275 )  ;
assign n25638 =  ( n97 ) & ( n24277 )  ;
assign n25639 =  ( n97 ) & ( n24279 )  ;
assign n25640 =  ( n97 ) & ( n24281 )  ;
assign n25641 =  ( n97 ) & ( n24283 )  ;
assign n25642 =  ( n97 ) & ( n24285 )  ;
assign n25643 =  ( n97 ) & ( n24287 )  ;
assign n25644 =  ( n97 ) & ( n24289 )  ;
assign n25645 =  ( n98 ) & ( n24259 )  ;
assign n25646 =  ( n98 ) & ( n24261 )  ;
assign n25647 =  ( n98 ) & ( n24263 )  ;
assign n25648 =  ( n98 ) & ( n24265 )  ;
assign n25649 =  ( n98 ) & ( n24267 )  ;
assign n25650 =  ( n98 ) & ( n24269 )  ;
assign n25651 =  ( n98 ) & ( n24271 )  ;
assign n25652 =  ( n98 ) & ( n24273 )  ;
assign n25653 =  ( n98 ) & ( n24275 )  ;
assign n25654 =  ( n98 ) & ( n24277 )  ;
assign n25655 =  ( n98 ) & ( n24279 )  ;
assign n25656 =  ( n98 ) & ( n24281 )  ;
assign n25657 =  ( n98 ) & ( n24283 )  ;
assign n25658 =  ( n98 ) & ( n24285 )  ;
assign n25659 =  ( n98 ) & ( n24287 )  ;
assign n25660 =  ( n98 ) & ( n24289 )  ;
assign n25661 =  ( n99 ) & ( n24259 )  ;
assign n25662 =  ( n99 ) & ( n24261 )  ;
assign n25663 =  ( n99 ) & ( n24263 )  ;
assign n25664 =  ( n99 ) & ( n24265 )  ;
assign n25665 =  ( n99 ) & ( n24267 )  ;
assign n25666 =  ( n99 ) & ( n24269 )  ;
assign n25667 =  ( n99 ) & ( n24271 )  ;
assign n25668 =  ( n99 ) & ( n24273 )  ;
assign n25669 =  ( n99 ) & ( n24275 )  ;
assign n25670 =  ( n99 ) & ( n24277 )  ;
assign n25671 =  ( n99 ) & ( n24279 )  ;
assign n25672 =  ( n99 ) & ( n24281 )  ;
assign n25673 =  ( n99 ) & ( n24283 )  ;
assign n25674 =  ( n99 ) & ( n24285 )  ;
assign n25675 =  ( n99 ) & ( n24287 )  ;
assign n25676 =  ( n99 ) & ( n24289 )  ;
assign n25677 =  ( n100 ) & ( n24259 )  ;
assign n25678 =  ( n100 ) & ( n24261 )  ;
assign n25679 =  ( n100 ) & ( n24263 )  ;
assign n25680 =  ( n100 ) & ( n24265 )  ;
assign n25681 =  ( n100 ) & ( n24267 )  ;
assign n25682 =  ( n100 ) & ( n24269 )  ;
assign n25683 =  ( n100 ) & ( n24271 )  ;
assign n25684 =  ( n100 ) & ( n24273 )  ;
assign n25685 =  ( n100 ) & ( n24275 )  ;
assign n25686 =  ( n100 ) & ( n24277 )  ;
assign n25687 =  ( n100 ) & ( n24279 )  ;
assign n25688 =  ( n100 ) & ( n24281 )  ;
assign n25689 =  ( n100 ) & ( n24283 )  ;
assign n25690 =  ( n100 ) & ( n24285 )  ;
assign n25691 =  ( n100 ) & ( n24287 )  ;
assign n25692 =  ( n100 ) & ( n24289 )  ;
assign n25693 =  ( n101 ) & ( n24259 )  ;
assign n25694 =  ( n101 ) & ( n24261 )  ;
assign n25695 =  ( n101 ) & ( n24263 )  ;
assign n25696 =  ( n101 ) & ( n24265 )  ;
assign n25697 =  ( n101 ) & ( n24267 )  ;
assign n25698 =  ( n101 ) & ( n24269 )  ;
assign n25699 =  ( n101 ) & ( n24271 )  ;
assign n25700 =  ( n101 ) & ( n24273 )  ;
assign n25701 =  ( n101 ) & ( n24275 )  ;
assign n25702 =  ( n101 ) & ( n24277 )  ;
assign n25703 =  ( n101 ) & ( n24279 )  ;
assign n25704 =  ( n101 ) & ( n24281 )  ;
assign n25705 =  ( n101 ) & ( n24283 )  ;
assign n25706 =  ( n101 ) & ( n24285 )  ;
assign n25707 =  ( n101 ) & ( n24287 )  ;
assign n25708 =  ( n101 ) & ( n24289 )  ;
assign n25709 =  ( n102 ) & ( n24259 )  ;
assign n25710 =  ( n102 ) & ( n24261 )  ;
assign n25711 =  ( n102 ) & ( n24263 )  ;
assign n25712 =  ( n102 ) & ( n24265 )  ;
assign n25713 =  ( n102 ) & ( n24267 )  ;
assign n25714 =  ( n102 ) & ( n24269 )  ;
assign n25715 =  ( n102 ) & ( n24271 )  ;
assign n25716 =  ( n102 ) & ( n24273 )  ;
assign n25717 =  ( n102 ) & ( n24275 )  ;
assign n25718 =  ( n102 ) & ( n24277 )  ;
assign n25719 =  ( n102 ) & ( n24279 )  ;
assign n25720 =  ( n102 ) & ( n24281 )  ;
assign n25721 =  ( n102 ) & ( n24283 )  ;
assign n25722 =  ( n102 ) & ( n24285 )  ;
assign n25723 =  ( n102 ) & ( n24287 )  ;
assign n25724 =  ( n102 ) & ( n24289 )  ;
assign n25725 =  ( n103 ) & ( n24259 )  ;
assign n25726 =  ( n103 ) & ( n24261 )  ;
assign n25727 =  ( n103 ) & ( n24263 )  ;
assign n25728 =  ( n103 ) & ( n24265 )  ;
assign n25729 =  ( n103 ) & ( n24267 )  ;
assign n25730 =  ( n103 ) & ( n24269 )  ;
assign n25731 =  ( n103 ) & ( n24271 )  ;
assign n25732 =  ( n103 ) & ( n24273 )  ;
assign n25733 =  ( n103 ) & ( n24275 )  ;
assign n25734 =  ( n103 ) & ( n24277 )  ;
assign n25735 =  ( n103 ) & ( n24279 )  ;
assign n25736 =  ( n103 ) & ( n24281 )  ;
assign n25737 =  ( n103 ) & ( n24283 )  ;
assign n25738 =  ( n103 ) & ( n24285 )  ;
assign n25739 =  ( n103 ) & ( n24287 )  ;
assign n25740 =  ( n103 ) & ( n24289 )  ;
assign n25741 =  ( n104 ) & ( n24259 )  ;
assign n25742 =  ( n104 ) & ( n24261 )  ;
assign n25743 =  ( n104 ) & ( n24263 )  ;
assign n25744 =  ( n104 ) & ( n24265 )  ;
assign n25745 =  ( n104 ) & ( n24267 )  ;
assign n25746 =  ( n104 ) & ( n24269 )  ;
assign n25747 =  ( n104 ) & ( n24271 )  ;
assign n25748 =  ( n104 ) & ( n24273 )  ;
assign n25749 =  ( n104 ) & ( n24275 )  ;
assign n25750 =  ( n104 ) & ( n24277 )  ;
assign n25751 =  ( n104 ) & ( n24279 )  ;
assign n25752 =  ( n104 ) & ( n24281 )  ;
assign n25753 =  ( n104 ) & ( n24283 )  ;
assign n25754 =  ( n104 ) & ( n24285 )  ;
assign n25755 =  ( n104 ) & ( n24287 )  ;
assign n25756 =  ( n104 ) & ( n24289 )  ;
assign n25757 =  ( n105 ) & ( n24259 )  ;
assign n25758 =  ( n105 ) & ( n24261 )  ;
assign n25759 =  ( n105 ) & ( n24263 )  ;
assign n25760 =  ( n105 ) & ( n24265 )  ;
assign n25761 =  ( n105 ) & ( n24267 )  ;
assign n25762 =  ( n105 ) & ( n24269 )  ;
assign n25763 =  ( n105 ) & ( n24271 )  ;
assign n25764 =  ( n105 ) & ( n24273 )  ;
assign n25765 =  ( n105 ) & ( n24275 )  ;
assign n25766 =  ( n105 ) & ( n24277 )  ;
assign n25767 =  ( n105 ) & ( n24279 )  ;
assign n25768 =  ( n105 ) & ( n24281 )  ;
assign n25769 =  ( n105 ) & ( n24283 )  ;
assign n25770 =  ( n105 ) & ( n24285 )  ;
assign n25771 =  ( n105 ) & ( n24287 )  ;
assign n25772 =  ( n105 ) & ( n24289 )  ;
assign n25773 =  ( n106 ) & ( n24259 )  ;
assign n25774 =  ( n106 ) & ( n24261 )  ;
assign n25775 =  ( n106 ) & ( n24263 )  ;
assign n25776 =  ( n106 ) & ( n24265 )  ;
assign n25777 =  ( n106 ) & ( n24267 )  ;
assign n25778 =  ( n106 ) & ( n24269 )  ;
assign n25779 =  ( n106 ) & ( n24271 )  ;
assign n25780 =  ( n106 ) & ( n24273 )  ;
assign n25781 =  ( n106 ) & ( n24275 )  ;
assign n25782 =  ( n106 ) & ( n24277 )  ;
assign n25783 =  ( n106 ) & ( n24279 )  ;
assign n25784 =  ( n106 ) & ( n24281 )  ;
assign n25785 =  ( n106 ) & ( n24283 )  ;
assign n25786 =  ( n106 ) & ( n24285 )  ;
assign n25787 =  ( n106 ) & ( n24287 )  ;
assign n25788 =  ( n106 ) & ( n24289 )  ;
assign n25789 =  ( n107 ) & ( n24259 )  ;
assign n25790 =  ( n107 ) & ( n24261 )  ;
assign n25791 =  ( n107 ) & ( n24263 )  ;
assign n25792 =  ( n107 ) & ( n24265 )  ;
assign n25793 =  ( n107 ) & ( n24267 )  ;
assign n25794 =  ( n107 ) & ( n24269 )  ;
assign n25795 =  ( n107 ) & ( n24271 )  ;
assign n25796 =  ( n107 ) & ( n24273 )  ;
assign n25797 =  ( n107 ) & ( n24275 )  ;
assign n25798 =  ( n107 ) & ( n24277 )  ;
assign n25799 =  ( n107 ) & ( n24279 )  ;
assign n25800 =  ( n107 ) & ( n24281 )  ;
assign n25801 =  ( n107 ) & ( n24283 )  ;
assign n25802 =  ( n107 ) & ( n24285 )  ;
assign n25803 =  ( n107 ) & ( n24287 )  ;
assign n25804 =  ( n107 ) & ( n24289 )  ;
assign n25805 =  ( n108 ) & ( n24259 )  ;
assign n25806 =  ( n108 ) & ( n24261 )  ;
assign n25807 =  ( n108 ) & ( n24263 )  ;
assign n25808 =  ( n108 ) & ( n24265 )  ;
assign n25809 =  ( n108 ) & ( n24267 )  ;
assign n25810 =  ( n108 ) & ( n24269 )  ;
assign n25811 =  ( n108 ) & ( n24271 )  ;
assign n25812 =  ( n108 ) & ( n24273 )  ;
assign n25813 =  ( n108 ) & ( n24275 )  ;
assign n25814 =  ( n108 ) & ( n24277 )  ;
assign n25815 =  ( n108 ) & ( n24279 )  ;
assign n25816 =  ( n108 ) & ( n24281 )  ;
assign n25817 =  ( n108 ) & ( n24283 )  ;
assign n25818 =  ( n108 ) & ( n24285 )  ;
assign n25819 =  ( n108 ) & ( n24287 )  ;
assign n25820 =  ( n108 ) & ( n24289 )  ;
assign n25821 =  ( n25820 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n25822 =  ( n25819 ) ? ( VREG_0_1 ) : ( n25821 ) ;
assign n25823 =  ( n25818 ) ? ( VREG_0_2 ) : ( n25822 ) ;
assign n25824 =  ( n25817 ) ? ( VREG_0_3 ) : ( n25823 ) ;
assign n25825 =  ( n25816 ) ? ( VREG_0_4 ) : ( n25824 ) ;
assign n25826 =  ( n25815 ) ? ( VREG_0_5 ) : ( n25825 ) ;
assign n25827 =  ( n25814 ) ? ( VREG_0_6 ) : ( n25826 ) ;
assign n25828 =  ( n25813 ) ? ( VREG_0_7 ) : ( n25827 ) ;
assign n25829 =  ( n25812 ) ? ( VREG_0_8 ) : ( n25828 ) ;
assign n25830 =  ( n25811 ) ? ( VREG_0_9 ) : ( n25829 ) ;
assign n25831 =  ( n25810 ) ? ( VREG_0_10 ) : ( n25830 ) ;
assign n25832 =  ( n25809 ) ? ( VREG_0_11 ) : ( n25831 ) ;
assign n25833 =  ( n25808 ) ? ( VREG_0_12 ) : ( n25832 ) ;
assign n25834 =  ( n25807 ) ? ( VREG_0_13 ) : ( n25833 ) ;
assign n25835 =  ( n25806 ) ? ( VREG_0_14 ) : ( n25834 ) ;
assign n25836 =  ( n25805 ) ? ( VREG_0_15 ) : ( n25835 ) ;
assign n25837 =  ( n25804 ) ? ( VREG_1_0 ) : ( n25836 ) ;
assign n25838 =  ( n25803 ) ? ( VREG_1_1 ) : ( n25837 ) ;
assign n25839 =  ( n25802 ) ? ( VREG_1_2 ) : ( n25838 ) ;
assign n25840 =  ( n25801 ) ? ( VREG_1_3 ) : ( n25839 ) ;
assign n25841 =  ( n25800 ) ? ( VREG_1_4 ) : ( n25840 ) ;
assign n25842 =  ( n25799 ) ? ( VREG_1_5 ) : ( n25841 ) ;
assign n25843 =  ( n25798 ) ? ( VREG_1_6 ) : ( n25842 ) ;
assign n25844 =  ( n25797 ) ? ( VREG_1_7 ) : ( n25843 ) ;
assign n25845 =  ( n25796 ) ? ( VREG_1_8 ) : ( n25844 ) ;
assign n25846 =  ( n25795 ) ? ( VREG_1_9 ) : ( n25845 ) ;
assign n25847 =  ( n25794 ) ? ( VREG_1_10 ) : ( n25846 ) ;
assign n25848 =  ( n25793 ) ? ( VREG_1_11 ) : ( n25847 ) ;
assign n25849 =  ( n25792 ) ? ( VREG_1_12 ) : ( n25848 ) ;
assign n25850 =  ( n25791 ) ? ( VREG_1_13 ) : ( n25849 ) ;
assign n25851 =  ( n25790 ) ? ( VREG_1_14 ) : ( n25850 ) ;
assign n25852 =  ( n25789 ) ? ( VREG_1_15 ) : ( n25851 ) ;
assign n25853 =  ( n25788 ) ? ( VREG_2_0 ) : ( n25852 ) ;
assign n25854 =  ( n25787 ) ? ( VREG_2_1 ) : ( n25853 ) ;
assign n25855 =  ( n25786 ) ? ( VREG_2_2 ) : ( n25854 ) ;
assign n25856 =  ( n25785 ) ? ( VREG_2_3 ) : ( n25855 ) ;
assign n25857 =  ( n25784 ) ? ( VREG_2_4 ) : ( n25856 ) ;
assign n25858 =  ( n25783 ) ? ( VREG_2_5 ) : ( n25857 ) ;
assign n25859 =  ( n25782 ) ? ( VREG_2_6 ) : ( n25858 ) ;
assign n25860 =  ( n25781 ) ? ( VREG_2_7 ) : ( n25859 ) ;
assign n25861 =  ( n25780 ) ? ( VREG_2_8 ) : ( n25860 ) ;
assign n25862 =  ( n25779 ) ? ( VREG_2_9 ) : ( n25861 ) ;
assign n25863 =  ( n25778 ) ? ( VREG_2_10 ) : ( n25862 ) ;
assign n25864 =  ( n25777 ) ? ( VREG_2_11 ) : ( n25863 ) ;
assign n25865 =  ( n25776 ) ? ( VREG_2_12 ) : ( n25864 ) ;
assign n25866 =  ( n25775 ) ? ( VREG_2_13 ) : ( n25865 ) ;
assign n25867 =  ( n25774 ) ? ( VREG_2_14 ) : ( n25866 ) ;
assign n25868 =  ( n25773 ) ? ( VREG_2_15 ) : ( n25867 ) ;
assign n25869 =  ( n25772 ) ? ( VREG_3_0 ) : ( n25868 ) ;
assign n25870 =  ( n25771 ) ? ( VREG_3_1 ) : ( n25869 ) ;
assign n25871 =  ( n25770 ) ? ( VREG_3_2 ) : ( n25870 ) ;
assign n25872 =  ( n25769 ) ? ( VREG_3_3 ) : ( n25871 ) ;
assign n25873 =  ( n25768 ) ? ( VREG_3_4 ) : ( n25872 ) ;
assign n25874 =  ( n25767 ) ? ( VREG_3_5 ) : ( n25873 ) ;
assign n25875 =  ( n25766 ) ? ( VREG_3_6 ) : ( n25874 ) ;
assign n25876 =  ( n25765 ) ? ( VREG_3_7 ) : ( n25875 ) ;
assign n25877 =  ( n25764 ) ? ( VREG_3_8 ) : ( n25876 ) ;
assign n25878 =  ( n25763 ) ? ( VREG_3_9 ) : ( n25877 ) ;
assign n25879 =  ( n25762 ) ? ( VREG_3_10 ) : ( n25878 ) ;
assign n25880 =  ( n25761 ) ? ( VREG_3_11 ) : ( n25879 ) ;
assign n25881 =  ( n25760 ) ? ( VREG_3_12 ) : ( n25880 ) ;
assign n25882 =  ( n25759 ) ? ( VREG_3_13 ) : ( n25881 ) ;
assign n25883 =  ( n25758 ) ? ( VREG_3_14 ) : ( n25882 ) ;
assign n25884 =  ( n25757 ) ? ( VREG_3_15 ) : ( n25883 ) ;
assign n25885 =  ( n25756 ) ? ( VREG_4_0 ) : ( n25884 ) ;
assign n25886 =  ( n25755 ) ? ( VREG_4_1 ) : ( n25885 ) ;
assign n25887 =  ( n25754 ) ? ( VREG_4_2 ) : ( n25886 ) ;
assign n25888 =  ( n25753 ) ? ( VREG_4_3 ) : ( n25887 ) ;
assign n25889 =  ( n25752 ) ? ( VREG_4_4 ) : ( n25888 ) ;
assign n25890 =  ( n25751 ) ? ( VREG_4_5 ) : ( n25889 ) ;
assign n25891 =  ( n25750 ) ? ( VREG_4_6 ) : ( n25890 ) ;
assign n25892 =  ( n25749 ) ? ( VREG_4_7 ) : ( n25891 ) ;
assign n25893 =  ( n25748 ) ? ( VREG_4_8 ) : ( n25892 ) ;
assign n25894 =  ( n25747 ) ? ( VREG_4_9 ) : ( n25893 ) ;
assign n25895 =  ( n25746 ) ? ( VREG_4_10 ) : ( n25894 ) ;
assign n25896 =  ( n25745 ) ? ( VREG_4_11 ) : ( n25895 ) ;
assign n25897 =  ( n25744 ) ? ( VREG_4_12 ) : ( n25896 ) ;
assign n25898 =  ( n25743 ) ? ( VREG_4_13 ) : ( n25897 ) ;
assign n25899 =  ( n25742 ) ? ( VREG_4_14 ) : ( n25898 ) ;
assign n25900 =  ( n25741 ) ? ( VREG_4_15 ) : ( n25899 ) ;
assign n25901 =  ( n25740 ) ? ( VREG_5_0 ) : ( n25900 ) ;
assign n25902 =  ( n25739 ) ? ( VREG_5_1 ) : ( n25901 ) ;
assign n25903 =  ( n25738 ) ? ( VREG_5_2 ) : ( n25902 ) ;
assign n25904 =  ( n25737 ) ? ( VREG_5_3 ) : ( n25903 ) ;
assign n25905 =  ( n25736 ) ? ( VREG_5_4 ) : ( n25904 ) ;
assign n25906 =  ( n25735 ) ? ( VREG_5_5 ) : ( n25905 ) ;
assign n25907 =  ( n25734 ) ? ( VREG_5_6 ) : ( n25906 ) ;
assign n25908 =  ( n25733 ) ? ( VREG_5_7 ) : ( n25907 ) ;
assign n25909 =  ( n25732 ) ? ( VREG_5_8 ) : ( n25908 ) ;
assign n25910 =  ( n25731 ) ? ( VREG_5_9 ) : ( n25909 ) ;
assign n25911 =  ( n25730 ) ? ( VREG_5_10 ) : ( n25910 ) ;
assign n25912 =  ( n25729 ) ? ( VREG_5_11 ) : ( n25911 ) ;
assign n25913 =  ( n25728 ) ? ( VREG_5_12 ) : ( n25912 ) ;
assign n25914 =  ( n25727 ) ? ( VREG_5_13 ) : ( n25913 ) ;
assign n25915 =  ( n25726 ) ? ( VREG_5_14 ) : ( n25914 ) ;
assign n25916 =  ( n25725 ) ? ( VREG_5_15 ) : ( n25915 ) ;
assign n25917 =  ( n25724 ) ? ( VREG_6_0 ) : ( n25916 ) ;
assign n25918 =  ( n25723 ) ? ( VREG_6_1 ) : ( n25917 ) ;
assign n25919 =  ( n25722 ) ? ( VREG_6_2 ) : ( n25918 ) ;
assign n25920 =  ( n25721 ) ? ( VREG_6_3 ) : ( n25919 ) ;
assign n25921 =  ( n25720 ) ? ( VREG_6_4 ) : ( n25920 ) ;
assign n25922 =  ( n25719 ) ? ( VREG_6_5 ) : ( n25921 ) ;
assign n25923 =  ( n25718 ) ? ( VREG_6_6 ) : ( n25922 ) ;
assign n25924 =  ( n25717 ) ? ( VREG_6_7 ) : ( n25923 ) ;
assign n25925 =  ( n25716 ) ? ( VREG_6_8 ) : ( n25924 ) ;
assign n25926 =  ( n25715 ) ? ( VREG_6_9 ) : ( n25925 ) ;
assign n25927 =  ( n25714 ) ? ( VREG_6_10 ) : ( n25926 ) ;
assign n25928 =  ( n25713 ) ? ( VREG_6_11 ) : ( n25927 ) ;
assign n25929 =  ( n25712 ) ? ( VREG_6_12 ) : ( n25928 ) ;
assign n25930 =  ( n25711 ) ? ( VREG_6_13 ) : ( n25929 ) ;
assign n25931 =  ( n25710 ) ? ( VREG_6_14 ) : ( n25930 ) ;
assign n25932 =  ( n25709 ) ? ( VREG_6_15 ) : ( n25931 ) ;
assign n25933 =  ( n25708 ) ? ( VREG_7_0 ) : ( n25932 ) ;
assign n25934 =  ( n25707 ) ? ( VREG_7_1 ) : ( n25933 ) ;
assign n25935 =  ( n25706 ) ? ( VREG_7_2 ) : ( n25934 ) ;
assign n25936 =  ( n25705 ) ? ( VREG_7_3 ) : ( n25935 ) ;
assign n25937 =  ( n25704 ) ? ( VREG_7_4 ) : ( n25936 ) ;
assign n25938 =  ( n25703 ) ? ( VREG_7_5 ) : ( n25937 ) ;
assign n25939 =  ( n25702 ) ? ( VREG_7_6 ) : ( n25938 ) ;
assign n25940 =  ( n25701 ) ? ( VREG_7_7 ) : ( n25939 ) ;
assign n25941 =  ( n25700 ) ? ( VREG_7_8 ) : ( n25940 ) ;
assign n25942 =  ( n25699 ) ? ( VREG_7_9 ) : ( n25941 ) ;
assign n25943 =  ( n25698 ) ? ( VREG_7_10 ) : ( n25942 ) ;
assign n25944 =  ( n25697 ) ? ( VREG_7_11 ) : ( n25943 ) ;
assign n25945 =  ( n25696 ) ? ( VREG_7_12 ) : ( n25944 ) ;
assign n25946 =  ( n25695 ) ? ( VREG_7_13 ) : ( n25945 ) ;
assign n25947 =  ( n25694 ) ? ( VREG_7_14 ) : ( n25946 ) ;
assign n25948 =  ( n25693 ) ? ( VREG_7_15 ) : ( n25947 ) ;
assign n25949 =  ( n25692 ) ? ( VREG_8_0 ) : ( n25948 ) ;
assign n25950 =  ( n25691 ) ? ( VREG_8_1 ) : ( n25949 ) ;
assign n25951 =  ( n25690 ) ? ( VREG_8_2 ) : ( n25950 ) ;
assign n25952 =  ( n25689 ) ? ( VREG_8_3 ) : ( n25951 ) ;
assign n25953 =  ( n25688 ) ? ( VREG_8_4 ) : ( n25952 ) ;
assign n25954 =  ( n25687 ) ? ( VREG_8_5 ) : ( n25953 ) ;
assign n25955 =  ( n25686 ) ? ( VREG_8_6 ) : ( n25954 ) ;
assign n25956 =  ( n25685 ) ? ( VREG_8_7 ) : ( n25955 ) ;
assign n25957 =  ( n25684 ) ? ( VREG_8_8 ) : ( n25956 ) ;
assign n25958 =  ( n25683 ) ? ( VREG_8_9 ) : ( n25957 ) ;
assign n25959 =  ( n25682 ) ? ( VREG_8_10 ) : ( n25958 ) ;
assign n25960 =  ( n25681 ) ? ( VREG_8_11 ) : ( n25959 ) ;
assign n25961 =  ( n25680 ) ? ( VREG_8_12 ) : ( n25960 ) ;
assign n25962 =  ( n25679 ) ? ( VREG_8_13 ) : ( n25961 ) ;
assign n25963 =  ( n25678 ) ? ( VREG_8_14 ) : ( n25962 ) ;
assign n25964 =  ( n25677 ) ? ( VREG_8_15 ) : ( n25963 ) ;
assign n25965 =  ( n25676 ) ? ( VREG_9_0 ) : ( n25964 ) ;
assign n25966 =  ( n25675 ) ? ( VREG_9_1 ) : ( n25965 ) ;
assign n25967 =  ( n25674 ) ? ( VREG_9_2 ) : ( n25966 ) ;
assign n25968 =  ( n25673 ) ? ( VREG_9_3 ) : ( n25967 ) ;
assign n25969 =  ( n25672 ) ? ( VREG_9_4 ) : ( n25968 ) ;
assign n25970 =  ( n25671 ) ? ( VREG_9_5 ) : ( n25969 ) ;
assign n25971 =  ( n25670 ) ? ( VREG_9_6 ) : ( n25970 ) ;
assign n25972 =  ( n25669 ) ? ( VREG_9_7 ) : ( n25971 ) ;
assign n25973 =  ( n25668 ) ? ( VREG_9_8 ) : ( n25972 ) ;
assign n25974 =  ( n25667 ) ? ( VREG_9_9 ) : ( n25973 ) ;
assign n25975 =  ( n25666 ) ? ( VREG_9_10 ) : ( n25974 ) ;
assign n25976 =  ( n25665 ) ? ( VREG_9_11 ) : ( n25975 ) ;
assign n25977 =  ( n25664 ) ? ( VREG_9_12 ) : ( n25976 ) ;
assign n25978 =  ( n25663 ) ? ( VREG_9_13 ) : ( n25977 ) ;
assign n25979 =  ( n25662 ) ? ( VREG_9_14 ) : ( n25978 ) ;
assign n25980 =  ( n25661 ) ? ( VREG_9_15 ) : ( n25979 ) ;
assign n25981 =  ( n25660 ) ? ( VREG_10_0 ) : ( n25980 ) ;
assign n25982 =  ( n25659 ) ? ( VREG_10_1 ) : ( n25981 ) ;
assign n25983 =  ( n25658 ) ? ( VREG_10_2 ) : ( n25982 ) ;
assign n25984 =  ( n25657 ) ? ( VREG_10_3 ) : ( n25983 ) ;
assign n25985 =  ( n25656 ) ? ( VREG_10_4 ) : ( n25984 ) ;
assign n25986 =  ( n25655 ) ? ( VREG_10_5 ) : ( n25985 ) ;
assign n25987 =  ( n25654 ) ? ( VREG_10_6 ) : ( n25986 ) ;
assign n25988 =  ( n25653 ) ? ( VREG_10_7 ) : ( n25987 ) ;
assign n25989 =  ( n25652 ) ? ( VREG_10_8 ) : ( n25988 ) ;
assign n25990 =  ( n25651 ) ? ( VREG_10_9 ) : ( n25989 ) ;
assign n25991 =  ( n25650 ) ? ( VREG_10_10 ) : ( n25990 ) ;
assign n25992 =  ( n25649 ) ? ( VREG_10_11 ) : ( n25991 ) ;
assign n25993 =  ( n25648 ) ? ( VREG_10_12 ) : ( n25992 ) ;
assign n25994 =  ( n25647 ) ? ( VREG_10_13 ) : ( n25993 ) ;
assign n25995 =  ( n25646 ) ? ( VREG_10_14 ) : ( n25994 ) ;
assign n25996 =  ( n25645 ) ? ( VREG_10_15 ) : ( n25995 ) ;
assign n25997 =  ( n25644 ) ? ( VREG_11_0 ) : ( n25996 ) ;
assign n25998 =  ( n25643 ) ? ( VREG_11_1 ) : ( n25997 ) ;
assign n25999 =  ( n25642 ) ? ( VREG_11_2 ) : ( n25998 ) ;
assign n26000 =  ( n25641 ) ? ( VREG_11_3 ) : ( n25999 ) ;
assign n26001 =  ( n25640 ) ? ( VREG_11_4 ) : ( n26000 ) ;
assign n26002 =  ( n25639 ) ? ( VREG_11_5 ) : ( n26001 ) ;
assign n26003 =  ( n25638 ) ? ( VREG_11_6 ) : ( n26002 ) ;
assign n26004 =  ( n25637 ) ? ( VREG_11_7 ) : ( n26003 ) ;
assign n26005 =  ( n25636 ) ? ( VREG_11_8 ) : ( n26004 ) ;
assign n26006 =  ( n25635 ) ? ( VREG_11_9 ) : ( n26005 ) ;
assign n26007 =  ( n25634 ) ? ( VREG_11_10 ) : ( n26006 ) ;
assign n26008 =  ( n25633 ) ? ( VREG_11_11 ) : ( n26007 ) ;
assign n26009 =  ( n25632 ) ? ( VREG_11_12 ) : ( n26008 ) ;
assign n26010 =  ( n25631 ) ? ( VREG_11_13 ) : ( n26009 ) ;
assign n26011 =  ( n25630 ) ? ( VREG_11_14 ) : ( n26010 ) ;
assign n26012 =  ( n25629 ) ? ( VREG_11_15 ) : ( n26011 ) ;
assign n26013 =  ( n25628 ) ? ( VREG_12_0 ) : ( n26012 ) ;
assign n26014 =  ( n25627 ) ? ( VREG_12_1 ) : ( n26013 ) ;
assign n26015 =  ( n25626 ) ? ( VREG_12_2 ) : ( n26014 ) ;
assign n26016 =  ( n25625 ) ? ( VREG_12_3 ) : ( n26015 ) ;
assign n26017 =  ( n25624 ) ? ( VREG_12_4 ) : ( n26016 ) ;
assign n26018 =  ( n25623 ) ? ( VREG_12_5 ) : ( n26017 ) ;
assign n26019 =  ( n25622 ) ? ( VREG_12_6 ) : ( n26018 ) ;
assign n26020 =  ( n25621 ) ? ( VREG_12_7 ) : ( n26019 ) ;
assign n26021 =  ( n25620 ) ? ( VREG_12_8 ) : ( n26020 ) ;
assign n26022 =  ( n25619 ) ? ( VREG_12_9 ) : ( n26021 ) ;
assign n26023 =  ( n25618 ) ? ( VREG_12_10 ) : ( n26022 ) ;
assign n26024 =  ( n25617 ) ? ( VREG_12_11 ) : ( n26023 ) ;
assign n26025 =  ( n25616 ) ? ( VREG_12_12 ) : ( n26024 ) ;
assign n26026 =  ( n25615 ) ? ( VREG_12_13 ) : ( n26025 ) ;
assign n26027 =  ( n25614 ) ? ( VREG_12_14 ) : ( n26026 ) ;
assign n26028 =  ( n25613 ) ? ( VREG_12_15 ) : ( n26027 ) ;
assign n26029 =  ( n25612 ) ? ( VREG_13_0 ) : ( n26028 ) ;
assign n26030 =  ( n25611 ) ? ( VREG_13_1 ) : ( n26029 ) ;
assign n26031 =  ( n25610 ) ? ( VREG_13_2 ) : ( n26030 ) ;
assign n26032 =  ( n25609 ) ? ( VREG_13_3 ) : ( n26031 ) ;
assign n26033 =  ( n25608 ) ? ( VREG_13_4 ) : ( n26032 ) ;
assign n26034 =  ( n25607 ) ? ( VREG_13_5 ) : ( n26033 ) ;
assign n26035 =  ( n25606 ) ? ( VREG_13_6 ) : ( n26034 ) ;
assign n26036 =  ( n25605 ) ? ( VREG_13_7 ) : ( n26035 ) ;
assign n26037 =  ( n25604 ) ? ( VREG_13_8 ) : ( n26036 ) ;
assign n26038 =  ( n25603 ) ? ( VREG_13_9 ) : ( n26037 ) ;
assign n26039 =  ( n25602 ) ? ( VREG_13_10 ) : ( n26038 ) ;
assign n26040 =  ( n25601 ) ? ( VREG_13_11 ) : ( n26039 ) ;
assign n26041 =  ( n25600 ) ? ( VREG_13_12 ) : ( n26040 ) ;
assign n26042 =  ( n25599 ) ? ( VREG_13_13 ) : ( n26041 ) ;
assign n26043 =  ( n25598 ) ? ( VREG_13_14 ) : ( n26042 ) ;
assign n26044 =  ( n25597 ) ? ( VREG_13_15 ) : ( n26043 ) ;
assign n26045 =  ( n25596 ) ? ( VREG_14_0 ) : ( n26044 ) ;
assign n26046 =  ( n25595 ) ? ( VREG_14_1 ) : ( n26045 ) ;
assign n26047 =  ( n25594 ) ? ( VREG_14_2 ) : ( n26046 ) ;
assign n26048 =  ( n25593 ) ? ( VREG_14_3 ) : ( n26047 ) ;
assign n26049 =  ( n25592 ) ? ( VREG_14_4 ) : ( n26048 ) ;
assign n26050 =  ( n25591 ) ? ( VREG_14_5 ) : ( n26049 ) ;
assign n26051 =  ( n25590 ) ? ( VREG_14_6 ) : ( n26050 ) ;
assign n26052 =  ( n25589 ) ? ( VREG_14_7 ) : ( n26051 ) ;
assign n26053 =  ( n25588 ) ? ( VREG_14_8 ) : ( n26052 ) ;
assign n26054 =  ( n25587 ) ? ( VREG_14_9 ) : ( n26053 ) ;
assign n26055 =  ( n25586 ) ? ( VREG_14_10 ) : ( n26054 ) ;
assign n26056 =  ( n25585 ) ? ( VREG_14_11 ) : ( n26055 ) ;
assign n26057 =  ( n25584 ) ? ( VREG_14_12 ) : ( n26056 ) ;
assign n26058 =  ( n25583 ) ? ( VREG_14_13 ) : ( n26057 ) ;
assign n26059 =  ( n25582 ) ? ( VREG_14_14 ) : ( n26058 ) ;
assign n26060 =  ( n25581 ) ? ( VREG_14_15 ) : ( n26059 ) ;
assign n26061 =  ( n25580 ) ? ( VREG_15_0 ) : ( n26060 ) ;
assign n26062 =  ( n25579 ) ? ( VREG_15_1 ) : ( n26061 ) ;
assign n26063 =  ( n25578 ) ? ( VREG_15_2 ) : ( n26062 ) ;
assign n26064 =  ( n25577 ) ? ( VREG_15_3 ) : ( n26063 ) ;
assign n26065 =  ( n25576 ) ? ( VREG_15_4 ) : ( n26064 ) ;
assign n26066 =  ( n25575 ) ? ( VREG_15_5 ) : ( n26065 ) ;
assign n26067 =  ( n25574 ) ? ( VREG_15_6 ) : ( n26066 ) ;
assign n26068 =  ( n25573 ) ? ( VREG_15_7 ) : ( n26067 ) ;
assign n26069 =  ( n25572 ) ? ( VREG_15_8 ) : ( n26068 ) ;
assign n26070 =  ( n25571 ) ? ( VREG_15_9 ) : ( n26069 ) ;
assign n26071 =  ( n25570 ) ? ( VREG_15_10 ) : ( n26070 ) ;
assign n26072 =  ( n25569 ) ? ( VREG_15_11 ) : ( n26071 ) ;
assign n26073 =  ( n25568 ) ? ( VREG_15_12 ) : ( n26072 ) ;
assign n26074 =  ( n25567 ) ? ( VREG_15_13 ) : ( n26073 ) ;
assign n26075 =  ( n25566 ) ? ( VREG_15_14 ) : ( n26074 ) ;
assign n26076 =  ( n25565 ) ? ( VREG_15_15 ) : ( n26075 ) ;
assign n26077 =  ( n25564 ) ? ( VREG_16_0 ) : ( n26076 ) ;
assign n26078 =  ( n25563 ) ? ( VREG_16_1 ) : ( n26077 ) ;
assign n26079 =  ( n25562 ) ? ( VREG_16_2 ) : ( n26078 ) ;
assign n26080 =  ( n25561 ) ? ( VREG_16_3 ) : ( n26079 ) ;
assign n26081 =  ( n25560 ) ? ( VREG_16_4 ) : ( n26080 ) ;
assign n26082 =  ( n25559 ) ? ( VREG_16_5 ) : ( n26081 ) ;
assign n26083 =  ( n25558 ) ? ( VREG_16_6 ) : ( n26082 ) ;
assign n26084 =  ( n25557 ) ? ( VREG_16_7 ) : ( n26083 ) ;
assign n26085 =  ( n25556 ) ? ( VREG_16_8 ) : ( n26084 ) ;
assign n26086 =  ( n25555 ) ? ( VREG_16_9 ) : ( n26085 ) ;
assign n26087 =  ( n25554 ) ? ( VREG_16_10 ) : ( n26086 ) ;
assign n26088 =  ( n25553 ) ? ( VREG_16_11 ) : ( n26087 ) ;
assign n26089 =  ( n25552 ) ? ( VREG_16_12 ) : ( n26088 ) ;
assign n26090 =  ( n25551 ) ? ( VREG_16_13 ) : ( n26089 ) ;
assign n26091 =  ( n25550 ) ? ( VREG_16_14 ) : ( n26090 ) ;
assign n26092 =  ( n25549 ) ? ( VREG_16_15 ) : ( n26091 ) ;
assign n26093 =  ( n25548 ) ? ( VREG_17_0 ) : ( n26092 ) ;
assign n26094 =  ( n25547 ) ? ( VREG_17_1 ) : ( n26093 ) ;
assign n26095 =  ( n25546 ) ? ( VREG_17_2 ) : ( n26094 ) ;
assign n26096 =  ( n25545 ) ? ( VREG_17_3 ) : ( n26095 ) ;
assign n26097 =  ( n25544 ) ? ( VREG_17_4 ) : ( n26096 ) ;
assign n26098 =  ( n25543 ) ? ( VREG_17_5 ) : ( n26097 ) ;
assign n26099 =  ( n25542 ) ? ( VREG_17_6 ) : ( n26098 ) ;
assign n26100 =  ( n25541 ) ? ( VREG_17_7 ) : ( n26099 ) ;
assign n26101 =  ( n25540 ) ? ( VREG_17_8 ) : ( n26100 ) ;
assign n26102 =  ( n25539 ) ? ( VREG_17_9 ) : ( n26101 ) ;
assign n26103 =  ( n25538 ) ? ( VREG_17_10 ) : ( n26102 ) ;
assign n26104 =  ( n25537 ) ? ( VREG_17_11 ) : ( n26103 ) ;
assign n26105 =  ( n25536 ) ? ( VREG_17_12 ) : ( n26104 ) ;
assign n26106 =  ( n25535 ) ? ( VREG_17_13 ) : ( n26105 ) ;
assign n26107 =  ( n25534 ) ? ( VREG_17_14 ) : ( n26106 ) ;
assign n26108 =  ( n25533 ) ? ( VREG_17_15 ) : ( n26107 ) ;
assign n26109 =  ( n25532 ) ? ( VREG_18_0 ) : ( n26108 ) ;
assign n26110 =  ( n25531 ) ? ( VREG_18_1 ) : ( n26109 ) ;
assign n26111 =  ( n25530 ) ? ( VREG_18_2 ) : ( n26110 ) ;
assign n26112 =  ( n25529 ) ? ( VREG_18_3 ) : ( n26111 ) ;
assign n26113 =  ( n25528 ) ? ( VREG_18_4 ) : ( n26112 ) ;
assign n26114 =  ( n25527 ) ? ( VREG_18_5 ) : ( n26113 ) ;
assign n26115 =  ( n25526 ) ? ( VREG_18_6 ) : ( n26114 ) ;
assign n26116 =  ( n25525 ) ? ( VREG_18_7 ) : ( n26115 ) ;
assign n26117 =  ( n25524 ) ? ( VREG_18_8 ) : ( n26116 ) ;
assign n26118 =  ( n25523 ) ? ( VREG_18_9 ) : ( n26117 ) ;
assign n26119 =  ( n25522 ) ? ( VREG_18_10 ) : ( n26118 ) ;
assign n26120 =  ( n25521 ) ? ( VREG_18_11 ) : ( n26119 ) ;
assign n26121 =  ( n25520 ) ? ( VREG_18_12 ) : ( n26120 ) ;
assign n26122 =  ( n25519 ) ? ( VREG_18_13 ) : ( n26121 ) ;
assign n26123 =  ( n25518 ) ? ( VREG_18_14 ) : ( n26122 ) ;
assign n26124 =  ( n25517 ) ? ( VREG_18_15 ) : ( n26123 ) ;
assign n26125 =  ( n25516 ) ? ( VREG_19_0 ) : ( n26124 ) ;
assign n26126 =  ( n25515 ) ? ( VREG_19_1 ) : ( n26125 ) ;
assign n26127 =  ( n25514 ) ? ( VREG_19_2 ) : ( n26126 ) ;
assign n26128 =  ( n25513 ) ? ( VREG_19_3 ) : ( n26127 ) ;
assign n26129 =  ( n25512 ) ? ( VREG_19_4 ) : ( n26128 ) ;
assign n26130 =  ( n25511 ) ? ( VREG_19_5 ) : ( n26129 ) ;
assign n26131 =  ( n25510 ) ? ( VREG_19_6 ) : ( n26130 ) ;
assign n26132 =  ( n25509 ) ? ( VREG_19_7 ) : ( n26131 ) ;
assign n26133 =  ( n25508 ) ? ( VREG_19_8 ) : ( n26132 ) ;
assign n26134 =  ( n25507 ) ? ( VREG_19_9 ) : ( n26133 ) ;
assign n26135 =  ( n25506 ) ? ( VREG_19_10 ) : ( n26134 ) ;
assign n26136 =  ( n25505 ) ? ( VREG_19_11 ) : ( n26135 ) ;
assign n26137 =  ( n25504 ) ? ( VREG_19_12 ) : ( n26136 ) ;
assign n26138 =  ( n25503 ) ? ( VREG_19_13 ) : ( n26137 ) ;
assign n26139 =  ( n25502 ) ? ( VREG_19_14 ) : ( n26138 ) ;
assign n26140 =  ( n25501 ) ? ( VREG_19_15 ) : ( n26139 ) ;
assign n26141 =  ( n25500 ) ? ( VREG_20_0 ) : ( n26140 ) ;
assign n26142 =  ( n25499 ) ? ( VREG_20_1 ) : ( n26141 ) ;
assign n26143 =  ( n25498 ) ? ( VREG_20_2 ) : ( n26142 ) ;
assign n26144 =  ( n25497 ) ? ( VREG_20_3 ) : ( n26143 ) ;
assign n26145 =  ( n25496 ) ? ( VREG_20_4 ) : ( n26144 ) ;
assign n26146 =  ( n25495 ) ? ( VREG_20_5 ) : ( n26145 ) ;
assign n26147 =  ( n25494 ) ? ( VREG_20_6 ) : ( n26146 ) ;
assign n26148 =  ( n25493 ) ? ( VREG_20_7 ) : ( n26147 ) ;
assign n26149 =  ( n25492 ) ? ( VREG_20_8 ) : ( n26148 ) ;
assign n26150 =  ( n25491 ) ? ( VREG_20_9 ) : ( n26149 ) ;
assign n26151 =  ( n25490 ) ? ( VREG_20_10 ) : ( n26150 ) ;
assign n26152 =  ( n25489 ) ? ( VREG_20_11 ) : ( n26151 ) ;
assign n26153 =  ( n25488 ) ? ( VREG_20_12 ) : ( n26152 ) ;
assign n26154 =  ( n25487 ) ? ( VREG_20_13 ) : ( n26153 ) ;
assign n26155 =  ( n25486 ) ? ( VREG_20_14 ) : ( n26154 ) ;
assign n26156 =  ( n25485 ) ? ( VREG_20_15 ) : ( n26155 ) ;
assign n26157 =  ( n25484 ) ? ( VREG_21_0 ) : ( n26156 ) ;
assign n26158 =  ( n25483 ) ? ( VREG_21_1 ) : ( n26157 ) ;
assign n26159 =  ( n25482 ) ? ( VREG_21_2 ) : ( n26158 ) ;
assign n26160 =  ( n25481 ) ? ( VREG_21_3 ) : ( n26159 ) ;
assign n26161 =  ( n25480 ) ? ( VREG_21_4 ) : ( n26160 ) ;
assign n26162 =  ( n25479 ) ? ( VREG_21_5 ) : ( n26161 ) ;
assign n26163 =  ( n25478 ) ? ( VREG_21_6 ) : ( n26162 ) ;
assign n26164 =  ( n25477 ) ? ( VREG_21_7 ) : ( n26163 ) ;
assign n26165 =  ( n25476 ) ? ( VREG_21_8 ) : ( n26164 ) ;
assign n26166 =  ( n25475 ) ? ( VREG_21_9 ) : ( n26165 ) ;
assign n26167 =  ( n25474 ) ? ( VREG_21_10 ) : ( n26166 ) ;
assign n26168 =  ( n25473 ) ? ( VREG_21_11 ) : ( n26167 ) ;
assign n26169 =  ( n25472 ) ? ( VREG_21_12 ) : ( n26168 ) ;
assign n26170 =  ( n25471 ) ? ( VREG_21_13 ) : ( n26169 ) ;
assign n26171 =  ( n25470 ) ? ( VREG_21_14 ) : ( n26170 ) ;
assign n26172 =  ( n25469 ) ? ( VREG_21_15 ) : ( n26171 ) ;
assign n26173 =  ( n25468 ) ? ( VREG_22_0 ) : ( n26172 ) ;
assign n26174 =  ( n25467 ) ? ( VREG_22_1 ) : ( n26173 ) ;
assign n26175 =  ( n25466 ) ? ( VREG_22_2 ) : ( n26174 ) ;
assign n26176 =  ( n25465 ) ? ( VREG_22_3 ) : ( n26175 ) ;
assign n26177 =  ( n25464 ) ? ( VREG_22_4 ) : ( n26176 ) ;
assign n26178 =  ( n25463 ) ? ( VREG_22_5 ) : ( n26177 ) ;
assign n26179 =  ( n25462 ) ? ( VREG_22_6 ) : ( n26178 ) ;
assign n26180 =  ( n25461 ) ? ( VREG_22_7 ) : ( n26179 ) ;
assign n26181 =  ( n25460 ) ? ( VREG_22_8 ) : ( n26180 ) ;
assign n26182 =  ( n25459 ) ? ( VREG_22_9 ) : ( n26181 ) ;
assign n26183 =  ( n25458 ) ? ( VREG_22_10 ) : ( n26182 ) ;
assign n26184 =  ( n25457 ) ? ( VREG_22_11 ) : ( n26183 ) ;
assign n26185 =  ( n25456 ) ? ( VREG_22_12 ) : ( n26184 ) ;
assign n26186 =  ( n25455 ) ? ( VREG_22_13 ) : ( n26185 ) ;
assign n26187 =  ( n25454 ) ? ( VREG_22_14 ) : ( n26186 ) ;
assign n26188 =  ( n25453 ) ? ( VREG_22_15 ) : ( n26187 ) ;
assign n26189 =  ( n25452 ) ? ( VREG_23_0 ) : ( n26188 ) ;
assign n26190 =  ( n25451 ) ? ( VREG_23_1 ) : ( n26189 ) ;
assign n26191 =  ( n25450 ) ? ( VREG_23_2 ) : ( n26190 ) ;
assign n26192 =  ( n25449 ) ? ( VREG_23_3 ) : ( n26191 ) ;
assign n26193 =  ( n25448 ) ? ( VREG_23_4 ) : ( n26192 ) ;
assign n26194 =  ( n25447 ) ? ( VREG_23_5 ) : ( n26193 ) ;
assign n26195 =  ( n25446 ) ? ( VREG_23_6 ) : ( n26194 ) ;
assign n26196 =  ( n25445 ) ? ( VREG_23_7 ) : ( n26195 ) ;
assign n26197 =  ( n25444 ) ? ( VREG_23_8 ) : ( n26196 ) ;
assign n26198 =  ( n25443 ) ? ( VREG_23_9 ) : ( n26197 ) ;
assign n26199 =  ( n25442 ) ? ( VREG_23_10 ) : ( n26198 ) ;
assign n26200 =  ( n25441 ) ? ( VREG_23_11 ) : ( n26199 ) ;
assign n26201 =  ( n25440 ) ? ( VREG_23_12 ) : ( n26200 ) ;
assign n26202 =  ( n25439 ) ? ( VREG_23_13 ) : ( n26201 ) ;
assign n26203 =  ( n25438 ) ? ( VREG_23_14 ) : ( n26202 ) ;
assign n26204 =  ( n25437 ) ? ( VREG_23_15 ) : ( n26203 ) ;
assign n26205 =  ( n25436 ) ? ( VREG_24_0 ) : ( n26204 ) ;
assign n26206 =  ( n25435 ) ? ( VREG_24_1 ) : ( n26205 ) ;
assign n26207 =  ( n25434 ) ? ( VREG_24_2 ) : ( n26206 ) ;
assign n26208 =  ( n25433 ) ? ( VREG_24_3 ) : ( n26207 ) ;
assign n26209 =  ( n25432 ) ? ( VREG_24_4 ) : ( n26208 ) ;
assign n26210 =  ( n25431 ) ? ( VREG_24_5 ) : ( n26209 ) ;
assign n26211 =  ( n25430 ) ? ( VREG_24_6 ) : ( n26210 ) ;
assign n26212 =  ( n25429 ) ? ( VREG_24_7 ) : ( n26211 ) ;
assign n26213 =  ( n25428 ) ? ( VREG_24_8 ) : ( n26212 ) ;
assign n26214 =  ( n25427 ) ? ( VREG_24_9 ) : ( n26213 ) ;
assign n26215 =  ( n25426 ) ? ( VREG_24_10 ) : ( n26214 ) ;
assign n26216 =  ( n25425 ) ? ( VREG_24_11 ) : ( n26215 ) ;
assign n26217 =  ( n25424 ) ? ( VREG_24_12 ) : ( n26216 ) ;
assign n26218 =  ( n25423 ) ? ( VREG_24_13 ) : ( n26217 ) ;
assign n26219 =  ( n25422 ) ? ( VREG_24_14 ) : ( n26218 ) ;
assign n26220 =  ( n25421 ) ? ( VREG_24_15 ) : ( n26219 ) ;
assign n26221 =  ( n25420 ) ? ( VREG_25_0 ) : ( n26220 ) ;
assign n26222 =  ( n25419 ) ? ( VREG_25_1 ) : ( n26221 ) ;
assign n26223 =  ( n25418 ) ? ( VREG_25_2 ) : ( n26222 ) ;
assign n26224 =  ( n25417 ) ? ( VREG_25_3 ) : ( n26223 ) ;
assign n26225 =  ( n25416 ) ? ( VREG_25_4 ) : ( n26224 ) ;
assign n26226 =  ( n25415 ) ? ( VREG_25_5 ) : ( n26225 ) ;
assign n26227 =  ( n25414 ) ? ( VREG_25_6 ) : ( n26226 ) ;
assign n26228 =  ( n25413 ) ? ( VREG_25_7 ) : ( n26227 ) ;
assign n26229 =  ( n25412 ) ? ( VREG_25_8 ) : ( n26228 ) ;
assign n26230 =  ( n25411 ) ? ( VREG_25_9 ) : ( n26229 ) ;
assign n26231 =  ( n25410 ) ? ( VREG_25_10 ) : ( n26230 ) ;
assign n26232 =  ( n25409 ) ? ( VREG_25_11 ) : ( n26231 ) ;
assign n26233 =  ( n25408 ) ? ( VREG_25_12 ) : ( n26232 ) ;
assign n26234 =  ( n25407 ) ? ( VREG_25_13 ) : ( n26233 ) ;
assign n26235 =  ( n25406 ) ? ( VREG_25_14 ) : ( n26234 ) ;
assign n26236 =  ( n25405 ) ? ( VREG_25_15 ) : ( n26235 ) ;
assign n26237 =  ( n25404 ) ? ( VREG_26_0 ) : ( n26236 ) ;
assign n26238 =  ( n25403 ) ? ( VREG_26_1 ) : ( n26237 ) ;
assign n26239 =  ( n25402 ) ? ( VREG_26_2 ) : ( n26238 ) ;
assign n26240 =  ( n25401 ) ? ( VREG_26_3 ) : ( n26239 ) ;
assign n26241 =  ( n25400 ) ? ( VREG_26_4 ) : ( n26240 ) ;
assign n26242 =  ( n25399 ) ? ( VREG_26_5 ) : ( n26241 ) ;
assign n26243 =  ( n25398 ) ? ( VREG_26_6 ) : ( n26242 ) ;
assign n26244 =  ( n25397 ) ? ( VREG_26_7 ) : ( n26243 ) ;
assign n26245 =  ( n25396 ) ? ( VREG_26_8 ) : ( n26244 ) ;
assign n26246 =  ( n25395 ) ? ( VREG_26_9 ) : ( n26245 ) ;
assign n26247 =  ( n25394 ) ? ( VREG_26_10 ) : ( n26246 ) ;
assign n26248 =  ( n25393 ) ? ( VREG_26_11 ) : ( n26247 ) ;
assign n26249 =  ( n25392 ) ? ( VREG_26_12 ) : ( n26248 ) ;
assign n26250 =  ( n25391 ) ? ( VREG_26_13 ) : ( n26249 ) ;
assign n26251 =  ( n25390 ) ? ( VREG_26_14 ) : ( n26250 ) ;
assign n26252 =  ( n25389 ) ? ( VREG_26_15 ) : ( n26251 ) ;
assign n26253 =  ( n25388 ) ? ( VREG_27_0 ) : ( n26252 ) ;
assign n26254 =  ( n25387 ) ? ( VREG_27_1 ) : ( n26253 ) ;
assign n26255 =  ( n25386 ) ? ( VREG_27_2 ) : ( n26254 ) ;
assign n26256 =  ( n25385 ) ? ( VREG_27_3 ) : ( n26255 ) ;
assign n26257 =  ( n25384 ) ? ( VREG_27_4 ) : ( n26256 ) ;
assign n26258 =  ( n25383 ) ? ( VREG_27_5 ) : ( n26257 ) ;
assign n26259 =  ( n25382 ) ? ( VREG_27_6 ) : ( n26258 ) ;
assign n26260 =  ( n25381 ) ? ( VREG_27_7 ) : ( n26259 ) ;
assign n26261 =  ( n25380 ) ? ( VREG_27_8 ) : ( n26260 ) ;
assign n26262 =  ( n25379 ) ? ( VREG_27_9 ) : ( n26261 ) ;
assign n26263 =  ( n25378 ) ? ( VREG_27_10 ) : ( n26262 ) ;
assign n26264 =  ( n25377 ) ? ( VREG_27_11 ) : ( n26263 ) ;
assign n26265 =  ( n25376 ) ? ( VREG_27_12 ) : ( n26264 ) ;
assign n26266 =  ( n25375 ) ? ( VREG_27_13 ) : ( n26265 ) ;
assign n26267 =  ( n25374 ) ? ( VREG_27_14 ) : ( n26266 ) ;
assign n26268 =  ( n25373 ) ? ( VREG_27_15 ) : ( n26267 ) ;
assign n26269 =  ( n25372 ) ? ( VREG_28_0 ) : ( n26268 ) ;
assign n26270 =  ( n25371 ) ? ( VREG_28_1 ) : ( n26269 ) ;
assign n26271 =  ( n25370 ) ? ( VREG_28_2 ) : ( n26270 ) ;
assign n26272 =  ( n25369 ) ? ( VREG_28_3 ) : ( n26271 ) ;
assign n26273 =  ( n25368 ) ? ( VREG_28_4 ) : ( n26272 ) ;
assign n26274 =  ( n25367 ) ? ( VREG_28_5 ) : ( n26273 ) ;
assign n26275 =  ( n25366 ) ? ( VREG_28_6 ) : ( n26274 ) ;
assign n26276 =  ( n25365 ) ? ( VREG_28_7 ) : ( n26275 ) ;
assign n26277 =  ( n25364 ) ? ( VREG_28_8 ) : ( n26276 ) ;
assign n26278 =  ( n25363 ) ? ( VREG_28_9 ) : ( n26277 ) ;
assign n26279 =  ( n25362 ) ? ( VREG_28_10 ) : ( n26278 ) ;
assign n26280 =  ( n25361 ) ? ( VREG_28_11 ) : ( n26279 ) ;
assign n26281 =  ( n25360 ) ? ( VREG_28_12 ) : ( n26280 ) ;
assign n26282 =  ( n25359 ) ? ( VREG_28_13 ) : ( n26281 ) ;
assign n26283 =  ( n25358 ) ? ( VREG_28_14 ) : ( n26282 ) ;
assign n26284 =  ( n25357 ) ? ( VREG_28_15 ) : ( n26283 ) ;
assign n26285 =  ( n25356 ) ? ( VREG_29_0 ) : ( n26284 ) ;
assign n26286 =  ( n25355 ) ? ( VREG_29_1 ) : ( n26285 ) ;
assign n26287 =  ( n25354 ) ? ( VREG_29_2 ) : ( n26286 ) ;
assign n26288 =  ( n25353 ) ? ( VREG_29_3 ) : ( n26287 ) ;
assign n26289 =  ( n25352 ) ? ( VREG_29_4 ) : ( n26288 ) ;
assign n26290 =  ( n25351 ) ? ( VREG_29_5 ) : ( n26289 ) ;
assign n26291 =  ( n25350 ) ? ( VREG_29_6 ) : ( n26290 ) ;
assign n26292 =  ( n25349 ) ? ( VREG_29_7 ) : ( n26291 ) ;
assign n26293 =  ( n25348 ) ? ( VREG_29_8 ) : ( n26292 ) ;
assign n26294 =  ( n25347 ) ? ( VREG_29_9 ) : ( n26293 ) ;
assign n26295 =  ( n25346 ) ? ( VREG_29_10 ) : ( n26294 ) ;
assign n26296 =  ( n25345 ) ? ( VREG_29_11 ) : ( n26295 ) ;
assign n26297 =  ( n25344 ) ? ( VREG_29_12 ) : ( n26296 ) ;
assign n26298 =  ( n25343 ) ? ( VREG_29_13 ) : ( n26297 ) ;
assign n26299 =  ( n25342 ) ? ( VREG_29_14 ) : ( n26298 ) ;
assign n26300 =  ( n25341 ) ? ( VREG_29_15 ) : ( n26299 ) ;
assign n26301 =  ( n25340 ) ? ( VREG_30_0 ) : ( n26300 ) ;
assign n26302 =  ( n25339 ) ? ( VREG_30_1 ) : ( n26301 ) ;
assign n26303 =  ( n25338 ) ? ( VREG_30_2 ) : ( n26302 ) ;
assign n26304 =  ( n25337 ) ? ( VREG_30_3 ) : ( n26303 ) ;
assign n26305 =  ( n25336 ) ? ( VREG_30_4 ) : ( n26304 ) ;
assign n26306 =  ( n25335 ) ? ( VREG_30_5 ) : ( n26305 ) ;
assign n26307 =  ( n25334 ) ? ( VREG_30_6 ) : ( n26306 ) ;
assign n26308 =  ( n25333 ) ? ( VREG_30_7 ) : ( n26307 ) ;
assign n26309 =  ( n25332 ) ? ( VREG_30_8 ) : ( n26308 ) ;
assign n26310 =  ( n25331 ) ? ( VREG_30_9 ) : ( n26309 ) ;
assign n26311 =  ( n25330 ) ? ( VREG_30_10 ) : ( n26310 ) ;
assign n26312 =  ( n25329 ) ? ( VREG_30_11 ) : ( n26311 ) ;
assign n26313 =  ( n25328 ) ? ( VREG_30_12 ) : ( n26312 ) ;
assign n26314 =  ( n25327 ) ? ( VREG_30_13 ) : ( n26313 ) ;
assign n26315 =  ( n25326 ) ? ( VREG_30_14 ) : ( n26314 ) ;
assign n26316 =  ( n25325 ) ? ( VREG_30_15 ) : ( n26315 ) ;
assign n26317 =  ( n25324 ) ? ( VREG_31_0 ) : ( n26316 ) ;
assign n26318 =  ( n25323 ) ? ( VREG_31_1 ) : ( n26317 ) ;
assign n26319 =  ( n25322 ) ? ( VREG_31_2 ) : ( n26318 ) ;
assign n26320 =  ( n25321 ) ? ( VREG_31_3 ) : ( n26319 ) ;
assign n26321 =  ( n25320 ) ? ( VREG_31_4 ) : ( n26320 ) ;
assign n26322 =  ( n25319 ) ? ( VREG_31_5 ) : ( n26321 ) ;
assign n26323 =  ( n25318 ) ? ( VREG_31_6 ) : ( n26322 ) ;
assign n26324 =  ( n25317 ) ? ( VREG_31_7 ) : ( n26323 ) ;
assign n26325 =  ( n25316 ) ? ( VREG_31_8 ) : ( n26324 ) ;
assign n26326 =  ( n25315 ) ? ( VREG_31_9 ) : ( n26325 ) ;
assign n26327 =  ( n25314 ) ? ( VREG_31_10 ) : ( n26326 ) ;
assign n26328 =  ( n25313 ) ? ( VREG_31_11 ) : ( n26327 ) ;
assign n26329 =  ( n25312 ) ? ( VREG_31_12 ) : ( n26328 ) ;
assign n26330 =  ( n25311 ) ? ( VREG_31_13 ) : ( n26329 ) ;
assign n26331 =  ( n25310 ) ? ( VREG_31_14 ) : ( n26330 ) ;
assign n26332 =  ( n25309 ) ? ( VREG_31_15 ) : ( n26331 ) ;
assign n26333 =  ( n25298 ) + ( n26332 )  ;
assign n26334 =  ( n25298 ) - ( n26332 )  ;
assign n26335 =  ( n25298 ) & ( n26332 )  ;
assign n26336 =  ( n25298 ) | ( n26332 )  ;
assign n26337 =  ( ( n25298 ) * ( n26332 ))  ;
assign n26338 =  ( n148 ) ? ( n26337 ) : ( VREG_0_5 ) ;
assign n26339 =  ( n146 ) ? ( n26336 ) : ( n26338 ) ;
assign n26340 =  ( n144 ) ? ( n26335 ) : ( n26339 ) ;
assign n26341 =  ( n142 ) ? ( n26334 ) : ( n26340 ) ;
assign n26342 =  ( n10 ) ? ( n26333 ) : ( n26341 ) ;
assign n26343 = n3030[5:5] ;
assign n26344 =  ( n26343 ) == ( 1'd0 )  ;
assign n26345 =  ( n26344 ) ? ( VREG_0_5 ) : ( n25308 ) ;
assign n26346 =  ( n26344 ) ? ( VREG_0_5 ) : ( n26342 ) ;
assign n26347 =  ( n3034 ) ? ( n26346 ) : ( VREG_0_5 ) ;
assign n26348 =  ( n2965 ) ? ( n26345 ) : ( n26347 ) ;
assign n26349 =  ( n1930 ) ? ( n26342 ) : ( n26348 ) ;
assign n26350 =  ( n879 ) ? ( n25308 ) : ( n26349 ) ;
assign n26351 =  ( n25298 ) + ( n164 )  ;
assign n26352 =  ( n25298 ) - ( n164 )  ;
assign n26353 =  ( n25298 ) & ( n164 )  ;
assign n26354 =  ( n25298 ) | ( n164 )  ;
assign n26355 =  ( ( n25298 ) * ( n164 ))  ;
assign n26356 =  ( n172 ) ? ( n26355 ) : ( VREG_0_5 ) ;
assign n26357 =  ( n170 ) ? ( n26354 ) : ( n26356 ) ;
assign n26358 =  ( n168 ) ? ( n26353 ) : ( n26357 ) ;
assign n26359 =  ( n166 ) ? ( n26352 ) : ( n26358 ) ;
assign n26360 =  ( n162 ) ? ( n26351 ) : ( n26359 ) ;
assign n26361 =  ( n25298 ) + ( n180 )  ;
assign n26362 =  ( n25298 ) - ( n180 )  ;
assign n26363 =  ( n25298 ) & ( n180 )  ;
assign n26364 =  ( n25298 ) | ( n180 )  ;
assign n26365 =  ( ( n25298 ) * ( n180 ))  ;
assign n26366 =  ( n172 ) ? ( n26365 ) : ( VREG_0_5 ) ;
assign n26367 =  ( n170 ) ? ( n26364 ) : ( n26366 ) ;
assign n26368 =  ( n168 ) ? ( n26363 ) : ( n26367 ) ;
assign n26369 =  ( n166 ) ? ( n26362 ) : ( n26368 ) ;
assign n26370 =  ( n162 ) ? ( n26361 ) : ( n26369 ) ;
assign n26371 =  ( n26344 ) ? ( VREG_0_5 ) : ( n26370 ) ;
assign n26372 =  ( n3051 ) ? ( n26371 ) : ( VREG_0_5 ) ;
assign n26373 =  ( n3040 ) ? ( n26360 ) : ( n26372 ) ;
assign n26374 =  ( n192 ) ? ( VREG_0_5 ) : ( VREG_0_5 ) ;
assign n26375 =  ( n157 ) ? ( n26373 ) : ( n26374 ) ;
assign n26376 =  ( n6 ) ? ( n26350 ) : ( n26375 ) ;
assign n26377 =  ( n4 ) ? ( n26376 ) : ( VREG_0_5 ) ;
assign n26378 =  ( 32'd6 ) == ( 32'd15 )  ;
assign n26379 =  ( n12 ) & ( n26378 )  ;
assign n26380 =  ( 32'd6 ) == ( 32'd14 )  ;
assign n26381 =  ( n12 ) & ( n26380 )  ;
assign n26382 =  ( 32'd6 ) == ( 32'd13 )  ;
assign n26383 =  ( n12 ) & ( n26382 )  ;
assign n26384 =  ( 32'd6 ) == ( 32'd12 )  ;
assign n26385 =  ( n12 ) & ( n26384 )  ;
assign n26386 =  ( 32'd6 ) == ( 32'd11 )  ;
assign n26387 =  ( n12 ) & ( n26386 )  ;
assign n26388 =  ( 32'd6 ) == ( 32'd10 )  ;
assign n26389 =  ( n12 ) & ( n26388 )  ;
assign n26390 =  ( 32'd6 ) == ( 32'd9 )  ;
assign n26391 =  ( n12 ) & ( n26390 )  ;
assign n26392 =  ( 32'd6 ) == ( 32'd8 )  ;
assign n26393 =  ( n12 ) & ( n26392 )  ;
assign n26394 =  ( 32'd6 ) == ( 32'd7 )  ;
assign n26395 =  ( n12 ) & ( n26394 )  ;
assign n26396 =  ( 32'd6 ) == ( 32'd6 )  ;
assign n26397 =  ( n12 ) & ( n26396 )  ;
assign n26398 =  ( 32'd6 ) == ( 32'd5 )  ;
assign n26399 =  ( n12 ) & ( n26398 )  ;
assign n26400 =  ( 32'd6 ) == ( 32'd4 )  ;
assign n26401 =  ( n12 ) & ( n26400 )  ;
assign n26402 =  ( 32'd6 ) == ( 32'd3 )  ;
assign n26403 =  ( n12 ) & ( n26402 )  ;
assign n26404 =  ( 32'd6 ) == ( 32'd2 )  ;
assign n26405 =  ( n12 ) & ( n26404 )  ;
assign n26406 =  ( 32'd6 ) == ( 32'd1 )  ;
assign n26407 =  ( n12 ) & ( n26406 )  ;
assign n26408 =  ( 32'd6 ) == ( 32'd0 )  ;
assign n26409 =  ( n12 ) & ( n26408 )  ;
assign n26410 =  ( n13 ) & ( n26378 )  ;
assign n26411 =  ( n13 ) & ( n26380 )  ;
assign n26412 =  ( n13 ) & ( n26382 )  ;
assign n26413 =  ( n13 ) & ( n26384 )  ;
assign n26414 =  ( n13 ) & ( n26386 )  ;
assign n26415 =  ( n13 ) & ( n26388 )  ;
assign n26416 =  ( n13 ) & ( n26390 )  ;
assign n26417 =  ( n13 ) & ( n26392 )  ;
assign n26418 =  ( n13 ) & ( n26394 )  ;
assign n26419 =  ( n13 ) & ( n26396 )  ;
assign n26420 =  ( n13 ) & ( n26398 )  ;
assign n26421 =  ( n13 ) & ( n26400 )  ;
assign n26422 =  ( n13 ) & ( n26402 )  ;
assign n26423 =  ( n13 ) & ( n26404 )  ;
assign n26424 =  ( n13 ) & ( n26406 )  ;
assign n26425 =  ( n13 ) & ( n26408 )  ;
assign n26426 =  ( n14 ) & ( n26378 )  ;
assign n26427 =  ( n14 ) & ( n26380 )  ;
assign n26428 =  ( n14 ) & ( n26382 )  ;
assign n26429 =  ( n14 ) & ( n26384 )  ;
assign n26430 =  ( n14 ) & ( n26386 )  ;
assign n26431 =  ( n14 ) & ( n26388 )  ;
assign n26432 =  ( n14 ) & ( n26390 )  ;
assign n26433 =  ( n14 ) & ( n26392 )  ;
assign n26434 =  ( n14 ) & ( n26394 )  ;
assign n26435 =  ( n14 ) & ( n26396 )  ;
assign n26436 =  ( n14 ) & ( n26398 )  ;
assign n26437 =  ( n14 ) & ( n26400 )  ;
assign n26438 =  ( n14 ) & ( n26402 )  ;
assign n26439 =  ( n14 ) & ( n26404 )  ;
assign n26440 =  ( n14 ) & ( n26406 )  ;
assign n26441 =  ( n14 ) & ( n26408 )  ;
assign n26442 =  ( n15 ) & ( n26378 )  ;
assign n26443 =  ( n15 ) & ( n26380 )  ;
assign n26444 =  ( n15 ) & ( n26382 )  ;
assign n26445 =  ( n15 ) & ( n26384 )  ;
assign n26446 =  ( n15 ) & ( n26386 )  ;
assign n26447 =  ( n15 ) & ( n26388 )  ;
assign n26448 =  ( n15 ) & ( n26390 )  ;
assign n26449 =  ( n15 ) & ( n26392 )  ;
assign n26450 =  ( n15 ) & ( n26394 )  ;
assign n26451 =  ( n15 ) & ( n26396 )  ;
assign n26452 =  ( n15 ) & ( n26398 )  ;
assign n26453 =  ( n15 ) & ( n26400 )  ;
assign n26454 =  ( n15 ) & ( n26402 )  ;
assign n26455 =  ( n15 ) & ( n26404 )  ;
assign n26456 =  ( n15 ) & ( n26406 )  ;
assign n26457 =  ( n15 ) & ( n26408 )  ;
assign n26458 =  ( n16 ) & ( n26378 )  ;
assign n26459 =  ( n16 ) & ( n26380 )  ;
assign n26460 =  ( n16 ) & ( n26382 )  ;
assign n26461 =  ( n16 ) & ( n26384 )  ;
assign n26462 =  ( n16 ) & ( n26386 )  ;
assign n26463 =  ( n16 ) & ( n26388 )  ;
assign n26464 =  ( n16 ) & ( n26390 )  ;
assign n26465 =  ( n16 ) & ( n26392 )  ;
assign n26466 =  ( n16 ) & ( n26394 )  ;
assign n26467 =  ( n16 ) & ( n26396 )  ;
assign n26468 =  ( n16 ) & ( n26398 )  ;
assign n26469 =  ( n16 ) & ( n26400 )  ;
assign n26470 =  ( n16 ) & ( n26402 )  ;
assign n26471 =  ( n16 ) & ( n26404 )  ;
assign n26472 =  ( n16 ) & ( n26406 )  ;
assign n26473 =  ( n16 ) & ( n26408 )  ;
assign n26474 =  ( n17 ) & ( n26378 )  ;
assign n26475 =  ( n17 ) & ( n26380 )  ;
assign n26476 =  ( n17 ) & ( n26382 )  ;
assign n26477 =  ( n17 ) & ( n26384 )  ;
assign n26478 =  ( n17 ) & ( n26386 )  ;
assign n26479 =  ( n17 ) & ( n26388 )  ;
assign n26480 =  ( n17 ) & ( n26390 )  ;
assign n26481 =  ( n17 ) & ( n26392 )  ;
assign n26482 =  ( n17 ) & ( n26394 )  ;
assign n26483 =  ( n17 ) & ( n26396 )  ;
assign n26484 =  ( n17 ) & ( n26398 )  ;
assign n26485 =  ( n17 ) & ( n26400 )  ;
assign n26486 =  ( n17 ) & ( n26402 )  ;
assign n26487 =  ( n17 ) & ( n26404 )  ;
assign n26488 =  ( n17 ) & ( n26406 )  ;
assign n26489 =  ( n17 ) & ( n26408 )  ;
assign n26490 =  ( n18 ) & ( n26378 )  ;
assign n26491 =  ( n18 ) & ( n26380 )  ;
assign n26492 =  ( n18 ) & ( n26382 )  ;
assign n26493 =  ( n18 ) & ( n26384 )  ;
assign n26494 =  ( n18 ) & ( n26386 )  ;
assign n26495 =  ( n18 ) & ( n26388 )  ;
assign n26496 =  ( n18 ) & ( n26390 )  ;
assign n26497 =  ( n18 ) & ( n26392 )  ;
assign n26498 =  ( n18 ) & ( n26394 )  ;
assign n26499 =  ( n18 ) & ( n26396 )  ;
assign n26500 =  ( n18 ) & ( n26398 )  ;
assign n26501 =  ( n18 ) & ( n26400 )  ;
assign n26502 =  ( n18 ) & ( n26402 )  ;
assign n26503 =  ( n18 ) & ( n26404 )  ;
assign n26504 =  ( n18 ) & ( n26406 )  ;
assign n26505 =  ( n18 ) & ( n26408 )  ;
assign n26506 =  ( n19 ) & ( n26378 )  ;
assign n26507 =  ( n19 ) & ( n26380 )  ;
assign n26508 =  ( n19 ) & ( n26382 )  ;
assign n26509 =  ( n19 ) & ( n26384 )  ;
assign n26510 =  ( n19 ) & ( n26386 )  ;
assign n26511 =  ( n19 ) & ( n26388 )  ;
assign n26512 =  ( n19 ) & ( n26390 )  ;
assign n26513 =  ( n19 ) & ( n26392 )  ;
assign n26514 =  ( n19 ) & ( n26394 )  ;
assign n26515 =  ( n19 ) & ( n26396 )  ;
assign n26516 =  ( n19 ) & ( n26398 )  ;
assign n26517 =  ( n19 ) & ( n26400 )  ;
assign n26518 =  ( n19 ) & ( n26402 )  ;
assign n26519 =  ( n19 ) & ( n26404 )  ;
assign n26520 =  ( n19 ) & ( n26406 )  ;
assign n26521 =  ( n19 ) & ( n26408 )  ;
assign n26522 =  ( n20 ) & ( n26378 )  ;
assign n26523 =  ( n20 ) & ( n26380 )  ;
assign n26524 =  ( n20 ) & ( n26382 )  ;
assign n26525 =  ( n20 ) & ( n26384 )  ;
assign n26526 =  ( n20 ) & ( n26386 )  ;
assign n26527 =  ( n20 ) & ( n26388 )  ;
assign n26528 =  ( n20 ) & ( n26390 )  ;
assign n26529 =  ( n20 ) & ( n26392 )  ;
assign n26530 =  ( n20 ) & ( n26394 )  ;
assign n26531 =  ( n20 ) & ( n26396 )  ;
assign n26532 =  ( n20 ) & ( n26398 )  ;
assign n26533 =  ( n20 ) & ( n26400 )  ;
assign n26534 =  ( n20 ) & ( n26402 )  ;
assign n26535 =  ( n20 ) & ( n26404 )  ;
assign n26536 =  ( n20 ) & ( n26406 )  ;
assign n26537 =  ( n20 ) & ( n26408 )  ;
assign n26538 =  ( n21 ) & ( n26378 )  ;
assign n26539 =  ( n21 ) & ( n26380 )  ;
assign n26540 =  ( n21 ) & ( n26382 )  ;
assign n26541 =  ( n21 ) & ( n26384 )  ;
assign n26542 =  ( n21 ) & ( n26386 )  ;
assign n26543 =  ( n21 ) & ( n26388 )  ;
assign n26544 =  ( n21 ) & ( n26390 )  ;
assign n26545 =  ( n21 ) & ( n26392 )  ;
assign n26546 =  ( n21 ) & ( n26394 )  ;
assign n26547 =  ( n21 ) & ( n26396 )  ;
assign n26548 =  ( n21 ) & ( n26398 )  ;
assign n26549 =  ( n21 ) & ( n26400 )  ;
assign n26550 =  ( n21 ) & ( n26402 )  ;
assign n26551 =  ( n21 ) & ( n26404 )  ;
assign n26552 =  ( n21 ) & ( n26406 )  ;
assign n26553 =  ( n21 ) & ( n26408 )  ;
assign n26554 =  ( n22 ) & ( n26378 )  ;
assign n26555 =  ( n22 ) & ( n26380 )  ;
assign n26556 =  ( n22 ) & ( n26382 )  ;
assign n26557 =  ( n22 ) & ( n26384 )  ;
assign n26558 =  ( n22 ) & ( n26386 )  ;
assign n26559 =  ( n22 ) & ( n26388 )  ;
assign n26560 =  ( n22 ) & ( n26390 )  ;
assign n26561 =  ( n22 ) & ( n26392 )  ;
assign n26562 =  ( n22 ) & ( n26394 )  ;
assign n26563 =  ( n22 ) & ( n26396 )  ;
assign n26564 =  ( n22 ) & ( n26398 )  ;
assign n26565 =  ( n22 ) & ( n26400 )  ;
assign n26566 =  ( n22 ) & ( n26402 )  ;
assign n26567 =  ( n22 ) & ( n26404 )  ;
assign n26568 =  ( n22 ) & ( n26406 )  ;
assign n26569 =  ( n22 ) & ( n26408 )  ;
assign n26570 =  ( n23 ) & ( n26378 )  ;
assign n26571 =  ( n23 ) & ( n26380 )  ;
assign n26572 =  ( n23 ) & ( n26382 )  ;
assign n26573 =  ( n23 ) & ( n26384 )  ;
assign n26574 =  ( n23 ) & ( n26386 )  ;
assign n26575 =  ( n23 ) & ( n26388 )  ;
assign n26576 =  ( n23 ) & ( n26390 )  ;
assign n26577 =  ( n23 ) & ( n26392 )  ;
assign n26578 =  ( n23 ) & ( n26394 )  ;
assign n26579 =  ( n23 ) & ( n26396 )  ;
assign n26580 =  ( n23 ) & ( n26398 )  ;
assign n26581 =  ( n23 ) & ( n26400 )  ;
assign n26582 =  ( n23 ) & ( n26402 )  ;
assign n26583 =  ( n23 ) & ( n26404 )  ;
assign n26584 =  ( n23 ) & ( n26406 )  ;
assign n26585 =  ( n23 ) & ( n26408 )  ;
assign n26586 =  ( n24 ) & ( n26378 )  ;
assign n26587 =  ( n24 ) & ( n26380 )  ;
assign n26588 =  ( n24 ) & ( n26382 )  ;
assign n26589 =  ( n24 ) & ( n26384 )  ;
assign n26590 =  ( n24 ) & ( n26386 )  ;
assign n26591 =  ( n24 ) & ( n26388 )  ;
assign n26592 =  ( n24 ) & ( n26390 )  ;
assign n26593 =  ( n24 ) & ( n26392 )  ;
assign n26594 =  ( n24 ) & ( n26394 )  ;
assign n26595 =  ( n24 ) & ( n26396 )  ;
assign n26596 =  ( n24 ) & ( n26398 )  ;
assign n26597 =  ( n24 ) & ( n26400 )  ;
assign n26598 =  ( n24 ) & ( n26402 )  ;
assign n26599 =  ( n24 ) & ( n26404 )  ;
assign n26600 =  ( n24 ) & ( n26406 )  ;
assign n26601 =  ( n24 ) & ( n26408 )  ;
assign n26602 =  ( n25 ) & ( n26378 )  ;
assign n26603 =  ( n25 ) & ( n26380 )  ;
assign n26604 =  ( n25 ) & ( n26382 )  ;
assign n26605 =  ( n25 ) & ( n26384 )  ;
assign n26606 =  ( n25 ) & ( n26386 )  ;
assign n26607 =  ( n25 ) & ( n26388 )  ;
assign n26608 =  ( n25 ) & ( n26390 )  ;
assign n26609 =  ( n25 ) & ( n26392 )  ;
assign n26610 =  ( n25 ) & ( n26394 )  ;
assign n26611 =  ( n25 ) & ( n26396 )  ;
assign n26612 =  ( n25 ) & ( n26398 )  ;
assign n26613 =  ( n25 ) & ( n26400 )  ;
assign n26614 =  ( n25 ) & ( n26402 )  ;
assign n26615 =  ( n25 ) & ( n26404 )  ;
assign n26616 =  ( n25 ) & ( n26406 )  ;
assign n26617 =  ( n25 ) & ( n26408 )  ;
assign n26618 =  ( n26 ) & ( n26378 )  ;
assign n26619 =  ( n26 ) & ( n26380 )  ;
assign n26620 =  ( n26 ) & ( n26382 )  ;
assign n26621 =  ( n26 ) & ( n26384 )  ;
assign n26622 =  ( n26 ) & ( n26386 )  ;
assign n26623 =  ( n26 ) & ( n26388 )  ;
assign n26624 =  ( n26 ) & ( n26390 )  ;
assign n26625 =  ( n26 ) & ( n26392 )  ;
assign n26626 =  ( n26 ) & ( n26394 )  ;
assign n26627 =  ( n26 ) & ( n26396 )  ;
assign n26628 =  ( n26 ) & ( n26398 )  ;
assign n26629 =  ( n26 ) & ( n26400 )  ;
assign n26630 =  ( n26 ) & ( n26402 )  ;
assign n26631 =  ( n26 ) & ( n26404 )  ;
assign n26632 =  ( n26 ) & ( n26406 )  ;
assign n26633 =  ( n26 ) & ( n26408 )  ;
assign n26634 =  ( n27 ) & ( n26378 )  ;
assign n26635 =  ( n27 ) & ( n26380 )  ;
assign n26636 =  ( n27 ) & ( n26382 )  ;
assign n26637 =  ( n27 ) & ( n26384 )  ;
assign n26638 =  ( n27 ) & ( n26386 )  ;
assign n26639 =  ( n27 ) & ( n26388 )  ;
assign n26640 =  ( n27 ) & ( n26390 )  ;
assign n26641 =  ( n27 ) & ( n26392 )  ;
assign n26642 =  ( n27 ) & ( n26394 )  ;
assign n26643 =  ( n27 ) & ( n26396 )  ;
assign n26644 =  ( n27 ) & ( n26398 )  ;
assign n26645 =  ( n27 ) & ( n26400 )  ;
assign n26646 =  ( n27 ) & ( n26402 )  ;
assign n26647 =  ( n27 ) & ( n26404 )  ;
assign n26648 =  ( n27 ) & ( n26406 )  ;
assign n26649 =  ( n27 ) & ( n26408 )  ;
assign n26650 =  ( n28 ) & ( n26378 )  ;
assign n26651 =  ( n28 ) & ( n26380 )  ;
assign n26652 =  ( n28 ) & ( n26382 )  ;
assign n26653 =  ( n28 ) & ( n26384 )  ;
assign n26654 =  ( n28 ) & ( n26386 )  ;
assign n26655 =  ( n28 ) & ( n26388 )  ;
assign n26656 =  ( n28 ) & ( n26390 )  ;
assign n26657 =  ( n28 ) & ( n26392 )  ;
assign n26658 =  ( n28 ) & ( n26394 )  ;
assign n26659 =  ( n28 ) & ( n26396 )  ;
assign n26660 =  ( n28 ) & ( n26398 )  ;
assign n26661 =  ( n28 ) & ( n26400 )  ;
assign n26662 =  ( n28 ) & ( n26402 )  ;
assign n26663 =  ( n28 ) & ( n26404 )  ;
assign n26664 =  ( n28 ) & ( n26406 )  ;
assign n26665 =  ( n28 ) & ( n26408 )  ;
assign n26666 =  ( n29 ) & ( n26378 )  ;
assign n26667 =  ( n29 ) & ( n26380 )  ;
assign n26668 =  ( n29 ) & ( n26382 )  ;
assign n26669 =  ( n29 ) & ( n26384 )  ;
assign n26670 =  ( n29 ) & ( n26386 )  ;
assign n26671 =  ( n29 ) & ( n26388 )  ;
assign n26672 =  ( n29 ) & ( n26390 )  ;
assign n26673 =  ( n29 ) & ( n26392 )  ;
assign n26674 =  ( n29 ) & ( n26394 )  ;
assign n26675 =  ( n29 ) & ( n26396 )  ;
assign n26676 =  ( n29 ) & ( n26398 )  ;
assign n26677 =  ( n29 ) & ( n26400 )  ;
assign n26678 =  ( n29 ) & ( n26402 )  ;
assign n26679 =  ( n29 ) & ( n26404 )  ;
assign n26680 =  ( n29 ) & ( n26406 )  ;
assign n26681 =  ( n29 ) & ( n26408 )  ;
assign n26682 =  ( n30 ) & ( n26378 )  ;
assign n26683 =  ( n30 ) & ( n26380 )  ;
assign n26684 =  ( n30 ) & ( n26382 )  ;
assign n26685 =  ( n30 ) & ( n26384 )  ;
assign n26686 =  ( n30 ) & ( n26386 )  ;
assign n26687 =  ( n30 ) & ( n26388 )  ;
assign n26688 =  ( n30 ) & ( n26390 )  ;
assign n26689 =  ( n30 ) & ( n26392 )  ;
assign n26690 =  ( n30 ) & ( n26394 )  ;
assign n26691 =  ( n30 ) & ( n26396 )  ;
assign n26692 =  ( n30 ) & ( n26398 )  ;
assign n26693 =  ( n30 ) & ( n26400 )  ;
assign n26694 =  ( n30 ) & ( n26402 )  ;
assign n26695 =  ( n30 ) & ( n26404 )  ;
assign n26696 =  ( n30 ) & ( n26406 )  ;
assign n26697 =  ( n30 ) & ( n26408 )  ;
assign n26698 =  ( n31 ) & ( n26378 )  ;
assign n26699 =  ( n31 ) & ( n26380 )  ;
assign n26700 =  ( n31 ) & ( n26382 )  ;
assign n26701 =  ( n31 ) & ( n26384 )  ;
assign n26702 =  ( n31 ) & ( n26386 )  ;
assign n26703 =  ( n31 ) & ( n26388 )  ;
assign n26704 =  ( n31 ) & ( n26390 )  ;
assign n26705 =  ( n31 ) & ( n26392 )  ;
assign n26706 =  ( n31 ) & ( n26394 )  ;
assign n26707 =  ( n31 ) & ( n26396 )  ;
assign n26708 =  ( n31 ) & ( n26398 )  ;
assign n26709 =  ( n31 ) & ( n26400 )  ;
assign n26710 =  ( n31 ) & ( n26402 )  ;
assign n26711 =  ( n31 ) & ( n26404 )  ;
assign n26712 =  ( n31 ) & ( n26406 )  ;
assign n26713 =  ( n31 ) & ( n26408 )  ;
assign n26714 =  ( n32 ) & ( n26378 )  ;
assign n26715 =  ( n32 ) & ( n26380 )  ;
assign n26716 =  ( n32 ) & ( n26382 )  ;
assign n26717 =  ( n32 ) & ( n26384 )  ;
assign n26718 =  ( n32 ) & ( n26386 )  ;
assign n26719 =  ( n32 ) & ( n26388 )  ;
assign n26720 =  ( n32 ) & ( n26390 )  ;
assign n26721 =  ( n32 ) & ( n26392 )  ;
assign n26722 =  ( n32 ) & ( n26394 )  ;
assign n26723 =  ( n32 ) & ( n26396 )  ;
assign n26724 =  ( n32 ) & ( n26398 )  ;
assign n26725 =  ( n32 ) & ( n26400 )  ;
assign n26726 =  ( n32 ) & ( n26402 )  ;
assign n26727 =  ( n32 ) & ( n26404 )  ;
assign n26728 =  ( n32 ) & ( n26406 )  ;
assign n26729 =  ( n32 ) & ( n26408 )  ;
assign n26730 =  ( n33 ) & ( n26378 )  ;
assign n26731 =  ( n33 ) & ( n26380 )  ;
assign n26732 =  ( n33 ) & ( n26382 )  ;
assign n26733 =  ( n33 ) & ( n26384 )  ;
assign n26734 =  ( n33 ) & ( n26386 )  ;
assign n26735 =  ( n33 ) & ( n26388 )  ;
assign n26736 =  ( n33 ) & ( n26390 )  ;
assign n26737 =  ( n33 ) & ( n26392 )  ;
assign n26738 =  ( n33 ) & ( n26394 )  ;
assign n26739 =  ( n33 ) & ( n26396 )  ;
assign n26740 =  ( n33 ) & ( n26398 )  ;
assign n26741 =  ( n33 ) & ( n26400 )  ;
assign n26742 =  ( n33 ) & ( n26402 )  ;
assign n26743 =  ( n33 ) & ( n26404 )  ;
assign n26744 =  ( n33 ) & ( n26406 )  ;
assign n26745 =  ( n33 ) & ( n26408 )  ;
assign n26746 =  ( n34 ) & ( n26378 )  ;
assign n26747 =  ( n34 ) & ( n26380 )  ;
assign n26748 =  ( n34 ) & ( n26382 )  ;
assign n26749 =  ( n34 ) & ( n26384 )  ;
assign n26750 =  ( n34 ) & ( n26386 )  ;
assign n26751 =  ( n34 ) & ( n26388 )  ;
assign n26752 =  ( n34 ) & ( n26390 )  ;
assign n26753 =  ( n34 ) & ( n26392 )  ;
assign n26754 =  ( n34 ) & ( n26394 )  ;
assign n26755 =  ( n34 ) & ( n26396 )  ;
assign n26756 =  ( n34 ) & ( n26398 )  ;
assign n26757 =  ( n34 ) & ( n26400 )  ;
assign n26758 =  ( n34 ) & ( n26402 )  ;
assign n26759 =  ( n34 ) & ( n26404 )  ;
assign n26760 =  ( n34 ) & ( n26406 )  ;
assign n26761 =  ( n34 ) & ( n26408 )  ;
assign n26762 =  ( n35 ) & ( n26378 )  ;
assign n26763 =  ( n35 ) & ( n26380 )  ;
assign n26764 =  ( n35 ) & ( n26382 )  ;
assign n26765 =  ( n35 ) & ( n26384 )  ;
assign n26766 =  ( n35 ) & ( n26386 )  ;
assign n26767 =  ( n35 ) & ( n26388 )  ;
assign n26768 =  ( n35 ) & ( n26390 )  ;
assign n26769 =  ( n35 ) & ( n26392 )  ;
assign n26770 =  ( n35 ) & ( n26394 )  ;
assign n26771 =  ( n35 ) & ( n26396 )  ;
assign n26772 =  ( n35 ) & ( n26398 )  ;
assign n26773 =  ( n35 ) & ( n26400 )  ;
assign n26774 =  ( n35 ) & ( n26402 )  ;
assign n26775 =  ( n35 ) & ( n26404 )  ;
assign n26776 =  ( n35 ) & ( n26406 )  ;
assign n26777 =  ( n35 ) & ( n26408 )  ;
assign n26778 =  ( n36 ) & ( n26378 )  ;
assign n26779 =  ( n36 ) & ( n26380 )  ;
assign n26780 =  ( n36 ) & ( n26382 )  ;
assign n26781 =  ( n36 ) & ( n26384 )  ;
assign n26782 =  ( n36 ) & ( n26386 )  ;
assign n26783 =  ( n36 ) & ( n26388 )  ;
assign n26784 =  ( n36 ) & ( n26390 )  ;
assign n26785 =  ( n36 ) & ( n26392 )  ;
assign n26786 =  ( n36 ) & ( n26394 )  ;
assign n26787 =  ( n36 ) & ( n26396 )  ;
assign n26788 =  ( n36 ) & ( n26398 )  ;
assign n26789 =  ( n36 ) & ( n26400 )  ;
assign n26790 =  ( n36 ) & ( n26402 )  ;
assign n26791 =  ( n36 ) & ( n26404 )  ;
assign n26792 =  ( n36 ) & ( n26406 )  ;
assign n26793 =  ( n36 ) & ( n26408 )  ;
assign n26794 =  ( n37 ) & ( n26378 )  ;
assign n26795 =  ( n37 ) & ( n26380 )  ;
assign n26796 =  ( n37 ) & ( n26382 )  ;
assign n26797 =  ( n37 ) & ( n26384 )  ;
assign n26798 =  ( n37 ) & ( n26386 )  ;
assign n26799 =  ( n37 ) & ( n26388 )  ;
assign n26800 =  ( n37 ) & ( n26390 )  ;
assign n26801 =  ( n37 ) & ( n26392 )  ;
assign n26802 =  ( n37 ) & ( n26394 )  ;
assign n26803 =  ( n37 ) & ( n26396 )  ;
assign n26804 =  ( n37 ) & ( n26398 )  ;
assign n26805 =  ( n37 ) & ( n26400 )  ;
assign n26806 =  ( n37 ) & ( n26402 )  ;
assign n26807 =  ( n37 ) & ( n26404 )  ;
assign n26808 =  ( n37 ) & ( n26406 )  ;
assign n26809 =  ( n37 ) & ( n26408 )  ;
assign n26810 =  ( n38 ) & ( n26378 )  ;
assign n26811 =  ( n38 ) & ( n26380 )  ;
assign n26812 =  ( n38 ) & ( n26382 )  ;
assign n26813 =  ( n38 ) & ( n26384 )  ;
assign n26814 =  ( n38 ) & ( n26386 )  ;
assign n26815 =  ( n38 ) & ( n26388 )  ;
assign n26816 =  ( n38 ) & ( n26390 )  ;
assign n26817 =  ( n38 ) & ( n26392 )  ;
assign n26818 =  ( n38 ) & ( n26394 )  ;
assign n26819 =  ( n38 ) & ( n26396 )  ;
assign n26820 =  ( n38 ) & ( n26398 )  ;
assign n26821 =  ( n38 ) & ( n26400 )  ;
assign n26822 =  ( n38 ) & ( n26402 )  ;
assign n26823 =  ( n38 ) & ( n26404 )  ;
assign n26824 =  ( n38 ) & ( n26406 )  ;
assign n26825 =  ( n38 ) & ( n26408 )  ;
assign n26826 =  ( n39 ) & ( n26378 )  ;
assign n26827 =  ( n39 ) & ( n26380 )  ;
assign n26828 =  ( n39 ) & ( n26382 )  ;
assign n26829 =  ( n39 ) & ( n26384 )  ;
assign n26830 =  ( n39 ) & ( n26386 )  ;
assign n26831 =  ( n39 ) & ( n26388 )  ;
assign n26832 =  ( n39 ) & ( n26390 )  ;
assign n26833 =  ( n39 ) & ( n26392 )  ;
assign n26834 =  ( n39 ) & ( n26394 )  ;
assign n26835 =  ( n39 ) & ( n26396 )  ;
assign n26836 =  ( n39 ) & ( n26398 )  ;
assign n26837 =  ( n39 ) & ( n26400 )  ;
assign n26838 =  ( n39 ) & ( n26402 )  ;
assign n26839 =  ( n39 ) & ( n26404 )  ;
assign n26840 =  ( n39 ) & ( n26406 )  ;
assign n26841 =  ( n39 ) & ( n26408 )  ;
assign n26842 =  ( n40 ) & ( n26378 )  ;
assign n26843 =  ( n40 ) & ( n26380 )  ;
assign n26844 =  ( n40 ) & ( n26382 )  ;
assign n26845 =  ( n40 ) & ( n26384 )  ;
assign n26846 =  ( n40 ) & ( n26386 )  ;
assign n26847 =  ( n40 ) & ( n26388 )  ;
assign n26848 =  ( n40 ) & ( n26390 )  ;
assign n26849 =  ( n40 ) & ( n26392 )  ;
assign n26850 =  ( n40 ) & ( n26394 )  ;
assign n26851 =  ( n40 ) & ( n26396 )  ;
assign n26852 =  ( n40 ) & ( n26398 )  ;
assign n26853 =  ( n40 ) & ( n26400 )  ;
assign n26854 =  ( n40 ) & ( n26402 )  ;
assign n26855 =  ( n40 ) & ( n26404 )  ;
assign n26856 =  ( n40 ) & ( n26406 )  ;
assign n26857 =  ( n40 ) & ( n26408 )  ;
assign n26858 =  ( n41 ) & ( n26378 )  ;
assign n26859 =  ( n41 ) & ( n26380 )  ;
assign n26860 =  ( n41 ) & ( n26382 )  ;
assign n26861 =  ( n41 ) & ( n26384 )  ;
assign n26862 =  ( n41 ) & ( n26386 )  ;
assign n26863 =  ( n41 ) & ( n26388 )  ;
assign n26864 =  ( n41 ) & ( n26390 )  ;
assign n26865 =  ( n41 ) & ( n26392 )  ;
assign n26866 =  ( n41 ) & ( n26394 )  ;
assign n26867 =  ( n41 ) & ( n26396 )  ;
assign n26868 =  ( n41 ) & ( n26398 )  ;
assign n26869 =  ( n41 ) & ( n26400 )  ;
assign n26870 =  ( n41 ) & ( n26402 )  ;
assign n26871 =  ( n41 ) & ( n26404 )  ;
assign n26872 =  ( n41 ) & ( n26406 )  ;
assign n26873 =  ( n41 ) & ( n26408 )  ;
assign n26874 =  ( n42 ) & ( n26378 )  ;
assign n26875 =  ( n42 ) & ( n26380 )  ;
assign n26876 =  ( n42 ) & ( n26382 )  ;
assign n26877 =  ( n42 ) & ( n26384 )  ;
assign n26878 =  ( n42 ) & ( n26386 )  ;
assign n26879 =  ( n42 ) & ( n26388 )  ;
assign n26880 =  ( n42 ) & ( n26390 )  ;
assign n26881 =  ( n42 ) & ( n26392 )  ;
assign n26882 =  ( n42 ) & ( n26394 )  ;
assign n26883 =  ( n42 ) & ( n26396 )  ;
assign n26884 =  ( n42 ) & ( n26398 )  ;
assign n26885 =  ( n42 ) & ( n26400 )  ;
assign n26886 =  ( n42 ) & ( n26402 )  ;
assign n26887 =  ( n42 ) & ( n26404 )  ;
assign n26888 =  ( n42 ) & ( n26406 )  ;
assign n26889 =  ( n42 ) & ( n26408 )  ;
assign n26890 =  ( n43 ) & ( n26378 )  ;
assign n26891 =  ( n43 ) & ( n26380 )  ;
assign n26892 =  ( n43 ) & ( n26382 )  ;
assign n26893 =  ( n43 ) & ( n26384 )  ;
assign n26894 =  ( n43 ) & ( n26386 )  ;
assign n26895 =  ( n43 ) & ( n26388 )  ;
assign n26896 =  ( n43 ) & ( n26390 )  ;
assign n26897 =  ( n43 ) & ( n26392 )  ;
assign n26898 =  ( n43 ) & ( n26394 )  ;
assign n26899 =  ( n43 ) & ( n26396 )  ;
assign n26900 =  ( n43 ) & ( n26398 )  ;
assign n26901 =  ( n43 ) & ( n26400 )  ;
assign n26902 =  ( n43 ) & ( n26402 )  ;
assign n26903 =  ( n43 ) & ( n26404 )  ;
assign n26904 =  ( n43 ) & ( n26406 )  ;
assign n26905 =  ( n43 ) & ( n26408 )  ;
assign n26906 =  ( n26905 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n26907 =  ( n26904 ) ? ( VREG_0_1 ) : ( n26906 ) ;
assign n26908 =  ( n26903 ) ? ( VREG_0_2 ) : ( n26907 ) ;
assign n26909 =  ( n26902 ) ? ( VREG_0_3 ) : ( n26908 ) ;
assign n26910 =  ( n26901 ) ? ( VREG_0_4 ) : ( n26909 ) ;
assign n26911 =  ( n26900 ) ? ( VREG_0_5 ) : ( n26910 ) ;
assign n26912 =  ( n26899 ) ? ( VREG_0_6 ) : ( n26911 ) ;
assign n26913 =  ( n26898 ) ? ( VREG_0_7 ) : ( n26912 ) ;
assign n26914 =  ( n26897 ) ? ( VREG_0_8 ) : ( n26913 ) ;
assign n26915 =  ( n26896 ) ? ( VREG_0_9 ) : ( n26914 ) ;
assign n26916 =  ( n26895 ) ? ( VREG_0_10 ) : ( n26915 ) ;
assign n26917 =  ( n26894 ) ? ( VREG_0_11 ) : ( n26916 ) ;
assign n26918 =  ( n26893 ) ? ( VREG_0_12 ) : ( n26917 ) ;
assign n26919 =  ( n26892 ) ? ( VREG_0_13 ) : ( n26918 ) ;
assign n26920 =  ( n26891 ) ? ( VREG_0_14 ) : ( n26919 ) ;
assign n26921 =  ( n26890 ) ? ( VREG_0_15 ) : ( n26920 ) ;
assign n26922 =  ( n26889 ) ? ( VREG_1_0 ) : ( n26921 ) ;
assign n26923 =  ( n26888 ) ? ( VREG_1_1 ) : ( n26922 ) ;
assign n26924 =  ( n26887 ) ? ( VREG_1_2 ) : ( n26923 ) ;
assign n26925 =  ( n26886 ) ? ( VREG_1_3 ) : ( n26924 ) ;
assign n26926 =  ( n26885 ) ? ( VREG_1_4 ) : ( n26925 ) ;
assign n26927 =  ( n26884 ) ? ( VREG_1_5 ) : ( n26926 ) ;
assign n26928 =  ( n26883 ) ? ( VREG_1_6 ) : ( n26927 ) ;
assign n26929 =  ( n26882 ) ? ( VREG_1_7 ) : ( n26928 ) ;
assign n26930 =  ( n26881 ) ? ( VREG_1_8 ) : ( n26929 ) ;
assign n26931 =  ( n26880 ) ? ( VREG_1_9 ) : ( n26930 ) ;
assign n26932 =  ( n26879 ) ? ( VREG_1_10 ) : ( n26931 ) ;
assign n26933 =  ( n26878 ) ? ( VREG_1_11 ) : ( n26932 ) ;
assign n26934 =  ( n26877 ) ? ( VREG_1_12 ) : ( n26933 ) ;
assign n26935 =  ( n26876 ) ? ( VREG_1_13 ) : ( n26934 ) ;
assign n26936 =  ( n26875 ) ? ( VREG_1_14 ) : ( n26935 ) ;
assign n26937 =  ( n26874 ) ? ( VREG_1_15 ) : ( n26936 ) ;
assign n26938 =  ( n26873 ) ? ( VREG_2_0 ) : ( n26937 ) ;
assign n26939 =  ( n26872 ) ? ( VREG_2_1 ) : ( n26938 ) ;
assign n26940 =  ( n26871 ) ? ( VREG_2_2 ) : ( n26939 ) ;
assign n26941 =  ( n26870 ) ? ( VREG_2_3 ) : ( n26940 ) ;
assign n26942 =  ( n26869 ) ? ( VREG_2_4 ) : ( n26941 ) ;
assign n26943 =  ( n26868 ) ? ( VREG_2_5 ) : ( n26942 ) ;
assign n26944 =  ( n26867 ) ? ( VREG_2_6 ) : ( n26943 ) ;
assign n26945 =  ( n26866 ) ? ( VREG_2_7 ) : ( n26944 ) ;
assign n26946 =  ( n26865 ) ? ( VREG_2_8 ) : ( n26945 ) ;
assign n26947 =  ( n26864 ) ? ( VREG_2_9 ) : ( n26946 ) ;
assign n26948 =  ( n26863 ) ? ( VREG_2_10 ) : ( n26947 ) ;
assign n26949 =  ( n26862 ) ? ( VREG_2_11 ) : ( n26948 ) ;
assign n26950 =  ( n26861 ) ? ( VREG_2_12 ) : ( n26949 ) ;
assign n26951 =  ( n26860 ) ? ( VREG_2_13 ) : ( n26950 ) ;
assign n26952 =  ( n26859 ) ? ( VREG_2_14 ) : ( n26951 ) ;
assign n26953 =  ( n26858 ) ? ( VREG_2_15 ) : ( n26952 ) ;
assign n26954 =  ( n26857 ) ? ( VREG_3_0 ) : ( n26953 ) ;
assign n26955 =  ( n26856 ) ? ( VREG_3_1 ) : ( n26954 ) ;
assign n26956 =  ( n26855 ) ? ( VREG_3_2 ) : ( n26955 ) ;
assign n26957 =  ( n26854 ) ? ( VREG_3_3 ) : ( n26956 ) ;
assign n26958 =  ( n26853 ) ? ( VREG_3_4 ) : ( n26957 ) ;
assign n26959 =  ( n26852 ) ? ( VREG_3_5 ) : ( n26958 ) ;
assign n26960 =  ( n26851 ) ? ( VREG_3_6 ) : ( n26959 ) ;
assign n26961 =  ( n26850 ) ? ( VREG_3_7 ) : ( n26960 ) ;
assign n26962 =  ( n26849 ) ? ( VREG_3_8 ) : ( n26961 ) ;
assign n26963 =  ( n26848 ) ? ( VREG_3_9 ) : ( n26962 ) ;
assign n26964 =  ( n26847 ) ? ( VREG_3_10 ) : ( n26963 ) ;
assign n26965 =  ( n26846 ) ? ( VREG_3_11 ) : ( n26964 ) ;
assign n26966 =  ( n26845 ) ? ( VREG_3_12 ) : ( n26965 ) ;
assign n26967 =  ( n26844 ) ? ( VREG_3_13 ) : ( n26966 ) ;
assign n26968 =  ( n26843 ) ? ( VREG_3_14 ) : ( n26967 ) ;
assign n26969 =  ( n26842 ) ? ( VREG_3_15 ) : ( n26968 ) ;
assign n26970 =  ( n26841 ) ? ( VREG_4_0 ) : ( n26969 ) ;
assign n26971 =  ( n26840 ) ? ( VREG_4_1 ) : ( n26970 ) ;
assign n26972 =  ( n26839 ) ? ( VREG_4_2 ) : ( n26971 ) ;
assign n26973 =  ( n26838 ) ? ( VREG_4_3 ) : ( n26972 ) ;
assign n26974 =  ( n26837 ) ? ( VREG_4_4 ) : ( n26973 ) ;
assign n26975 =  ( n26836 ) ? ( VREG_4_5 ) : ( n26974 ) ;
assign n26976 =  ( n26835 ) ? ( VREG_4_6 ) : ( n26975 ) ;
assign n26977 =  ( n26834 ) ? ( VREG_4_7 ) : ( n26976 ) ;
assign n26978 =  ( n26833 ) ? ( VREG_4_8 ) : ( n26977 ) ;
assign n26979 =  ( n26832 ) ? ( VREG_4_9 ) : ( n26978 ) ;
assign n26980 =  ( n26831 ) ? ( VREG_4_10 ) : ( n26979 ) ;
assign n26981 =  ( n26830 ) ? ( VREG_4_11 ) : ( n26980 ) ;
assign n26982 =  ( n26829 ) ? ( VREG_4_12 ) : ( n26981 ) ;
assign n26983 =  ( n26828 ) ? ( VREG_4_13 ) : ( n26982 ) ;
assign n26984 =  ( n26827 ) ? ( VREG_4_14 ) : ( n26983 ) ;
assign n26985 =  ( n26826 ) ? ( VREG_4_15 ) : ( n26984 ) ;
assign n26986 =  ( n26825 ) ? ( VREG_5_0 ) : ( n26985 ) ;
assign n26987 =  ( n26824 ) ? ( VREG_5_1 ) : ( n26986 ) ;
assign n26988 =  ( n26823 ) ? ( VREG_5_2 ) : ( n26987 ) ;
assign n26989 =  ( n26822 ) ? ( VREG_5_3 ) : ( n26988 ) ;
assign n26990 =  ( n26821 ) ? ( VREG_5_4 ) : ( n26989 ) ;
assign n26991 =  ( n26820 ) ? ( VREG_5_5 ) : ( n26990 ) ;
assign n26992 =  ( n26819 ) ? ( VREG_5_6 ) : ( n26991 ) ;
assign n26993 =  ( n26818 ) ? ( VREG_5_7 ) : ( n26992 ) ;
assign n26994 =  ( n26817 ) ? ( VREG_5_8 ) : ( n26993 ) ;
assign n26995 =  ( n26816 ) ? ( VREG_5_9 ) : ( n26994 ) ;
assign n26996 =  ( n26815 ) ? ( VREG_5_10 ) : ( n26995 ) ;
assign n26997 =  ( n26814 ) ? ( VREG_5_11 ) : ( n26996 ) ;
assign n26998 =  ( n26813 ) ? ( VREG_5_12 ) : ( n26997 ) ;
assign n26999 =  ( n26812 ) ? ( VREG_5_13 ) : ( n26998 ) ;
assign n27000 =  ( n26811 ) ? ( VREG_5_14 ) : ( n26999 ) ;
assign n27001 =  ( n26810 ) ? ( VREG_5_15 ) : ( n27000 ) ;
assign n27002 =  ( n26809 ) ? ( VREG_6_0 ) : ( n27001 ) ;
assign n27003 =  ( n26808 ) ? ( VREG_6_1 ) : ( n27002 ) ;
assign n27004 =  ( n26807 ) ? ( VREG_6_2 ) : ( n27003 ) ;
assign n27005 =  ( n26806 ) ? ( VREG_6_3 ) : ( n27004 ) ;
assign n27006 =  ( n26805 ) ? ( VREG_6_4 ) : ( n27005 ) ;
assign n27007 =  ( n26804 ) ? ( VREG_6_5 ) : ( n27006 ) ;
assign n27008 =  ( n26803 ) ? ( VREG_6_6 ) : ( n27007 ) ;
assign n27009 =  ( n26802 ) ? ( VREG_6_7 ) : ( n27008 ) ;
assign n27010 =  ( n26801 ) ? ( VREG_6_8 ) : ( n27009 ) ;
assign n27011 =  ( n26800 ) ? ( VREG_6_9 ) : ( n27010 ) ;
assign n27012 =  ( n26799 ) ? ( VREG_6_10 ) : ( n27011 ) ;
assign n27013 =  ( n26798 ) ? ( VREG_6_11 ) : ( n27012 ) ;
assign n27014 =  ( n26797 ) ? ( VREG_6_12 ) : ( n27013 ) ;
assign n27015 =  ( n26796 ) ? ( VREG_6_13 ) : ( n27014 ) ;
assign n27016 =  ( n26795 ) ? ( VREG_6_14 ) : ( n27015 ) ;
assign n27017 =  ( n26794 ) ? ( VREG_6_15 ) : ( n27016 ) ;
assign n27018 =  ( n26793 ) ? ( VREG_7_0 ) : ( n27017 ) ;
assign n27019 =  ( n26792 ) ? ( VREG_7_1 ) : ( n27018 ) ;
assign n27020 =  ( n26791 ) ? ( VREG_7_2 ) : ( n27019 ) ;
assign n27021 =  ( n26790 ) ? ( VREG_7_3 ) : ( n27020 ) ;
assign n27022 =  ( n26789 ) ? ( VREG_7_4 ) : ( n27021 ) ;
assign n27023 =  ( n26788 ) ? ( VREG_7_5 ) : ( n27022 ) ;
assign n27024 =  ( n26787 ) ? ( VREG_7_6 ) : ( n27023 ) ;
assign n27025 =  ( n26786 ) ? ( VREG_7_7 ) : ( n27024 ) ;
assign n27026 =  ( n26785 ) ? ( VREG_7_8 ) : ( n27025 ) ;
assign n27027 =  ( n26784 ) ? ( VREG_7_9 ) : ( n27026 ) ;
assign n27028 =  ( n26783 ) ? ( VREG_7_10 ) : ( n27027 ) ;
assign n27029 =  ( n26782 ) ? ( VREG_7_11 ) : ( n27028 ) ;
assign n27030 =  ( n26781 ) ? ( VREG_7_12 ) : ( n27029 ) ;
assign n27031 =  ( n26780 ) ? ( VREG_7_13 ) : ( n27030 ) ;
assign n27032 =  ( n26779 ) ? ( VREG_7_14 ) : ( n27031 ) ;
assign n27033 =  ( n26778 ) ? ( VREG_7_15 ) : ( n27032 ) ;
assign n27034 =  ( n26777 ) ? ( VREG_8_0 ) : ( n27033 ) ;
assign n27035 =  ( n26776 ) ? ( VREG_8_1 ) : ( n27034 ) ;
assign n27036 =  ( n26775 ) ? ( VREG_8_2 ) : ( n27035 ) ;
assign n27037 =  ( n26774 ) ? ( VREG_8_3 ) : ( n27036 ) ;
assign n27038 =  ( n26773 ) ? ( VREG_8_4 ) : ( n27037 ) ;
assign n27039 =  ( n26772 ) ? ( VREG_8_5 ) : ( n27038 ) ;
assign n27040 =  ( n26771 ) ? ( VREG_8_6 ) : ( n27039 ) ;
assign n27041 =  ( n26770 ) ? ( VREG_8_7 ) : ( n27040 ) ;
assign n27042 =  ( n26769 ) ? ( VREG_8_8 ) : ( n27041 ) ;
assign n27043 =  ( n26768 ) ? ( VREG_8_9 ) : ( n27042 ) ;
assign n27044 =  ( n26767 ) ? ( VREG_8_10 ) : ( n27043 ) ;
assign n27045 =  ( n26766 ) ? ( VREG_8_11 ) : ( n27044 ) ;
assign n27046 =  ( n26765 ) ? ( VREG_8_12 ) : ( n27045 ) ;
assign n27047 =  ( n26764 ) ? ( VREG_8_13 ) : ( n27046 ) ;
assign n27048 =  ( n26763 ) ? ( VREG_8_14 ) : ( n27047 ) ;
assign n27049 =  ( n26762 ) ? ( VREG_8_15 ) : ( n27048 ) ;
assign n27050 =  ( n26761 ) ? ( VREG_9_0 ) : ( n27049 ) ;
assign n27051 =  ( n26760 ) ? ( VREG_9_1 ) : ( n27050 ) ;
assign n27052 =  ( n26759 ) ? ( VREG_9_2 ) : ( n27051 ) ;
assign n27053 =  ( n26758 ) ? ( VREG_9_3 ) : ( n27052 ) ;
assign n27054 =  ( n26757 ) ? ( VREG_9_4 ) : ( n27053 ) ;
assign n27055 =  ( n26756 ) ? ( VREG_9_5 ) : ( n27054 ) ;
assign n27056 =  ( n26755 ) ? ( VREG_9_6 ) : ( n27055 ) ;
assign n27057 =  ( n26754 ) ? ( VREG_9_7 ) : ( n27056 ) ;
assign n27058 =  ( n26753 ) ? ( VREG_9_8 ) : ( n27057 ) ;
assign n27059 =  ( n26752 ) ? ( VREG_9_9 ) : ( n27058 ) ;
assign n27060 =  ( n26751 ) ? ( VREG_9_10 ) : ( n27059 ) ;
assign n27061 =  ( n26750 ) ? ( VREG_9_11 ) : ( n27060 ) ;
assign n27062 =  ( n26749 ) ? ( VREG_9_12 ) : ( n27061 ) ;
assign n27063 =  ( n26748 ) ? ( VREG_9_13 ) : ( n27062 ) ;
assign n27064 =  ( n26747 ) ? ( VREG_9_14 ) : ( n27063 ) ;
assign n27065 =  ( n26746 ) ? ( VREG_9_15 ) : ( n27064 ) ;
assign n27066 =  ( n26745 ) ? ( VREG_10_0 ) : ( n27065 ) ;
assign n27067 =  ( n26744 ) ? ( VREG_10_1 ) : ( n27066 ) ;
assign n27068 =  ( n26743 ) ? ( VREG_10_2 ) : ( n27067 ) ;
assign n27069 =  ( n26742 ) ? ( VREG_10_3 ) : ( n27068 ) ;
assign n27070 =  ( n26741 ) ? ( VREG_10_4 ) : ( n27069 ) ;
assign n27071 =  ( n26740 ) ? ( VREG_10_5 ) : ( n27070 ) ;
assign n27072 =  ( n26739 ) ? ( VREG_10_6 ) : ( n27071 ) ;
assign n27073 =  ( n26738 ) ? ( VREG_10_7 ) : ( n27072 ) ;
assign n27074 =  ( n26737 ) ? ( VREG_10_8 ) : ( n27073 ) ;
assign n27075 =  ( n26736 ) ? ( VREG_10_9 ) : ( n27074 ) ;
assign n27076 =  ( n26735 ) ? ( VREG_10_10 ) : ( n27075 ) ;
assign n27077 =  ( n26734 ) ? ( VREG_10_11 ) : ( n27076 ) ;
assign n27078 =  ( n26733 ) ? ( VREG_10_12 ) : ( n27077 ) ;
assign n27079 =  ( n26732 ) ? ( VREG_10_13 ) : ( n27078 ) ;
assign n27080 =  ( n26731 ) ? ( VREG_10_14 ) : ( n27079 ) ;
assign n27081 =  ( n26730 ) ? ( VREG_10_15 ) : ( n27080 ) ;
assign n27082 =  ( n26729 ) ? ( VREG_11_0 ) : ( n27081 ) ;
assign n27083 =  ( n26728 ) ? ( VREG_11_1 ) : ( n27082 ) ;
assign n27084 =  ( n26727 ) ? ( VREG_11_2 ) : ( n27083 ) ;
assign n27085 =  ( n26726 ) ? ( VREG_11_3 ) : ( n27084 ) ;
assign n27086 =  ( n26725 ) ? ( VREG_11_4 ) : ( n27085 ) ;
assign n27087 =  ( n26724 ) ? ( VREG_11_5 ) : ( n27086 ) ;
assign n27088 =  ( n26723 ) ? ( VREG_11_6 ) : ( n27087 ) ;
assign n27089 =  ( n26722 ) ? ( VREG_11_7 ) : ( n27088 ) ;
assign n27090 =  ( n26721 ) ? ( VREG_11_8 ) : ( n27089 ) ;
assign n27091 =  ( n26720 ) ? ( VREG_11_9 ) : ( n27090 ) ;
assign n27092 =  ( n26719 ) ? ( VREG_11_10 ) : ( n27091 ) ;
assign n27093 =  ( n26718 ) ? ( VREG_11_11 ) : ( n27092 ) ;
assign n27094 =  ( n26717 ) ? ( VREG_11_12 ) : ( n27093 ) ;
assign n27095 =  ( n26716 ) ? ( VREG_11_13 ) : ( n27094 ) ;
assign n27096 =  ( n26715 ) ? ( VREG_11_14 ) : ( n27095 ) ;
assign n27097 =  ( n26714 ) ? ( VREG_11_15 ) : ( n27096 ) ;
assign n27098 =  ( n26713 ) ? ( VREG_12_0 ) : ( n27097 ) ;
assign n27099 =  ( n26712 ) ? ( VREG_12_1 ) : ( n27098 ) ;
assign n27100 =  ( n26711 ) ? ( VREG_12_2 ) : ( n27099 ) ;
assign n27101 =  ( n26710 ) ? ( VREG_12_3 ) : ( n27100 ) ;
assign n27102 =  ( n26709 ) ? ( VREG_12_4 ) : ( n27101 ) ;
assign n27103 =  ( n26708 ) ? ( VREG_12_5 ) : ( n27102 ) ;
assign n27104 =  ( n26707 ) ? ( VREG_12_6 ) : ( n27103 ) ;
assign n27105 =  ( n26706 ) ? ( VREG_12_7 ) : ( n27104 ) ;
assign n27106 =  ( n26705 ) ? ( VREG_12_8 ) : ( n27105 ) ;
assign n27107 =  ( n26704 ) ? ( VREG_12_9 ) : ( n27106 ) ;
assign n27108 =  ( n26703 ) ? ( VREG_12_10 ) : ( n27107 ) ;
assign n27109 =  ( n26702 ) ? ( VREG_12_11 ) : ( n27108 ) ;
assign n27110 =  ( n26701 ) ? ( VREG_12_12 ) : ( n27109 ) ;
assign n27111 =  ( n26700 ) ? ( VREG_12_13 ) : ( n27110 ) ;
assign n27112 =  ( n26699 ) ? ( VREG_12_14 ) : ( n27111 ) ;
assign n27113 =  ( n26698 ) ? ( VREG_12_15 ) : ( n27112 ) ;
assign n27114 =  ( n26697 ) ? ( VREG_13_0 ) : ( n27113 ) ;
assign n27115 =  ( n26696 ) ? ( VREG_13_1 ) : ( n27114 ) ;
assign n27116 =  ( n26695 ) ? ( VREG_13_2 ) : ( n27115 ) ;
assign n27117 =  ( n26694 ) ? ( VREG_13_3 ) : ( n27116 ) ;
assign n27118 =  ( n26693 ) ? ( VREG_13_4 ) : ( n27117 ) ;
assign n27119 =  ( n26692 ) ? ( VREG_13_5 ) : ( n27118 ) ;
assign n27120 =  ( n26691 ) ? ( VREG_13_6 ) : ( n27119 ) ;
assign n27121 =  ( n26690 ) ? ( VREG_13_7 ) : ( n27120 ) ;
assign n27122 =  ( n26689 ) ? ( VREG_13_8 ) : ( n27121 ) ;
assign n27123 =  ( n26688 ) ? ( VREG_13_9 ) : ( n27122 ) ;
assign n27124 =  ( n26687 ) ? ( VREG_13_10 ) : ( n27123 ) ;
assign n27125 =  ( n26686 ) ? ( VREG_13_11 ) : ( n27124 ) ;
assign n27126 =  ( n26685 ) ? ( VREG_13_12 ) : ( n27125 ) ;
assign n27127 =  ( n26684 ) ? ( VREG_13_13 ) : ( n27126 ) ;
assign n27128 =  ( n26683 ) ? ( VREG_13_14 ) : ( n27127 ) ;
assign n27129 =  ( n26682 ) ? ( VREG_13_15 ) : ( n27128 ) ;
assign n27130 =  ( n26681 ) ? ( VREG_14_0 ) : ( n27129 ) ;
assign n27131 =  ( n26680 ) ? ( VREG_14_1 ) : ( n27130 ) ;
assign n27132 =  ( n26679 ) ? ( VREG_14_2 ) : ( n27131 ) ;
assign n27133 =  ( n26678 ) ? ( VREG_14_3 ) : ( n27132 ) ;
assign n27134 =  ( n26677 ) ? ( VREG_14_4 ) : ( n27133 ) ;
assign n27135 =  ( n26676 ) ? ( VREG_14_5 ) : ( n27134 ) ;
assign n27136 =  ( n26675 ) ? ( VREG_14_6 ) : ( n27135 ) ;
assign n27137 =  ( n26674 ) ? ( VREG_14_7 ) : ( n27136 ) ;
assign n27138 =  ( n26673 ) ? ( VREG_14_8 ) : ( n27137 ) ;
assign n27139 =  ( n26672 ) ? ( VREG_14_9 ) : ( n27138 ) ;
assign n27140 =  ( n26671 ) ? ( VREG_14_10 ) : ( n27139 ) ;
assign n27141 =  ( n26670 ) ? ( VREG_14_11 ) : ( n27140 ) ;
assign n27142 =  ( n26669 ) ? ( VREG_14_12 ) : ( n27141 ) ;
assign n27143 =  ( n26668 ) ? ( VREG_14_13 ) : ( n27142 ) ;
assign n27144 =  ( n26667 ) ? ( VREG_14_14 ) : ( n27143 ) ;
assign n27145 =  ( n26666 ) ? ( VREG_14_15 ) : ( n27144 ) ;
assign n27146 =  ( n26665 ) ? ( VREG_15_0 ) : ( n27145 ) ;
assign n27147 =  ( n26664 ) ? ( VREG_15_1 ) : ( n27146 ) ;
assign n27148 =  ( n26663 ) ? ( VREG_15_2 ) : ( n27147 ) ;
assign n27149 =  ( n26662 ) ? ( VREG_15_3 ) : ( n27148 ) ;
assign n27150 =  ( n26661 ) ? ( VREG_15_4 ) : ( n27149 ) ;
assign n27151 =  ( n26660 ) ? ( VREG_15_5 ) : ( n27150 ) ;
assign n27152 =  ( n26659 ) ? ( VREG_15_6 ) : ( n27151 ) ;
assign n27153 =  ( n26658 ) ? ( VREG_15_7 ) : ( n27152 ) ;
assign n27154 =  ( n26657 ) ? ( VREG_15_8 ) : ( n27153 ) ;
assign n27155 =  ( n26656 ) ? ( VREG_15_9 ) : ( n27154 ) ;
assign n27156 =  ( n26655 ) ? ( VREG_15_10 ) : ( n27155 ) ;
assign n27157 =  ( n26654 ) ? ( VREG_15_11 ) : ( n27156 ) ;
assign n27158 =  ( n26653 ) ? ( VREG_15_12 ) : ( n27157 ) ;
assign n27159 =  ( n26652 ) ? ( VREG_15_13 ) : ( n27158 ) ;
assign n27160 =  ( n26651 ) ? ( VREG_15_14 ) : ( n27159 ) ;
assign n27161 =  ( n26650 ) ? ( VREG_15_15 ) : ( n27160 ) ;
assign n27162 =  ( n26649 ) ? ( VREG_16_0 ) : ( n27161 ) ;
assign n27163 =  ( n26648 ) ? ( VREG_16_1 ) : ( n27162 ) ;
assign n27164 =  ( n26647 ) ? ( VREG_16_2 ) : ( n27163 ) ;
assign n27165 =  ( n26646 ) ? ( VREG_16_3 ) : ( n27164 ) ;
assign n27166 =  ( n26645 ) ? ( VREG_16_4 ) : ( n27165 ) ;
assign n27167 =  ( n26644 ) ? ( VREG_16_5 ) : ( n27166 ) ;
assign n27168 =  ( n26643 ) ? ( VREG_16_6 ) : ( n27167 ) ;
assign n27169 =  ( n26642 ) ? ( VREG_16_7 ) : ( n27168 ) ;
assign n27170 =  ( n26641 ) ? ( VREG_16_8 ) : ( n27169 ) ;
assign n27171 =  ( n26640 ) ? ( VREG_16_9 ) : ( n27170 ) ;
assign n27172 =  ( n26639 ) ? ( VREG_16_10 ) : ( n27171 ) ;
assign n27173 =  ( n26638 ) ? ( VREG_16_11 ) : ( n27172 ) ;
assign n27174 =  ( n26637 ) ? ( VREG_16_12 ) : ( n27173 ) ;
assign n27175 =  ( n26636 ) ? ( VREG_16_13 ) : ( n27174 ) ;
assign n27176 =  ( n26635 ) ? ( VREG_16_14 ) : ( n27175 ) ;
assign n27177 =  ( n26634 ) ? ( VREG_16_15 ) : ( n27176 ) ;
assign n27178 =  ( n26633 ) ? ( VREG_17_0 ) : ( n27177 ) ;
assign n27179 =  ( n26632 ) ? ( VREG_17_1 ) : ( n27178 ) ;
assign n27180 =  ( n26631 ) ? ( VREG_17_2 ) : ( n27179 ) ;
assign n27181 =  ( n26630 ) ? ( VREG_17_3 ) : ( n27180 ) ;
assign n27182 =  ( n26629 ) ? ( VREG_17_4 ) : ( n27181 ) ;
assign n27183 =  ( n26628 ) ? ( VREG_17_5 ) : ( n27182 ) ;
assign n27184 =  ( n26627 ) ? ( VREG_17_6 ) : ( n27183 ) ;
assign n27185 =  ( n26626 ) ? ( VREG_17_7 ) : ( n27184 ) ;
assign n27186 =  ( n26625 ) ? ( VREG_17_8 ) : ( n27185 ) ;
assign n27187 =  ( n26624 ) ? ( VREG_17_9 ) : ( n27186 ) ;
assign n27188 =  ( n26623 ) ? ( VREG_17_10 ) : ( n27187 ) ;
assign n27189 =  ( n26622 ) ? ( VREG_17_11 ) : ( n27188 ) ;
assign n27190 =  ( n26621 ) ? ( VREG_17_12 ) : ( n27189 ) ;
assign n27191 =  ( n26620 ) ? ( VREG_17_13 ) : ( n27190 ) ;
assign n27192 =  ( n26619 ) ? ( VREG_17_14 ) : ( n27191 ) ;
assign n27193 =  ( n26618 ) ? ( VREG_17_15 ) : ( n27192 ) ;
assign n27194 =  ( n26617 ) ? ( VREG_18_0 ) : ( n27193 ) ;
assign n27195 =  ( n26616 ) ? ( VREG_18_1 ) : ( n27194 ) ;
assign n27196 =  ( n26615 ) ? ( VREG_18_2 ) : ( n27195 ) ;
assign n27197 =  ( n26614 ) ? ( VREG_18_3 ) : ( n27196 ) ;
assign n27198 =  ( n26613 ) ? ( VREG_18_4 ) : ( n27197 ) ;
assign n27199 =  ( n26612 ) ? ( VREG_18_5 ) : ( n27198 ) ;
assign n27200 =  ( n26611 ) ? ( VREG_18_6 ) : ( n27199 ) ;
assign n27201 =  ( n26610 ) ? ( VREG_18_7 ) : ( n27200 ) ;
assign n27202 =  ( n26609 ) ? ( VREG_18_8 ) : ( n27201 ) ;
assign n27203 =  ( n26608 ) ? ( VREG_18_9 ) : ( n27202 ) ;
assign n27204 =  ( n26607 ) ? ( VREG_18_10 ) : ( n27203 ) ;
assign n27205 =  ( n26606 ) ? ( VREG_18_11 ) : ( n27204 ) ;
assign n27206 =  ( n26605 ) ? ( VREG_18_12 ) : ( n27205 ) ;
assign n27207 =  ( n26604 ) ? ( VREG_18_13 ) : ( n27206 ) ;
assign n27208 =  ( n26603 ) ? ( VREG_18_14 ) : ( n27207 ) ;
assign n27209 =  ( n26602 ) ? ( VREG_18_15 ) : ( n27208 ) ;
assign n27210 =  ( n26601 ) ? ( VREG_19_0 ) : ( n27209 ) ;
assign n27211 =  ( n26600 ) ? ( VREG_19_1 ) : ( n27210 ) ;
assign n27212 =  ( n26599 ) ? ( VREG_19_2 ) : ( n27211 ) ;
assign n27213 =  ( n26598 ) ? ( VREG_19_3 ) : ( n27212 ) ;
assign n27214 =  ( n26597 ) ? ( VREG_19_4 ) : ( n27213 ) ;
assign n27215 =  ( n26596 ) ? ( VREG_19_5 ) : ( n27214 ) ;
assign n27216 =  ( n26595 ) ? ( VREG_19_6 ) : ( n27215 ) ;
assign n27217 =  ( n26594 ) ? ( VREG_19_7 ) : ( n27216 ) ;
assign n27218 =  ( n26593 ) ? ( VREG_19_8 ) : ( n27217 ) ;
assign n27219 =  ( n26592 ) ? ( VREG_19_9 ) : ( n27218 ) ;
assign n27220 =  ( n26591 ) ? ( VREG_19_10 ) : ( n27219 ) ;
assign n27221 =  ( n26590 ) ? ( VREG_19_11 ) : ( n27220 ) ;
assign n27222 =  ( n26589 ) ? ( VREG_19_12 ) : ( n27221 ) ;
assign n27223 =  ( n26588 ) ? ( VREG_19_13 ) : ( n27222 ) ;
assign n27224 =  ( n26587 ) ? ( VREG_19_14 ) : ( n27223 ) ;
assign n27225 =  ( n26586 ) ? ( VREG_19_15 ) : ( n27224 ) ;
assign n27226 =  ( n26585 ) ? ( VREG_20_0 ) : ( n27225 ) ;
assign n27227 =  ( n26584 ) ? ( VREG_20_1 ) : ( n27226 ) ;
assign n27228 =  ( n26583 ) ? ( VREG_20_2 ) : ( n27227 ) ;
assign n27229 =  ( n26582 ) ? ( VREG_20_3 ) : ( n27228 ) ;
assign n27230 =  ( n26581 ) ? ( VREG_20_4 ) : ( n27229 ) ;
assign n27231 =  ( n26580 ) ? ( VREG_20_5 ) : ( n27230 ) ;
assign n27232 =  ( n26579 ) ? ( VREG_20_6 ) : ( n27231 ) ;
assign n27233 =  ( n26578 ) ? ( VREG_20_7 ) : ( n27232 ) ;
assign n27234 =  ( n26577 ) ? ( VREG_20_8 ) : ( n27233 ) ;
assign n27235 =  ( n26576 ) ? ( VREG_20_9 ) : ( n27234 ) ;
assign n27236 =  ( n26575 ) ? ( VREG_20_10 ) : ( n27235 ) ;
assign n27237 =  ( n26574 ) ? ( VREG_20_11 ) : ( n27236 ) ;
assign n27238 =  ( n26573 ) ? ( VREG_20_12 ) : ( n27237 ) ;
assign n27239 =  ( n26572 ) ? ( VREG_20_13 ) : ( n27238 ) ;
assign n27240 =  ( n26571 ) ? ( VREG_20_14 ) : ( n27239 ) ;
assign n27241 =  ( n26570 ) ? ( VREG_20_15 ) : ( n27240 ) ;
assign n27242 =  ( n26569 ) ? ( VREG_21_0 ) : ( n27241 ) ;
assign n27243 =  ( n26568 ) ? ( VREG_21_1 ) : ( n27242 ) ;
assign n27244 =  ( n26567 ) ? ( VREG_21_2 ) : ( n27243 ) ;
assign n27245 =  ( n26566 ) ? ( VREG_21_3 ) : ( n27244 ) ;
assign n27246 =  ( n26565 ) ? ( VREG_21_4 ) : ( n27245 ) ;
assign n27247 =  ( n26564 ) ? ( VREG_21_5 ) : ( n27246 ) ;
assign n27248 =  ( n26563 ) ? ( VREG_21_6 ) : ( n27247 ) ;
assign n27249 =  ( n26562 ) ? ( VREG_21_7 ) : ( n27248 ) ;
assign n27250 =  ( n26561 ) ? ( VREG_21_8 ) : ( n27249 ) ;
assign n27251 =  ( n26560 ) ? ( VREG_21_9 ) : ( n27250 ) ;
assign n27252 =  ( n26559 ) ? ( VREG_21_10 ) : ( n27251 ) ;
assign n27253 =  ( n26558 ) ? ( VREG_21_11 ) : ( n27252 ) ;
assign n27254 =  ( n26557 ) ? ( VREG_21_12 ) : ( n27253 ) ;
assign n27255 =  ( n26556 ) ? ( VREG_21_13 ) : ( n27254 ) ;
assign n27256 =  ( n26555 ) ? ( VREG_21_14 ) : ( n27255 ) ;
assign n27257 =  ( n26554 ) ? ( VREG_21_15 ) : ( n27256 ) ;
assign n27258 =  ( n26553 ) ? ( VREG_22_0 ) : ( n27257 ) ;
assign n27259 =  ( n26552 ) ? ( VREG_22_1 ) : ( n27258 ) ;
assign n27260 =  ( n26551 ) ? ( VREG_22_2 ) : ( n27259 ) ;
assign n27261 =  ( n26550 ) ? ( VREG_22_3 ) : ( n27260 ) ;
assign n27262 =  ( n26549 ) ? ( VREG_22_4 ) : ( n27261 ) ;
assign n27263 =  ( n26548 ) ? ( VREG_22_5 ) : ( n27262 ) ;
assign n27264 =  ( n26547 ) ? ( VREG_22_6 ) : ( n27263 ) ;
assign n27265 =  ( n26546 ) ? ( VREG_22_7 ) : ( n27264 ) ;
assign n27266 =  ( n26545 ) ? ( VREG_22_8 ) : ( n27265 ) ;
assign n27267 =  ( n26544 ) ? ( VREG_22_9 ) : ( n27266 ) ;
assign n27268 =  ( n26543 ) ? ( VREG_22_10 ) : ( n27267 ) ;
assign n27269 =  ( n26542 ) ? ( VREG_22_11 ) : ( n27268 ) ;
assign n27270 =  ( n26541 ) ? ( VREG_22_12 ) : ( n27269 ) ;
assign n27271 =  ( n26540 ) ? ( VREG_22_13 ) : ( n27270 ) ;
assign n27272 =  ( n26539 ) ? ( VREG_22_14 ) : ( n27271 ) ;
assign n27273 =  ( n26538 ) ? ( VREG_22_15 ) : ( n27272 ) ;
assign n27274 =  ( n26537 ) ? ( VREG_23_0 ) : ( n27273 ) ;
assign n27275 =  ( n26536 ) ? ( VREG_23_1 ) : ( n27274 ) ;
assign n27276 =  ( n26535 ) ? ( VREG_23_2 ) : ( n27275 ) ;
assign n27277 =  ( n26534 ) ? ( VREG_23_3 ) : ( n27276 ) ;
assign n27278 =  ( n26533 ) ? ( VREG_23_4 ) : ( n27277 ) ;
assign n27279 =  ( n26532 ) ? ( VREG_23_5 ) : ( n27278 ) ;
assign n27280 =  ( n26531 ) ? ( VREG_23_6 ) : ( n27279 ) ;
assign n27281 =  ( n26530 ) ? ( VREG_23_7 ) : ( n27280 ) ;
assign n27282 =  ( n26529 ) ? ( VREG_23_8 ) : ( n27281 ) ;
assign n27283 =  ( n26528 ) ? ( VREG_23_9 ) : ( n27282 ) ;
assign n27284 =  ( n26527 ) ? ( VREG_23_10 ) : ( n27283 ) ;
assign n27285 =  ( n26526 ) ? ( VREG_23_11 ) : ( n27284 ) ;
assign n27286 =  ( n26525 ) ? ( VREG_23_12 ) : ( n27285 ) ;
assign n27287 =  ( n26524 ) ? ( VREG_23_13 ) : ( n27286 ) ;
assign n27288 =  ( n26523 ) ? ( VREG_23_14 ) : ( n27287 ) ;
assign n27289 =  ( n26522 ) ? ( VREG_23_15 ) : ( n27288 ) ;
assign n27290 =  ( n26521 ) ? ( VREG_24_0 ) : ( n27289 ) ;
assign n27291 =  ( n26520 ) ? ( VREG_24_1 ) : ( n27290 ) ;
assign n27292 =  ( n26519 ) ? ( VREG_24_2 ) : ( n27291 ) ;
assign n27293 =  ( n26518 ) ? ( VREG_24_3 ) : ( n27292 ) ;
assign n27294 =  ( n26517 ) ? ( VREG_24_4 ) : ( n27293 ) ;
assign n27295 =  ( n26516 ) ? ( VREG_24_5 ) : ( n27294 ) ;
assign n27296 =  ( n26515 ) ? ( VREG_24_6 ) : ( n27295 ) ;
assign n27297 =  ( n26514 ) ? ( VREG_24_7 ) : ( n27296 ) ;
assign n27298 =  ( n26513 ) ? ( VREG_24_8 ) : ( n27297 ) ;
assign n27299 =  ( n26512 ) ? ( VREG_24_9 ) : ( n27298 ) ;
assign n27300 =  ( n26511 ) ? ( VREG_24_10 ) : ( n27299 ) ;
assign n27301 =  ( n26510 ) ? ( VREG_24_11 ) : ( n27300 ) ;
assign n27302 =  ( n26509 ) ? ( VREG_24_12 ) : ( n27301 ) ;
assign n27303 =  ( n26508 ) ? ( VREG_24_13 ) : ( n27302 ) ;
assign n27304 =  ( n26507 ) ? ( VREG_24_14 ) : ( n27303 ) ;
assign n27305 =  ( n26506 ) ? ( VREG_24_15 ) : ( n27304 ) ;
assign n27306 =  ( n26505 ) ? ( VREG_25_0 ) : ( n27305 ) ;
assign n27307 =  ( n26504 ) ? ( VREG_25_1 ) : ( n27306 ) ;
assign n27308 =  ( n26503 ) ? ( VREG_25_2 ) : ( n27307 ) ;
assign n27309 =  ( n26502 ) ? ( VREG_25_3 ) : ( n27308 ) ;
assign n27310 =  ( n26501 ) ? ( VREG_25_4 ) : ( n27309 ) ;
assign n27311 =  ( n26500 ) ? ( VREG_25_5 ) : ( n27310 ) ;
assign n27312 =  ( n26499 ) ? ( VREG_25_6 ) : ( n27311 ) ;
assign n27313 =  ( n26498 ) ? ( VREG_25_7 ) : ( n27312 ) ;
assign n27314 =  ( n26497 ) ? ( VREG_25_8 ) : ( n27313 ) ;
assign n27315 =  ( n26496 ) ? ( VREG_25_9 ) : ( n27314 ) ;
assign n27316 =  ( n26495 ) ? ( VREG_25_10 ) : ( n27315 ) ;
assign n27317 =  ( n26494 ) ? ( VREG_25_11 ) : ( n27316 ) ;
assign n27318 =  ( n26493 ) ? ( VREG_25_12 ) : ( n27317 ) ;
assign n27319 =  ( n26492 ) ? ( VREG_25_13 ) : ( n27318 ) ;
assign n27320 =  ( n26491 ) ? ( VREG_25_14 ) : ( n27319 ) ;
assign n27321 =  ( n26490 ) ? ( VREG_25_15 ) : ( n27320 ) ;
assign n27322 =  ( n26489 ) ? ( VREG_26_0 ) : ( n27321 ) ;
assign n27323 =  ( n26488 ) ? ( VREG_26_1 ) : ( n27322 ) ;
assign n27324 =  ( n26487 ) ? ( VREG_26_2 ) : ( n27323 ) ;
assign n27325 =  ( n26486 ) ? ( VREG_26_3 ) : ( n27324 ) ;
assign n27326 =  ( n26485 ) ? ( VREG_26_4 ) : ( n27325 ) ;
assign n27327 =  ( n26484 ) ? ( VREG_26_5 ) : ( n27326 ) ;
assign n27328 =  ( n26483 ) ? ( VREG_26_6 ) : ( n27327 ) ;
assign n27329 =  ( n26482 ) ? ( VREG_26_7 ) : ( n27328 ) ;
assign n27330 =  ( n26481 ) ? ( VREG_26_8 ) : ( n27329 ) ;
assign n27331 =  ( n26480 ) ? ( VREG_26_9 ) : ( n27330 ) ;
assign n27332 =  ( n26479 ) ? ( VREG_26_10 ) : ( n27331 ) ;
assign n27333 =  ( n26478 ) ? ( VREG_26_11 ) : ( n27332 ) ;
assign n27334 =  ( n26477 ) ? ( VREG_26_12 ) : ( n27333 ) ;
assign n27335 =  ( n26476 ) ? ( VREG_26_13 ) : ( n27334 ) ;
assign n27336 =  ( n26475 ) ? ( VREG_26_14 ) : ( n27335 ) ;
assign n27337 =  ( n26474 ) ? ( VREG_26_15 ) : ( n27336 ) ;
assign n27338 =  ( n26473 ) ? ( VREG_27_0 ) : ( n27337 ) ;
assign n27339 =  ( n26472 ) ? ( VREG_27_1 ) : ( n27338 ) ;
assign n27340 =  ( n26471 ) ? ( VREG_27_2 ) : ( n27339 ) ;
assign n27341 =  ( n26470 ) ? ( VREG_27_3 ) : ( n27340 ) ;
assign n27342 =  ( n26469 ) ? ( VREG_27_4 ) : ( n27341 ) ;
assign n27343 =  ( n26468 ) ? ( VREG_27_5 ) : ( n27342 ) ;
assign n27344 =  ( n26467 ) ? ( VREG_27_6 ) : ( n27343 ) ;
assign n27345 =  ( n26466 ) ? ( VREG_27_7 ) : ( n27344 ) ;
assign n27346 =  ( n26465 ) ? ( VREG_27_8 ) : ( n27345 ) ;
assign n27347 =  ( n26464 ) ? ( VREG_27_9 ) : ( n27346 ) ;
assign n27348 =  ( n26463 ) ? ( VREG_27_10 ) : ( n27347 ) ;
assign n27349 =  ( n26462 ) ? ( VREG_27_11 ) : ( n27348 ) ;
assign n27350 =  ( n26461 ) ? ( VREG_27_12 ) : ( n27349 ) ;
assign n27351 =  ( n26460 ) ? ( VREG_27_13 ) : ( n27350 ) ;
assign n27352 =  ( n26459 ) ? ( VREG_27_14 ) : ( n27351 ) ;
assign n27353 =  ( n26458 ) ? ( VREG_27_15 ) : ( n27352 ) ;
assign n27354 =  ( n26457 ) ? ( VREG_28_0 ) : ( n27353 ) ;
assign n27355 =  ( n26456 ) ? ( VREG_28_1 ) : ( n27354 ) ;
assign n27356 =  ( n26455 ) ? ( VREG_28_2 ) : ( n27355 ) ;
assign n27357 =  ( n26454 ) ? ( VREG_28_3 ) : ( n27356 ) ;
assign n27358 =  ( n26453 ) ? ( VREG_28_4 ) : ( n27357 ) ;
assign n27359 =  ( n26452 ) ? ( VREG_28_5 ) : ( n27358 ) ;
assign n27360 =  ( n26451 ) ? ( VREG_28_6 ) : ( n27359 ) ;
assign n27361 =  ( n26450 ) ? ( VREG_28_7 ) : ( n27360 ) ;
assign n27362 =  ( n26449 ) ? ( VREG_28_8 ) : ( n27361 ) ;
assign n27363 =  ( n26448 ) ? ( VREG_28_9 ) : ( n27362 ) ;
assign n27364 =  ( n26447 ) ? ( VREG_28_10 ) : ( n27363 ) ;
assign n27365 =  ( n26446 ) ? ( VREG_28_11 ) : ( n27364 ) ;
assign n27366 =  ( n26445 ) ? ( VREG_28_12 ) : ( n27365 ) ;
assign n27367 =  ( n26444 ) ? ( VREG_28_13 ) : ( n27366 ) ;
assign n27368 =  ( n26443 ) ? ( VREG_28_14 ) : ( n27367 ) ;
assign n27369 =  ( n26442 ) ? ( VREG_28_15 ) : ( n27368 ) ;
assign n27370 =  ( n26441 ) ? ( VREG_29_0 ) : ( n27369 ) ;
assign n27371 =  ( n26440 ) ? ( VREG_29_1 ) : ( n27370 ) ;
assign n27372 =  ( n26439 ) ? ( VREG_29_2 ) : ( n27371 ) ;
assign n27373 =  ( n26438 ) ? ( VREG_29_3 ) : ( n27372 ) ;
assign n27374 =  ( n26437 ) ? ( VREG_29_4 ) : ( n27373 ) ;
assign n27375 =  ( n26436 ) ? ( VREG_29_5 ) : ( n27374 ) ;
assign n27376 =  ( n26435 ) ? ( VREG_29_6 ) : ( n27375 ) ;
assign n27377 =  ( n26434 ) ? ( VREG_29_7 ) : ( n27376 ) ;
assign n27378 =  ( n26433 ) ? ( VREG_29_8 ) : ( n27377 ) ;
assign n27379 =  ( n26432 ) ? ( VREG_29_9 ) : ( n27378 ) ;
assign n27380 =  ( n26431 ) ? ( VREG_29_10 ) : ( n27379 ) ;
assign n27381 =  ( n26430 ) ? ( VREG_29_11 ) : ( n27380 ) ;
assign n27382 =  ( n26429 ) ? ( VREG_29_12 ) : ( n27381 ) ;
assign n27383 =  ( n26428 ) ? ( VREG_29_13 ) : ( n27382 ) ;
assign n27384 =  ( n26427 ) ? ( VREG_29_14 ) : ( n27383 ) ;
assign n27385 =  ( n26426 ) ? ( VREG_29_15 ) : ( n27384 ) ;
assign n27386 =  ( n26425 ) ? ( VREG_30_0 ) : ( n27385 ) ;
assign n27387 =  ( n26424 ) ? ( VREG_30_1 ) : ( n27386 ) ;
assign n27388 =  ( n26423 ) ? ( VREG_30_2 ) : ( n27387 ) ;
assign n27389 =  ( n26422 ) ? ( VREG_30_3 ) : ( n27388 ) ;
assign n27390 =  ( n26421 ) ? ( VREG_30_4 ) : ( n27389 ) ;
assign n27391 =  ( n26420 ) ? ( VREG_30_5 ) : ( n27390 ) ;
assign n27392 =  ( n26419 ) ? ( VREG_30_6 ) : ( n27391 ) ;
assign n27393 =  ( n26418 ) ? ( VREG_30_7 ) : ( n27392 ) ;
assign n27394 =  ( n26417 ) ? ( VREG_30_8 ) : ( n27393 ) ;
assign n27395 =  ( n26416 ) ? ( VREG_30_9 ) : ( n27394 ) ;
assign n27396 =  ( n26415 ) ? ( VREG_30_10 ) : ( n27395 ) ;
assign n27397 =  ( n26414 ) ? ( VREG_30_11 ) : ( n27396 ) ;
assign n27398 =  ( n26413 ) ? ( VREG_30_12 ) : ( n27397 ) ;
assign n27399 =  ( n26412 ) ? ( VREG_30_13 ) : ( n27398 ) ;
assign n27400 =  ( n26411 ) ? ( VREG_30_14 ) : ( n27399 ) ;
assign n27401 =  ( n26410 ) ? ( VREG_30_15 ) : ( n27400 ) ;
assign n27402 =  ( n26409 ) ? ( VREG_31_0 ) : ( n27401 ) ;
assign n27403 =  ( n26407 ) ? ( VREG_31_1 ) : ( n27402 ) ;
assign n27404 =  ( n26405 ) ? ( VREG_31_2 ) : ( n27403 ) ;
assign n27405 =  ( n26403 ) ? ( VREG_31_3 ) : ( n27404 ) ;
assign n27406 =  ( n26401 ) ? ( VREG_31_4 ) : ( n27405 ) ;
assign n27407 =  ( n26399 ) ? ( VREG_31_5 ) : ( n27406 ) ;
assign n27408 =  ( n26397 ) ? ( VREG_31_6 ) : ( n27407 ) ;
assign n27409 =  ( n26395 ) ? ( VREG_31_7 ) : ( n27408 ) ;
assign n27410 =  ( n26393 ) ? ( VREG_31_8 ) : ( n27409 ) ;
assign n27411 =  ( n26391 ) ? ( VREG_31_9 ) : ( n27410 ) ;
assign n27412 =  ( n26389 ) ? ( VREG_31_10 ) : ( n27411 ) ;
assign n27413 =  ( n26387 ) ? ( VREG_31_11 ) : ( n27412 ) ;
assign n27414 =  ( n26385 ) ? ( VREG_31_12 ) : ( n27413 ) ;
assign n27415 =  ( n26383 ) ? ( VREG_31_13 ) : ( n27414 ) ;
assign n27416 =  ( n26381 ) ? ( VREG_31_14 ) : ( n27415 ) ;
assign n27417 =  ( n26379 ) ? ( VREG_31_15 ) : ( n27416 ) ;
assign n27418 =  ( n27417 ) + ( n140 )  ;
assign n27419 =  ( n27417 ) - ( n140 )  ;
assign n27420 =  ( n27417 ) & ( n140 )  ;
assign n27421 =  ( n27417 ) | ( n140 )  ;
assign n27422 =  ( ( n27417 ) * ( n140 ))  ;
assign n27423 =  ( n148 ) ? ( n27422 ) : ( VREG_0_6 ) ;
assign n27424 =  ( n146 ) ? ( n27421 ) : ( n27423 ) ;
assign n27425 =  ( n144 ) ? ( n27420 ) : ( n27424 ) ;
assign n27426 =  ( n142 ) ? ( n27419 ) : ( n27425 ) ;
assign n27427 =  ( n10 ) ? ( n27418 ) : ( n27426 ) ;
assign n27428 =  ( n77 ) & ( n26378 )  ;
assign n27429 =  ( n77 ) & ( n26380 )  ;
assign n27430 =  ( n77 ) & ( n26382 )  ;
assign n27431 =  ( n77 ) & ( n26384 )  ;
assign n27432 =  ( n77 ) & ( n26386 )  ;
assign n27433 =  ( n77 ) & ( n26388 )  ;
assign n27434 =  ( n77 ) & ( n26390 )  ;
assign n27435 =  ( n77 ) & ( n26392 )  ;
assign n27436 =  ( n77 ) & ( n26394 )  ;
assign n27437 =  ( n77 ) & ( n26396 )  ;
assign n27438 =  ( n77 ) & ( n26398 )  ;
assign n27439 =  ( n77 ) & ( n26400 )  ;
assign n27440 =  ( n77 ) & ( n26402 )  ;
assign n27441 =  ( n77 ) & ( n26404 )  ;
assign n27442 =  ( n77 ) & ( n26406 )  ;
assign n27443 =  ( n77 ) & ( n26408 )  ;
assign n27444 =  ( n78 ) & ( n26378 )  ;
assign n27445 =  ( n78 ) & ( n26380 )  ;
assign n27446 =  ( n78 ) & ( n26382 )  ;
assign n27447 =  ( n78 ) & ( n26384 )  ;
assign n27448 =  ( n78 ) & ( n26386 )  ;
assign n27449 =  ( n78 ) & ( n26388 )  ;
assign n27450 =  ( n78 ) & ( n26390 )  ;
assign n27451 =  ( n78 ) & ( n26392 )  ;
assign n27452 =  ( n78 ) & ( n26394 )  ;
assign n27453 =  ( n78 ) & ( n26396 )  ;
assign n27454 =  ( n78 ) & ( n26398 )  ;
assign n27455 =  ( n78 ) & ( n26400 )  ;
assign n27456 =  ( n78 ) & ( n26402 )  ;
assign n27457 =  ( n78 ) & ( n26404 )  ;
assign n27458 =  ( n78 ) & ( n26406 )  ;
assign n27459 =  ( n78 ) & ( n26408 )  ;
assign n27460 =  ( n79 ) & ( n26378 )  ;
assign n27461 =  ( n79 ) & ( n26380 )  ;
assign n27462 =  ( n79 ) & ( n26382 )  ;
assign n27463 =  ( n79 ) & ( n26384 )  ;
assign n27464 =  ( n79 ) & ( n26386 )  ;
assign n27465 =  ( n79 ) & ( n26388 )  ;
assign n27466 =  ( n79 ) & ( n26390 )  ;
assign n27467 =  ( n79 ) & ( n26392 )  ;
assign n27468 =  ( n79 ) & ( n26394 )  ;
assign n27469 =  ( n79 ) & ( n26396 )  ;
assign n27470 =  ( n79 ) & ( n26398 )  ;
assign n27471 =  ( n79 ) & ( n26400 )  ;
assign n27472 =  ( n79 ) & ( n26402 )  ;
assign n27473 =  ( n79 ) & ( n26404 )  ;
assign n27474 =  ( n79 ) & ( n26406 )  ;
assign n27475 =  ( n79 ) & ( n26408 )  ;
assign n27476 =  ( n80 ) & ( n26378 )  ;
assign n27477 =  ( n80 ) & ( n26380 )  ;
assign n27478 =  ( n80 ) & ( n26382 )  ;
assign n27479 =  ( n80 ) & ( n26384 )  ;
assign n27480 =  ( n80 ) & ( n26386 )  ;
assign n27481 =  ( n80 ) & ( n26388 )  ;
assign n27482 =  ( n80 ) & ( n26390 )  ;
assign n27483 =  ( n80 ) & ( n26392 )  ;
assign n27484 =  ( n80 ) & ( n26394 )  ;
assign n27485 =  ( n80 ) & ( n26396 )  ;
assign n27486 =  ( n80 ) & ( n26398 )  ;
assign n27487 =  ( n80 ) & ( n26400 )  ;
assign n27488 =  ( n80 ) & ( n26402 )  ;
assign n27489 =  ( n80 ) & ( n26404 )  ;
assign n27490 =  ( n80 ) & ( n26406 )  ;
assign n27491 =  ( n80 ) & ( n26408 )  ;
assign n27492 =  ( n81 ) & ( n26378 )  ;
assign n27493 =  ( n81 ) & ( n26380 )  ;
assign n27494 =  ( n81 ) & ( n26382 )  ;
assign n27495 =  ( n81 ) & ( n26384 )  ;
assign n27496 =  ( n81 ) & ( n26386 )  ;
assign n27497 =  ( n81 ) & ( n26388 )  ;
assign n27498 =  ( n81 ) & ( n26390 )  ;
assign n27499 =  ( n81 ) & ( n26392 )  ;
assign n27500 =  ( n81 ) & ( n26394 )  ;
assign n27501 =  ( n81 ) & ( n26396 )  ;
assign n27502 =  ( n81 ) & ( n26398 )  ;
assign n27503 =  ( n81 ) & ( n26400 )  ;
assign n27504 =  ( n81 ) & ( n26402 )  ;
assign n27505 =  ( n81 ) & ( n26404 )  ;
assign n27506 =  ( n81 ) & ( n26406 )  ;
assign n27507 =  ( n81 ) & ( n26408 )  ;
assign n27508 =  ( n82 ) & ( n26378 )  ;
assign n27509 =  ( n82 ) & ( n26380 )  ;
assign n27510 =  ( n82 ) & ( n26382 )  ;
assign n27511 =  ( n82 ) & ( n26384 )  ;
assign n27512 =  ( n82 ) & ( n26386 )  ;
assign n27513 =  ( n82 ) & ( n26388 )  ;
assign n27514 =  ( n82 ) & ( n26390 )  ;
assign n27515 =  ( n82 ) & ( n26392 )  ;
assign n27516 =  ( n82 ) & ( n26394 )  ;
assign n27517 =  ( n82 ) & ( n26396 )  ;
assign n27518 =  ( n82 ) & ( n26398 )  ;
assign n27519 =  ( n82 ) & ( n26400 )  ;
assign n27520 =  ( n82 ) & ( n26402 )  ;
assign n27521 =  ( n82 ) & ( n26404 )  ;
assign n27522 =  ( n82 ) & ( n26406 )  ;
assign n27523 =  ( n82 ) & ( n26408 )  ;
assign n27524 =  ( n83 ) & ( n26378 )  ;
assign n27525 =  ( n83 ) & ( n26380 )  ;
assign n27526 =  ( n83 ) & ( n26382 )  ;
assign n27527 =  ( n83 ) & ( n26384 )  ;
assign n27528 =  ( n83 ) & ( n26386 )  ;
assign n27529 =  ( n83 ) & ( n26388 )  ;
assign n27530 =  ( n83 ) & ( n26390 )  ;
assign n27531 =  ( n83 ) & ( n26392 )  ;
assign n27532 =  ( n83 ) & ( n26394 )  ;
assign n27533 =  ( n83 ) & ( n26396 )  ;
assign n27534 =  ( n83 ) & ( n26398 )  ;
assign n27535 =  ( n83 ) & ( n26400 )  ;
assign n27536 =  ( n83 ) & ( n26402 )  ;
assign n27537 =  ( n83 ) & ( n26404 )  ;
assign n27538 =  ( n83 ) & ( n26406 )  ;
assign n27539 =  ( n83 ) & ( n26408 )  ;
assign n27540 =  ( n84 ) & ( n26378 )  ;
assign n27541 =  ( n84 ) & ( n26380 )  ;
assign n27542 =  ( n84 ) & ( n26382 )  ;
assign n27543 =  ( n84 ) & ( n26384 )  ;
assign n27544 =  ( n84 ) & ( n26386 )  ;
assign n27545 =  ( n84 ) & ( n26388 )  ;
assign n27546 =  ( n84 ) & ( n26390 )  ;
assign n27547 =  ( n84 ) & ( n26392 )  ;
assign n27548 =  ( n84 ) & ( n26394 )  ;
assign n27549 =  ( n84 ) & ( n26396 )  ;
assign n27550 =  ( n84 ) & ( n26398 )  ;
assign n27551 =  ( n84 ) & ( n26400 )  ;
assign n27552 =  ( n84 ) & ( n26402 )  ;
assign n27553 =  ( n84 ) & ( n26404 )  ;
assign n27554 =  ( n84 ) & ( n26406 )  ;
assign n27555 =  ( n84 ) & ( n26408 )  ;
assign n27556 =  ( n85 ) & ( n26378 )  ;
assign n27557 =  ( n85 ) & ( n26380 )  ;
assign n27558 =  ( n85 ) & ( n26382 )  ;
assign n27559 =  ( n85 ) & ( n26384 )  ;
assign n27560 =  ( n85 ) & ( n26386 )  ;
assign n27561 =  ( n85 ) & ( n26388 )  ;
assign n27562 =  ( n85 ) & ( n26390 )  ;
assign n27563 =  ( n85 ) & ( n26392 )  ;
assign n27564 =  ( n85 ) & ( n26394 )  ;
assign n27565 =  ( n85 ) & ( n26396 )  ;
assign n27566 =  ( n85 ) & ( n26398 )  ;
assign n27567 =  ( n85 ) & ( n26400 )  ;
assign n27568 =  ( n85 ) & ( n26402 )  ;
assign n27569 =  ( n85 ) & ( n26404 )  ;
assign n27570 =  ( n85 ) & ( n26406 )  ;
assign n27571 =  ( n85 ) & ( n26408 )  ;
assign n27572 =  ( n86 ) & ( n26378 )  ;
assign n27573 =  ( n86 ) & ( n26380 )  ;
assign n27574 =  ( n86 ) & ( n26382 )  ;
assign n27575 =  ( n86 ) & ( n26384 )  ;
assign n27576 =  ( n86 ) & ( n26386 )  ;
assign n27577 =  ( n86 ) & ( n26388 )  ;
assign n27578 =  ( n86 ) & ( n26390 )  ;
assign n27579 =  ( n86 ) & ( n26392 )  ;
assign n27580 =  ( n86 ) & ( n26394 )  ;
assign n27581 =  ( n86 ) & ( n26396 )  ;
assign n27582 =  ( n86 ) & ( n26398 )  ;
assign n27583 =  ( n86 ) & ( n26400 )  ;
assign n27584 =  ( n86 ) & ( n26402 )  ;
assign n27585 =  ( n86 ) & ( n26404 )  ;
assign n27586 =  ( n86 ) & ( n26406 )  ;
assign n27587 =  ( n86 ) & ( n26408 )  ;
assign n27588 =  ( n87 ) & ( n26378 )  ;
assign n27589 =  ( n87 ) & ( n26380 )  ;
assign n27590 =  ( n87 ) & ( n26382 )  ;
assign n27591 =  ( n87 ) & ( n26384 )  ;
assign n27592 =  ( n87 ) & ( n26386 )  ;
assign n27593 =  ( n87 ) & ( n26388 )  ;
assign n27594 =  ( n87 ) & ( n26390 )  ;
assign n27595 =  ( n87 ) & ( n26392 )  ;
assign n27596 =  ( n87 ) & ( n26394 )  ;
assign n27597 =  ( n87 ) & ( n26396 )  ;
assign n27598 =  ( n87 ) & ( n26398 )  ;
assign n27599 =  ( n87 ) & ( n26400 )  ;
assign n27600 =  ( n87 ) & ( n26402 )  ;
assign n27601 =  ( n87 ) & ( n26404 )  ;
assign n27602 =  ( n87 ) & ( n26406 )  ;
assign n27603 =  ( n87 ) & ( n26408 )  ;
assign n27604 =  ( n88 ) & ( n26378 )  ;
assign n27605 =  ( n88 ) & ( n26380 )  ;
assign n27606 =  ( n88 ) & ( n26382 )  ;
assign n27607 =  ( n88 ) & ( n26384 )  ;
assign n27608 =  ( n88 ) & ( n26386 )  ;
assign n27609 =  ( n88 ) & ( n26388 )  ;
assign n27610 =  ( n88 ) & ( n26390 )  ;
assign n27611 =  ( n88 ) & ( n26392 )  ;
assign n27612 =  ( n88 ) & ( n26394 )  ;
assign n27613 =  ( n88 ) & ( n26396 )  ;
assign n27614 =  ( n88 ) & ( n26398 )  ;
assign n27615 =  ( n88 ) & ( n26400 )  ;
assign n27616 =  ( n88 ) & ( n26402 )  ;
assign n27617 =  ( n88 ) & ( n26404 )  ;
assign n27618 =  ( n88 ) & ( n26406 )  ;
assign n27619 =  ( n88 ) & ( n26408 )  ;
assign n27620 =  ( n89 ) & ( n26378 )  ;
assign n27621 =  ( n89 ) & ( n26380 )  ;
assign n27622 =  ( n89 ) & ( n26382 )  ;
assign n27623 =  ( n89 ) & ( n26384 )  ;
assign n27624 =  ( n89 ) & ( n26386 )  ;
assign n27625 =  ( n89 ) & ( n26388 )  ;
assign n27626 =  ( n89 ) & ( n26390 )  ;
assign n27627 =  ( n89 ) & ( n26392 )  ;
assign n27628 =  ( n89 ) & ( n26394 )  ;
assign n27629 =  ( n89 ) & ( n26396 )  ;
assign n27630 =  ( n89 ) & ( n26398 )  ;
assign n27631 =  ( n89 ) & ( n26400 )  ;
assign n27632 =  ( n89 ) & ( n26402 )  ;
assign n27633 =  ( n89 ) & ( n26404 )  ;
assign n27634 =  ( n89 ) & ( n26406 )  ;
assign n27635 =  ( n89 ) & ( n26408 )  ;
assign n27636 =  ( n90 ) & ( n26378 )  ;
assign n27637 =  ( n90 ) & ( n26380 )  ;
assign n27638 =  ( n90 ) & ( n26382 )  ;
assign n27639 =  ( n90 ) & ( n26384 )  ;
assign n27640 =  ( n90 ) & ( n26386 )  ;
assign n27641 =  ( n90 ) & ( n26388 )  ;
assign n27642 =  ( n90 ) & ( n26390 )  ;
assign n27643 =  ( n90 ) & ( n26392 )  ;
assign n27644 =  ( n90 ) & ( n26394 )  ;
assign n27645 =  ( n90 ) & ( n26396 )  ;
assign n27646 =  ( n90 ) & ( n26398 )  ;
assign n27647 =  ( n90 ) & ( n26400 )  ;
assign n27648 =  ( n90 ) & ( n26402 )  ;
assign n27649 =  ( n90 ) & ( n26404 )  ;
assign n27650 =  ( n90 ) & ( n26406 )  ;
assign n27651 =  ( n90 ) & ( n26408 )  ;
assign n27652 =  ( n91 ) & ( n26378 )  ;
assign n27653 =  ( n91 ) & ( n26380 )  ;
assign n27654 =  ( n91 ) & ( n26382 )  ;
assign n27655 =  ( n91 ) & ( n26384 )  ;
assign n27656 =  ( n91 ) & ( n26386 )  ;
assign n27657 =  ( n91 ) & ( n26388 )  ;
assign n27658 =  ( n91 ) & ( n26390 )  ;
assign n27659 =  ( n91 ) & ( n26392 )  ;
assign n27660 =  ( n91 ) & ( n26394 )  ;
assign n27661 =  ( n91 ) & ( n26396 )  ;
assign n27662 =  ( n91 ) & ( n26398 )  ;
assign n27663 =  ( n91 ) & ( n26400 )  ;
assign n27664 =  ( n91 ) & ( n26402 )  ;
assign n27665 =  ( n91 ) & ( n26404 )  ;
assign n27666 =  ( n91 ) & ( n26406 )  ;
assign n27667 =  ( n91 ) & ( n26408 )  ;
assign n27668 =  ( n92 ) & ( n26378 )  ;
assign n27669 =  ( n92 ) & ( n26380 )  ;
assign n27670 =  ( n92 ) & ( n26382 )  ;
assign n27671 =  ( n92 ) & ( n26384 )  ;
assign n27672 =  ( n92 ) & ( n26386 )  ;
assign n27673 =  ( n92 ) & ( n26388 )  ;
assign n27674 =  ( n92 ) & ( n26390 )  ;
assign n27675 =  ( n92 ) & ( n26392 )  ;
assign n27676 =  ( n92 ) & ( n26394 )  ;
assign n27677 =  ( n92 ) & ( n26396 )  ;
assign n27678 =  ( n92 ) & ( n26398 )  ;
assign n27679 =  ( n92 ) & ( n26400 )  ;
assign n27680 =  ( n92 ) & ( n26402 )  ;
assign n27681 =  ( n92 ) & ( n26404 )  ;
assign n27682 =  ( n92 ) & ( n26406 )  ;
assign n27683 =  ( n92 ) & ( n26408 )  ;
assign n27684 =  ( n93 ) & ( n26378 )  ;
assign n27685 =  ( n93 ) & ( n26380 )  ;
assign n27686 =  ( n93 ) & ( n26382 )  ;
assign n27687 =  ( n93 ) & ( n26384 )  ;
assign n27688 =  ( n93 ) & ( n26386 )  ;
assign n27689 =  ( n93 ) & ( n26388 )  ;
assign n27690 =  ( n93 ) & ( n26390 )  ;
assign n27691 =  ( n93 ) & ( n26392 )  ;
assign n27692 =  ( n93 ) & ( n26394 )  ;
assign n27693 =  ( n93 ) & ( n26396 )  ;
assign n27694 =  ( n93 ) & ( n26398 )  ;
assign n27695 =  ( n93 ) & ( n26400 )  ;
assign n27696 =  ( n93 ) & ( n26402 )  ;
assign n27697 =  ( n93 ) & ( n26404 )  ;
assign n27698 =  ( n93 ) & ( n26406 )  ;
assign n27699 =  ( n93 ) & ( n26408 )  ;
assign n27700 =  ( n94 ) & ( n26378 )  ;
assign n27701 =  ( n94 ) & ( n26380 )  ;
assign n27702 =  ( n94 ) & ( n26382 )  ;
assign n27703 =  ( n94 ) & ( n26384 )  ;
assign n27704 =  ( n94 ) & ( n26386 )  ;
assign n27705 =  ( n94 ) & ( n26388 )  ;
assign n27706 =  ( n94 ) & ( n26390 )  ;
assign n27707 =  ( n94 ) & ( n26392 )  ;
assign n27708 =  ( n94 ) & ( n26394 )  ;
assign n27709 =  ( n94 ) & ( n26396 )  ;
assign n27710 =  ( n94 ) & ( n26398 )  ;
assign n27711 =  ( n94 ) & ( n26400 )  ;
assign n27712 =  ( n94 ) & ( n26402 )  ;
assign n27713 =  ( n94 ) & ( n26404 )  ;
assign n27714 =  ( n94 ) & ( n26406 )  ;
assign n27715 =  ( n94 ) & ( n26408 )  ;
assign n27716 =  ( n95 ) & ( n26378 )  ;
assign n27717 =  ( n95 ) & ( n26380 )  ;
assign n27718 =  ( n95 ) & ( n26382 )  ;
assign n27719 =  ( n95 ) & ( n26384 )  ;
assign n27720 =  ( n95 ) & ( n26386 )  ;
assign n27721 =  ( n95 ) & ( n26388 )  ;
assign n27722 =  ( n95 ) & ( n26390 )  ;
assign n27723 =  ( n95 ) & ( n26392 )  ;
assign n27724 =  ( n95 ) & ( n26394 )  ;
assign n27725 =  ( n95 ) & ( n26396 )  ;
assign n27726 =  ( n95 ) & ( n26398 )  ;
assign n27727 =  ( n95 ) & ( n26400 )  ;
assign n27728 =  ( n95 ) & ( n26402 )  ;
assign n27729 =  ( n95 ) & ( n26404 )  ;
assign n27730 =  ( n95 ) & ( n26406 )  ;
assign n27731 =  ( n95 ) & ( n26408 )  ;
assign n27732 =  ( n96 ) & ( n26378 )  ;
assign n27733 =  ( n96 ) & ( n26380 )  ;
assign n27734 =  ( n96 ) & ( n26382 )  ;
assign n27735 =  ( n96 ) & ( n26384 )  ;
assign n27736 =  ( n96 ) & ( n26386 )  ;
assign n27737 =  ( n96 ) & ( n26388 )  ;
assign n27738 =  ( n96 ) & ( n26390 )  ;
assign n27739 =  ( n96 ) & ( n26392 )  ;
assign n27740 =  ( n96 ) & ( n26394 )  ;
assign n27741 =  ( n96 ) & ( n26396 )  ;
assign n27742 =  ( n96 ) & ( n26398 )  ;
assign n27743 =  ( n96 ) & ( n26400 )  ;
assign n27744 =  ( n96 ) & ( n26402 )  ;
assign n27745 =  ( n96 ) & ( n26404 )  ;
assign n27746 =  ( n96 ) & ( n26406 )  ;
assign n27747 =  ( n96 ) & ( n26408 )  ;
assign n27748 =  ( n97 ) & ( n26378 )  ;
assign n27749 =  ( n97 ) & ( n26380 )  ;
assign n27750 =  ( n97 ) & ( n26382 )  ;
assign n27751 =  ( n97 ) & ( n26384 )  ;
assign n27752 =  ( n97 ) & ( n26386 )  ;
assign n27753 =  ( n97 ) & ( n26388 )  ;
assign n27754 =  ( n97 ) & ( n26390 )  ;
assign n27755 =  ( n97 ) & ( n26392 )  ;
assign n27756 =  ( n97 ) & ( n26394 )  ;
assign n27757 =  ( n97 ) & ( n26396 )  ;
assign n27758 =  ( n97 ) & ( n26398 )  ;
assign n27759 =  ( n97 ) & ( n26400 )  ;
assign n27760 =  ( n97 ) & ( n26402 )  ;
assign n27761 =  ( n97 ) & ( n26404 )  ;
assign n27762 =  ( n97 ) & ( n26406 )  ;
assign n27763 =  ( n97 ) & ( n26408 )  ;
assign n27764 =  ( n98 ) & ( n26378 )  ;
assign n27765 =  ( n98 ) & ( n26380 )  ;
assign n27766 =  ( n98 ) & ( n26382 )  ;
assign n27767 =  ( n98 ) & ( n26384 )  ;
assign n27768 =  ( n98 ) & ( n26386 )  ;
assign n27769 =  ( n98 ) & ( n26388 )  ;
assign n27770 =  ( n98 ) & ( n26390 )  ;
assign n27771 =  ( n98 ) & ( n26392 )  ;
assign n27772 =  ( n98 ) & ( n26394 )  ;
assign n27773 =  ( n98 ) & ( n26396 )  ;
assign n27774 =  ( n98 ) & ( n26398 )  ;
assign n27775 =  ( n98 ) & ( n26400 )  ;
assign n27776 =  ( n98 ) & ( n26402 )  ;
assign n27777 =  ( n98 ) & ( n26404 )  ;
assign n27778 =  ( n98 ) & ( n26406 )  ;
assign n27779 =  ( n98 ) & ( n26408 )  ;
assign n27780 =  ( n99 ) & ( n26378 )  ;
assign n27781 =  ( n99 ) & ( n26380 )  ;
assign n27782 =  ( n99 ) & ( n26382 )  ;
assign n27783 =  ( n99 ) & ( n26384 )  ;
assign n27784 =  ( n99 ) & ( n26386 )  ;
assign n27785 =  ( n99 ) & ( n26388 )  ;
assign n27786 =  ( n99 ) & ( n26390 )  ;
assign n27787 =  ( n99 ) & ( n26392 )  ;
assign n27788 =  ( n99 ) & ( n26394 )  ;
assign n27789 =  ( n99 ) & ( n26396 )  ;
assign n27790 =  ( n99 ) & ( n26398 )  ;
assign n27791 =  ( n99 ) & ( n26400 )  ;
assign n27792 =  ( n99 ) & ( n26402 )  ;
assign n27793 =  ( n99 ) & ( n26404 )  ;
assign n27794 =  ( n99 ) & ( n26406 )  ;
assign n27795 =  ( n99 ) & ( n26408 )  ;
assign n27796 =  ( n100 ) & ( n26378 )  ;
assign n27797 =  ( n100 ) & ( n26380 )  ;
assign n27798 =  ( n100 ) & ( n26382 )  ;
assign n27799 =  ( n100 ) & ( n26384 )  ;
assign n27800 =  ( n100 ) & ( n26386 )  ;
assign n27801 =  ( n100 ) & ( n26388 )  ;
assign n27802 =  ( n100 ) & ( n26390 )  ;
assign n27803 =  ( n100 ) & ( n26392 )  ;
assign n27804 =  ( n100 ) & ( n26394 )  ;
assign n27805 =  ( n100 ) & ( n26396 )  ;
assign n27806 =  ( n100 ) & ( n26398 )  ;
assign n27807 =  ( n100 ) & ( n26400 )  ;
assign n27808 =  ( n100 ) & ( n26402 )  ;
assign n27809 =  ( n100 ) & ( n26404 )  ;
assign n27810 =  ( n100 ) & ( n26406 )  ;
assign n27811 =  ( n100 ) & ( n26408 )  ;
assign n27812 =  ( n101 ) & ( n26378 )  ;
assign n27813 =  ( n101 ) & ( n26380 )  ;
assign n27814 =  ( n101 ) & ( n26382 )  ;
assign n27815 =  ( n101 ) & ( n26384 )  ;
assign n27816 =  ( n101 ) & ( n26386 )  ;
assign n27817 =  ( n101 ) & ( n26388 )  ;
assign n27818 =  ( n101 ) & ( n26390 )  ;
assign n27819 =  ( n101 ) & ( n26392 )  ;
assign n27820 =  ( n101 ) & ( n26394 )  ;
assign n27821 =  ( n101 ) & ( n26396 )  ;
assign n27822 =  ( n101 ) & ( n26398 )  ;
assign n27823 =  ( n101 ) & ( n26400 )  ;
assign n27824 =  ( n101 ) & ( n26402 )  ;
assign n27825 =  ( n101 ) & ( n26404 )  ;
assign n27826 =  ( n101 ) & ( n26406 )  ;
assign n27827 =  ( n101 ) & ( n26408 )  ;
assign n27828 =  ( n102 ) & ( n26378 )  ;
assign n27829 =  ( n102 ) & ( n26380 )  ;
assign n27830 =  ( n102 ) & ( n26382 )  ;
assign n27831 =  ( n102 ) & ( n26384 )  ;
assign n27832 =  ( n102 ) & ( n26386 )  ;
assign n27833 =  ( n102 ) & ( n26388 )  ;
assign n27834 =  ( n102 ) & ( n26390 )  ;
assign n27835 =  ( n102 ) & ( n26392 )  ;
assign n27836 =  ( n102 ) & ( n26394 )  ;
assign n27837 =  ( n102 ) & ( n26396 )  ;
assign n27838 =  ( n102 ) & ( n26398 )  ;
assign n27839 =  ( n102 ) & ( n26400 )  ;
assign n27840 =  ( n102 ) & ( n26402 )  ;
assign n27841 =  ( n102 ) & ( n26404 )  ;
assign n27842 =  ( n102 ) & ( n26406 )  ;
assign n27843 =  ( n102 ) & ( n26408 )  ;
assign n27844 =  ( n103 ) & ( n26378 )  ;
assign n27845 =  ( n103 ) & ( n26380 )  ;
assign n27846 =  ( n103 ) & ( n26382 )  ;
assign n27847 =  ( n103 ) & ( n26384 )  ;
assign n27848 =  ( n103 ) & ( n26386 )  ;
assign n27849 =  ( n103 ) & ( n26388 )  ;
assign n27850 =  ( n103 ) & ( n26390 )  ;
assign n27851 =  ( n103 ) & ( n26392 )  ;
assign n27852 =  ( n103 ) & ( n26394 )  ;
assign n27853 =  ( n103 ) & ( n26396 )  ;
assign n27854 =  ( n103 ) & ( n26398 )  ;
assign n27855 =  ( n103 ) & ( n26400 )  ;
assign n27856 =  ( n103 ) & ( n26402 )  ;
assign n27857 =  ( n103 ) & ( n26404 )  ;
assign n27858 =  ( n103 ) & ( n26406 )  ;
assign n27859 =  ( n103 ) & ( n26408 )  ;
assign n27860 =  ( n104 ) & ( n26378 )  ;
assign n27861 =  ( n104 ) & ( n26380 )  ;
assign n27862 =  ( n104 ) & ( n26382 )  ;
assign n27863 =  ( n104 ) & ( n26384 )  ;
assign n27864 =  ( n104 ) & ( n26386 )  ;
assign n27865 =  ( n104 ) & ( n26388 )  ;
assign n27866 =  ( n104 ) & ( n26390 )  ;
assign n27867 =  ( n104 ) & ( n26392 )  ;
assign n27868 =  ( n104 ) & ( n26394 )  ;
assign n27869 =  ( n104 ) & ( n26396 )  ;
assign n27870 =  ( n104 ) & ( n26398 )  ;
assign n27871 =  ( n104 ) & ( n26400 )  ;
assign n27872 =  ( n104 ) & ( n26402 )  ;
assign n27873 =  ( n104 ) & ( n26404 )  ;
assign n27874 =  ( n104 ) & ( n26406 )  ;
assign n27875 =  ( n104 ) & ( n26408 )  ;
assign n27876 =  ( n105 ) & ( n26378 )  ;
assign n27877 =  ( n105 ) & ( n26380 )  ;
assign n27878 =  ( n105 ) & ( n26382 )  ;
assign n27879 =  ( n105 ) & ( n26384 )  ;
assign n27880 =  ( n105 ) & ( n26386 )  ;
assign n27881 =  ( n105 ) & ( n26388 )  ;
assign n27882 =  ( n105 ) & ( n26390 )  ;
assign n27883 =  ( n105 ) & ( n26392 )  ;
assign n27884 =  ( n105 ) & ( n26394 )  ;
assign n27885 =  ( n105 ) & ( n26396 )  ;
assign n27886 =  ( n105 ) & ( n26398 )  ;
assign n27887 =  ( n105 ) & ( n26400 )  ;
assign n27888 =  ( n105 ) & ( n26402 )  ;
assign n27889 =  ( n105 ) & ( n26404 )  ;
assign n27890 =  ( n105 ) & ( n26406 )  ;
assign n27891 =  ( n105 ) & ( n26408 )  ;
assign n27892 =  ( n106 ) & ( n26378 )  ;
assign n27893 =  ( n106 ) & ( n26380 )  ;
assign n27894 =  ( n106 ) & ( n26382 )  ;
assign n27895 =  ( n106 ) & ( n26384 )  ;
assign n27896 =  ( n106 ) & ( n26386 )  ;
assign n27897 =  ( n106 ) & ( n26388 )  ;
assign n27898 =  ( n106 ) & ( n26390 )  ;
assign n27899 =  ( n106 ) & ( n26392 )  ;
assign n27900 =  ( n106 ) & ( n26394 )  ;
assign n27901 =  ( n106 ) & ( n26396 )  ;
assign n27902 =  ( n106 ) & ( n26398 )  ;
assign n27903 =  ( n106 ) & ( n26400 )  ;
assign n27904 =  ( n106 ) & ( n26402 )  ;
assign n27905 =  ( n106 ) & ( n26404 )  ;
assign n27906 =  ( n106 ) & ( n26406 )  ;
assign n27907 =  ( n106 ) & ( n26408 )  ;
assign n27908 =  ( n107 ) & ( n26378 )  ;
assign n27909 =  ( n107 ) & ( n26380 )  ;
assign n27910 =  ( n107 ) & ( n26382 )  ;
assign n27911 =  ( n107 ) & ( n26384 )  ;
assign n27912 =  ( n107 ) & ( n26386 )  ;
assign n27913 =  ( n107 ) & ( n26388 )  ;
assign n27914 =  ( n107 ) & ( n26390 )  ;
assign n27915 =  ( n107 ) & ( n26392 )  ;
assign n27916 =  ( n107 ) & ( n26394 )  ;
assign n27917 =  ( n107 ) & ( n26396 )  ;
assign n27918 =  ( n107 ) & ( n26398 )  ;
assign n27919 =  ( n107 ) & ( n26400 )  ;
assign n27920 =  ( n107 ) & ( n26402 )  ;
assign n27921 =  ( n107 ) & ( n26404 )  ;
assign n27922 =  ( n107 ) & ( n26406 )  ;
assign n27923 =  ( n107 ) & ( n26408 )  ;
assign n27924 =  ( n108 ) & ( n26378 )  ;
assign n27925 =  ( n108 ) & ( n26380 )  ;
assign n27926 =  ( n108 ) & ( n26382 )  ;
assign n27927 =  ( n108 ) & ( n26384 )  ;
assign n27928 =  ( n108 ) & ( n26386 )  ;
assign n27929 =  ( n108 ) & ( n26388 )  ;
assign n27930 =  ( n108 ) & ( n26390 )  ;
assign n27931 =  ( n108 ) & ( n26392 )  ;
assign n27932 =  ( n108 ) & ( n26394 )  ;
assign n27933 =  ( n108 ) & ( n26396 )  ;
assign n27934 =  ( n108 ) & ( n26398 )  ;
assign n27935 =  ( n108 ) & ( n26400 )  ;
assign n27936 =  ( n108 ) & ( n26402 )  ;
assign n27937 =  ( n108 ) & ( n26404 )  ;
assign n27938 =  ( n108 ) & ( n26406 )  ;
assign n27939 =  ( n108 ) & ( n26408 )  ;
assign n27940 =  ( n27939 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n27941 =  ( n27938 ) ? ( VREG_0_1 ) : ( n27940 ) ;
assign n27942 =  ( n27937 ) ? ( VREG_0_2 ) : ( n27941 ) ;
assign n27943 =  ( n27936 ) ? ( VREG_0_3 ) : ( n27942 ) ;
assign n27944 =  ( n27935 ) ? ( VREG_0_4 ) : ( n27943 ) ;
assign n27945 =  ( n27934 ) ? ( VREG_0_5 ) : ( n27944 ) ;
assign n27946 =  ( n27933 ) ? ( VREG_0_6 ) : ( n27945 ) ;
assign n27947 =  ( n27932 ) ? ( VREG_0_7 ) : ( n27946 ) ;
assign n27948 =  ( n27931 ) ? ( VREG_0_8 ) : ( n27947 ) ;
assign n27949 =  ( n27930 ) ? ( VREG_0_9 ) : ( n27948 ) ;
assign n27950 =  ( n27929 ) ? ( VREG_0_10 ) : ( n27949 ) ;
assign n27951 =  ( n27928 ) ? ( VREG_0_11 ) : ( n27950 ) ;
assign n27952 =  ( n27927 ) ? ( VREG_0_12 ) : ( n27951 ) ;
assign n27953 =  ( n27926 ) ? ( VREG_0_13 ) : ( n27952 ) ;
assign n27954 =  ( n27925 ) ? ( VREG_0_14 ) : ( n27953 ) ;
assign n27955 =  ( n27924 ) ? ( VREG_0_15 ) : ( n27954 ) ;
assign n27956 =  ( n27923 ) ? ( VREG_1_0 ) : ( n27955 ) ;
assign n27957 =  ( n27922 ) ? ( VREG_1_1 ) : ( n27956 ) ;
assign n27958 =  ( n27921 ) ? ( VREG_1_2 ) : ( n27957 ) ;
assign n27959 =  ( n27920 ) ? ( VREG_1_3 ) : ( n27958 ) ;
assign n27960 =  ( n27919 ) ? ( VREG_1_4 ) : ( n27959 ) ;
assign n27961 =  ( n27918 ) ? ( VREG_1_5 ) : ( n27960 ) ;
assign n27962 =  ( n27917 ) ? ( VREG_1_6 ) : ( n27961 ) ;
assign n27963 =  ( n27916 ) ? ( VREG_1_7 ) : ( n27962 ) ;
assign n27964 =  ( n27915 ) ? ( VREG_1_8 ) : ( n27963 ) ;
assign n27965 =  ( n27914 ) ? ( VREG_1_9 ) : ( n27964 ) ;
assign n27966 =  ( n27913 ) ? ( VREG_1_10 ) : ( n27965 ) ;
assign n27967 =  ( n27912 ) ? ( VREG_1_11 ) : ( n27966 ) ;
assign n27968 =  ( n27911 ) ? ( VREG_1_12 ) : ( n27967 ) ;
assign n27969 =  ( n27910 ) ? ( VREG_1_13 ) : ( n27968 ) ;
assign n27970 =  ( n27909 ) ? ( VREG_1_14 ) : ( n27969 ) ;
assign n27971 =  ( n27908 ) ? ( VREG_1_15 ) : ( n27970 ) ;
assign n27972 =  ( n27907 ) ? ( VREG_2_0 ) : ( n27971 ) ;
assign n27973 =  ( n27906 ) ? ( VREG_2_1 ) : ( n27972 ) ;
assign n27974 =  ( n27905 ) ? ( VREG_2_2 ) : ( n27973 ) ;
assign n27975 =  ( n27904 ) ? ( VREG_2_3 ) : ( n27974 ) ;
assign n27976 =  ( n27903 ) ? ( VREG_2_4 ) : ( n27975 ) ;
assign n27977 =  ( n27902 ) ? ( VREG_2_5 ) : ( n27976 ) ;
assign n27978 =  ( n27901 ) ? ( VREG_2_6 ) : ( n27977 ) ;
assign n27979 =  ( n27900 ) ? ( VREG_2_7 ) : ( n27978 ) ;
assign n27980 =  ( n27899 ) ? ( VREG_2_8 ) : ( n27979 ) ;
assign n27981 =  ( n27898 ) ? ( VREG_2_9 ) : ( n27980 ) ;
assign n27982 =  ( n27897 ) ? ( VREG_2_10 ) : ( n27981 ) ;
assign n27983 =  ( n27896 ) ? ( VREG_2_11 ) : ( n27982 ) ;
assign n27984 =  ( n27895 ) ? ( VREG_2_12 ) : ( n27983 ) ;
assign n27985 =  ( n27894 ) ? ( VREG_2_13 ) : ( n27984 ) ;
assign n27986 =  ( n27893 ) ? ( VREG_2_14 ) : ( n27985 ) ;
assign n27987 =  ( n27892 ) ? ( VREG_2_15 ) : ( n27986 ) ;
assign n27988 =  ( n27891 ) ? ( VREG_3_0 ) : ( n27987 ) ;
assign n27989 =  ( n27890 ) ? ( VREG_3_1 ) : ( n27988 ) ;
assign n27990 =  ( n27889 ) ? ( VREG_3_2 ) : ( n27989 ) ;
assign n27991 =  ( n27888 ) ? ( VREG_3_3 ) : ( n27990 ) ;
assign n27992 =  ( n27887 ) ? ( VREG_3_4 ) : ( n27991 ) ;
assign n27993 =  ( n27886 ) ? ( VREG_3_5 ) : ( n27992 ) ;
assign n27994 =  ( n27885 ) ? ( VREG_3_6 ) : ( n27993 ) ;
assign n27995 =  ( n27884 ) ? ( VREG_3_7 ) : ( n27994 ) ;
assign n27996 =  ( n27883 ) ? ( VREG_3_8 ) : ( n27995 ) ;
assign n27997 =  ( n27882 ) ? ( VREG_3_9 ) : ( n27996 ) ;
assign n27998 =  ( n27881 ) ? ( VREG_3_10 ) : ( n27997 ) ;
assign n27999 =  ( n27880 ) ? ( VREG_3_11 ) : ( n27998 ) ;
assign n28000 =  ( n27879 ) ? ( VREG_3_12 ) : ( n27999 ) ;
assign n28001 =  ( n27878 ) ? ( VREG_3_13 ) : ( n28000 ) ;
assign n28002 =  ( n27877 ) ? ( VREG_3_14 ) : ( n28001 ) ;
assign n28003 =  ( n27876 ) ? ( VREG_3_15 ) : ( n28002 ) ;
assign n28004 =  ( n27875 ) ? ( VREG_4_0 ) : ( n28003 ) ;
assign n28005 =  ( n27874 ) ? ( VREG_4_1 ) : ( n28004 ) ;
assign n28006 =  ( n27873 ) ? ( VREG_4_2 ) : ( n28005 ) ;
assign n28007 =  ( n27872 ) ? ( VREG_4_3 ) : ( n28006 ) ;
assign n28008 =  ( n27871 ) ? ( VREG_4_4 ) : ( n28007 ) ;
assign n28009 =  ( n27870 ) ? ( VREG_4_5 ) : ( n28008 ) ;
assign n28010 =  ( n27869 ) ? ( VREG_4_6 ) : ( n28009 ) ;
assign n28011 =  ( n27868 ) ? ( VREG_4_7 ) : ( n28010 ) ;
assign n28012 =  ( n27867 ) ? ( VREG_4_8 ) : ( n28011 ) ;
assign n28013 =  ( n27866 ) ? ( VREG_4_9 ) : ( n28012 ) ;
assign n28014 =  ( n27865 ) ? ( VREG_4_10 ) : ( n28013 ) ;
assign n28015 =  ( n27864 ) ? ( VREG_4_11 ) : ( n28014 ) ;
assign n28016 =  ( n27863 ) ? ( VREG_4_12 ) : ( n28015 ) ;
assign n28017 =  ( n27862 ) ? ( VREG_4_13 ) : ( n28016 ) ;
assign n28018 =  ( n27861 ) ? ( VREG_4_14 ) : ( n28017 ) ;
assign n28019 =  ( n27860 ) ? ( VREG_4_15 ) : ( n28018 ) ;
assign n28020 =  ( n27859 ) ? ( VREG_5_0 ) : ( n28019 ) ;
assign n28021 =  ( n27858 ) ? ( VREG_5_1 ) : ( n28020 ) ;
assign n28022 =  ( n27857 ) ? ( VREG_5_2 ) : ( n28021 ) ;
assign n28023 =  ( n27856 ) ? ( VREG_5_3 ) : ( n28022 ) ;
assign n28024 =  ( n27855 ) ? ( VREG_5_4 ) : ( n28023 ) ;
assign n28025 =  ( n27854 ) ? ( VREG_5_5 ) : ( n28024 ) ;
assign n28026 =  ( n27853 ) ? ( VREG_5_6 ) : ( n28025 ) ;
assign n28027 =  ( n27852 ) ? ( VREG_5_7 ) : ( n28026 ) ;
assign n28028 =  ( n27851 ) ? ( VREG_5_8 ) : ( n28027 ) ;
assign n28029 =  ( n27850 ) ? ( VREG_5_9 ) : ( n28028 ) ;
assign n28030 =  ( n27849 ) ? ( VREG_5_10 ) : ( n28029 ) ;
assign n28031 =  ( n27848 ) ? ( VREG_5_11 ) : ( n28030 ) ;
assign n28032 =  ( n27847 ) ? ( VREG_5_12 ) : ( n28031 ) ;
assign n28033 =  ( n27846 ) ? ( VREG_5_13 ) : ( n28032 ) ;
assign n28034 =  ( n27845 ) ? ( VREG_5_14 ) : ( n28033 ) ;
assign n28035 =  ( n27844 ) ? ( VREG_5_15 ) : ( n28034 ) ;
assign n28036 =  ( n27843 ) ? ( VREG_6_0 ) : ( n28035 ) ;
assign n28037 =  ( n27842 ) ? ( VREG_6_1 ) : ( n28036 ) ;
assign n28038 =  ( n27841 ) ? ( VREG_6_2 ) : ( n28037 ) ;
assign n28039 =  ( n27840 ) ? ( VREG_6_3 ) : ( n28038 ) ;
assign n28040 =  ( n27839 ) ? ( VREG_6_4 ) : ( n28039 ) ;
assign n28041 =  ( n27838 ) ? ( VREG_6_5 ) : ( n28040 ) ;
assign n28042 =  ( n27837 ) ? ( VREG_6_6 ) : ( n28041 ) ;
assign n28043 =  ( n27836 ) ? ( VREG_6_7 ) : ( n28042 ) ;
assign n28044 =  ( n27835 ) ? ( VREG_6_8 ) : ( n28043 ) ;
assign n28045 =  ( n27834 ) ? ( VREG_6_9 ) : ( n28044 ) ;
assign n28046 =  ( n27833 ) ? ( VREG_6_10 ) : ( n28045 ) ;
assign n28047 =  ( n27832 ) ? ( VREG_6_11 ) : ( n28046 ) ;
assign n28048 =  ( n27831 ) ? ( VREG_6_12 ) : ( n28047 ) ;
assign n28049 =  ( n27830 ) ? ( VREG_6_13 ) : ( n28048 ) ;
assign n28050 =  ( n27829 ) ? ( VREG_6_14 ) : ( n28049 ) ;
assign n28051 =  ( n27828 ) ? ( VREG_6_15 ) : ( n28050 ) ;
assign n28052 =  ( n27827 ) ? ( VREG_7_0 ) : ( n28051 ) ;
assign n28053 =  ( n27826 ) ? ( VREG_7_1 ) : ( n28052 ) ;
assign n28054 =  ( n27825 ) ? ( VREG_7_2 ) : ( n28053 ) ;
assign n28055 =  ( n27824 ) ? ( VREG_7_3 ) : ( n28054 ) ;
assign n28056 =  ( n27823 ) ? ( VREG_7_4 ) : ( n28055 ) ;
assign n28057 =  ( n27822 ) ? ( VREG_7_5 ) : ( n28056 ) ;
assign n28058 =  ( n27821 ) ? ( VREG_7_6 ) : ( n28057 ) ;
assign n28059 =  ( n27820 ) ? ( VREG_7_7 ) : ( n28058 ) ;
assign n28060 =  ( n27819 ) ? ( VREG_7_8 ) : ( n28059 ) ;
assign n28061 =  ( n27818 ) ? ( VREG_7_9 ) : ( n28060 ) ;
assign n28062 =  ( n27817 ) ? ( VREG_7_10 ) : ( n28061 ) ;
assign n28063 =  ( n27816 ) ? ( VREG_7_11 ) : ( n28062 ) ;
assign n28064 =  ( n27815 ) ? ( VREG_7_12 ) : ( n28063 ) ;
assign n28065 =  ( n27814 ) ? ( VREG_7_13 ) : ( n28064 ) ;
assign n28066 =  ( n27813 ) ? ( VREG_7_14 ) : ( n28065 ) ;
assign n28067 =  ( n27812 ) ? ( VREG_7_15 ) : ( n28066 ) ;
assign n28068 =  ( n27811 ) ? ( VREG_8_0 ) : ( n28067 ) ;
assign n28069 =  ( n27810 ) ? ( VREG_8_1 ) : ( n28068 ) ;
assign n28070 =  ( n27809 ) ? ( VREG_8_2 ) : ( n28069 ) ;
assign n28071 =  ( n27808 ) ? ( VREG_8_3 ) : ( n28070 ) ;
assign n28072 =  ( n27807 ) ? ( VREG_8_4 ) : ( n28071 ) ;
assign n28073 =  ( n27806 ) ? ( VREG_8_5 ) : ( n28072 ) ;
assign n28074 =  ( n27805 ) ? ( VREG_8_6 ) : ( n28073 ) ;
assign n28075 =  ( n27804 ) ? ( VREG_8_7 ) : ( n28074 ) ;
assign n28076 =  ( n27803 ) ? ( VREG_8_8 ) : ( n28075 ) ;
assign n28077 =  ( n27802 ) ? ( VREG_8_9 ) : ( n28076 ) ;
assign n28078 =  ( n27801 ) ? ( VREG_8_10 ) : ( n28077 ) ;
assign n28079 =  ( n27800 ) ? ( VREG_8_11 ) : ( n28078 ) ;
assign n28080 =  ( n27799 ) ? ( VREG_8_12 ) : ( n28079 ) ;
assign n28081 =  ( n27798 ) ? ( VREG_8_13 ) : ( n28080 ) ;
assign n28082 =  ( n27797 ) ? ( VREG_8_14 ) : ( n28081 ) ;
assign n28083 =  ( n27796 ) ? ( VREG_8_15 ) : ( n28082 ) ;
assign n28084 =  ( n27795 ) ? ( VREG_9_0 ) : ( n28083 ) ;
assign n28085 =  ( n27794 ) ? ( VREG_9_1 ) : ( n28084 ) ;
assign n28086 =  ( n27793 ) ? ( VREG_9_2 ) : ( n28085 ) ;
assign n28087 =  ( n27792 ) ? ( VREG_9_3 ) : ( n28086 ) ;
assign n28088 =  ( n27791 ) ? ( VREG_9_4 ) : ( n28087 ) ;
assign n28089 =  ( n27790 ) ? ( VREG_9_5 ) : ( n28088 ) ;
assign n28090 =  ( n27789 ) ? ( VREG_9_6 ) : ( n28089 ) ;
assign n28091 =  ( n27788 ) ? ( VREG_9_7 ) : ( n28090 ) ;
assign n28092 =  ( n27787 ) ? ( VREG_9_8 ) : ( n28091 ) ;
assign n28093 =  ( n27786 ) ? ( VREG_9_9 ) : ( n28092 ) ;
assign n28094 =  ( n27785 ) ? ( VREG_9_10 ) : ( n28093 ) ;
assign n28095 =  ( n27784 ) ? ( VREG_9_11 ) : ( n28094 ) ;
assign n28096 =  ( n27783 ) ? ( VREG_9_12 ) : ( n28095 ) ;
assign n28097 =  ( n27782 ) ? ( VREG_9_13 ) : ( n28096 ) ;
assign n28098 =  ( n27781 ) ? ( VREG_9_14 ) : ( n28097 ) ;
assign n28099 =  ( n27780 ) ? ( VREG_9_15 ) : ( n28098 ) ;
assign n28100 =  ( n27779 ) ? ( VREG_10_0 ) : ( n28099 ) ;
assign n28101 =  ( n27778 ) ? ( VREG_10_1 ) : ( n28100 ) ;
assign n28102 =  ( n27777 ) ? ( VREG_10_2 ) : ( n28101 ) ;
assign n28103 =  ( n27776 ) ? ( VREG_10_3 ) : ( n28102 ) ;
assign n28104 =  ( n27775 ) ? ( VREG_10_4 ) : ( n28103 ) ;
assign n28105 =  ( n27774 ) ? ( VREG_10_5 ) : ( n28104 ) ;
assign n28106 =  ( n27773 ) ? ( VREG_10_6 ) : ( n28105 ) ;
assign n28107 =  ( n27772 ) ? ( VREG_10_7 ) : ( n28106 ) ;
assign n28108 =  ( n27771 ) ? ( VREG_10_8 ) : ( n28107 ) ;
assign n28109 =  ( n27770 ) ? ( VREG_10_9 ) : ( n28108 ) ;
assign n28110 =  ( n27769 ) ? ( VREG_10_10 ) : ( n28109 ) ;
assign n28111 =  ( n27768 ) ? ( VREG_10_11 ) : ( n28110 ) ;
assign n28112 =  ( n27767 ) ? ( VREG_10_12 ) : ( n28111 ) ;
assign n28113 =  ( n27766 ) ? ( VREG_10_13 ) : ( n28112 ) ;
assign n28114 =  ( n27765 ) ? ( VREG_10_14 ) : ( n28113 ) ;
assign n28115 =  ( n27764 ) ? ( VREG_10_15 ) : ( n28114 ) ;
assign n28116 =  ( n27763 ) ? ( VREG_11_0 ) : ( n28115 ) ;
assign n28117 =  ( n27762 ) ? ( VREG_11_1 ) : ( n28116 ) ;
assign n28118 =  ( n27761 ) ? ( VREG_11_2 ) : ( n28117 ) ;
assign n28119 =  ( n27760 ) ? ( VREG_11_3 ) : ( n28118 ) ;
assign n28120 =  ( n27759 ) ? ( VREG_11_4 ) : ( n28119 ) ;
assign n28121 =  ( n27758 ) ? ( VREG_11_5 ) : ( n28120 ) ;
assign n28122 =  ( n27757 ) ? ( VREG_11_6 ) : ( n28121 ) ;
assign n28123 =  ( n27756 ) ? ( VREG_11_7 ) : ( n28122 ) ;
assign n28124 =  ( n27755 ) ? ( VREG_11_8 ) : ( n28123 ) ;
assign n28125 =  ( n27754 ) ? ( VREG_11_9 ) : ( n28124 ) ;
assign n28126 =  ( n27753 ) ? ( VREG_11_10 ) : ( n28125 ) ;
assign n28127 =  ( n27752 ) ? ( VREG_11_11 ) : ( n28126 ) ;
assign n28128 =  ( n27751 ) ? ( VREG_11_12 ) : ( n28127 ) ;
assign n28129 =  ( n27750 ) ? ( VREG_11_13 ) : ( n28128 ) ;
assign n28130 =  ( n27749 ) ? ( VREG_11_14 ) : ( n28129 ) ;
assign n28131 =  ( n27748 ) ? ( VREG_11_15 ) : ( n28130 ) ;
assign n28132 =  ( n27747 ) ? ( VREG_12_0 ) : ( n28131 ) ;
assign n28133 =  ( n27746 ) ? ( VREG_12_1 ) : ( n28132 ) ;
assign n28134 =  ( n27745 ) ? ( VREG_12_2 ) : ( n28133 ) ;
assign n28135 =  ( n27744 ) ? ( VREG_12_3 ) : ( n28134 ) ;
assign n28136 =  ( n27743 ) ? ( VREG_12_4 ) : ( n28135 ) ;
assign n28137 =  ( n27742 ) ? ( VREG_12_5 ) : ( n28136 ) ;
assign n28138 =  ( n27741 ) ? ( VREG_12_6 ) : ( n28137 ) ;
assign n28139 =  ( n27740 ) ? ( VREG_12_7 ) : ( n28138 ) ;
assign n28140 =  ( n27739 ) ? ( VREG_12_8 ) : ( n28139 ) ;
assign n28141 =  ( n27738 ) ? ( VREG_12_9 ) : ( n28140 ) ;
assign n28142 =  ( n27737 ) ? ( VREG_12_10 ) : ( n28141 ) ;
assign n28143 =  ( n27736 ) ? ( VREG_12_11 ) : ( n28142 ) ;
assign n28144 =  ( n27735 ) ? ( VREG_12_12 ) : ( n28143 ) ;
assign n28145 =  ( n27734 ) ? ( VREG_12_13 ) : ( n28144 ) ;
assign n28146 =  ( n27733 ) ? ( VREG_12_14 ) : ( n28145 ) ;
assign n28147 =  ( n27732 ) ? ( VREG_12_15 ) : ( n28146 ) ;
assign n28148 =  ( n27731 ) ? ( VREG_13_0 ) : ( n28147 ) ;
assign n28149 =  ( n27730 ) ? ( VREG_13_1 ) : ( n28148 ) ;
assign n28150 =  ( n27729 ) ? ( VREG_13_2 ) : ( n28149 ) ;
assign n28151 =  ( n27728 ) ? ( VREG_13_3 ) : ( n28150 ) ;
assign n28152 =  ( n27727 ) ? ( VREG_13_4 ) : ( n28151 ) ;
assign n28153 =  ( n27726 ) ? ( VREG_13_5 ) : ( n28152 ) ;
assign n28154 =  ( n27725 ) ? ( VREG_13_6 ) : ( n28153 ) ;
assign n28155 =  ( n27724 ) ? ( VREG_13_7 ) : ( n28154 ) ;
assign n28156 =  ( n27723 ) ? ( VREG_13_8 ) : ( n28155 ) ;
assign n28157 =  ( n27722 ) ? ( VREG_13_9 ) : ( n28156 ) ;
assign n28158 =  ( n27721 ) ? ( VREG_13_10 ) : ( n28157 ) ;
assign n28159 =  ( n27720 ) ? ( VREG_13_11 ) : ( n28158 ) ;
assign n28160 =  ( n27719 ) ? ( VREG_13_12 ) : ( n28159 ) ;
assign n28161 =  ( n27718 ) ? ( VREG_13_13 ) : ( n28160 ) ;
assign n28162 =  ( n27717 ) ? ( VREG_13_14 ) : ( n28161 ) ;
assign n28163 =  ( n27716 ) ? ( VREG_13_15 ) : ( n28162 ) ;
assign n28164 =  ( n27715 ) ? ( VREG_14_0 ) : ( n28163 ) ;
assign n28165 =  ( n27714 ) ? ( VREG_14_1 ) : ( n28164 ) ;
assign n28166 =  ( n27713 ) ? ( VREG_14_2 ) : ( n28165 ) ;
assign n28167 =  ( n27712 ) ? ( VREG_14_3 ) : ( n28166 ) ;
assign n28168 =  ( n27711 ) ? ( VREG_14_4 ) : ( n28167 ) ;
assign n28169 =  ( n27710 ) ? ( VREG_14_5 ) : ( n28168 ) ;
assign n28170 =  ( n27709 ) ? ( VREG_14_6 ) : ( n28169 ) ;
assign n28171 =  ( n27708 ) ? ( VREG_14_7 ) : ( n28170 ) ;
assign n28172 =  ( n27707 ) ? ( VREG_14_8 ) : ( n28171 ) ;
assign n28173 =  ( n27706 ) ? ( VREG_14_9 ) : ( n28172 ) ;
assign n28174 =  ( n27705 ) ? ( VREG_14_10 ) : ( n28173 ) ;
assign n28175 =  ( n27704 ) ? ( VREG_14_11 ) : ( n28174 ) ;
assign n28176 =  ( n27703 ) ? ( VREG_14_12 ) : ( n28175 ) ;
assign n28177 =  ( n27702 ) ? ( VREG_14_13 ) : ( n28176 ) ;
assign n28178 =  ( n27701 ) ? ( VREG_14_14 ) : ( n28177 ) ;
assign n28179 =  ( n27700 ) ? ( VREG_14_15 ) : ( n28178 ) ;
assign n28180 =  ( n27699 ) ? ( VREG_15_0 ) : ( n28179 ) ;
assign n28181 =  ( n27698 ) ? ( VREG_15_1 ) : ( n28180 ) ;
assign n28182 =  ( n27697 ) ? ( VREG_15_2 ) : ( n28181 ) ;
assign n28183 =  ( n27696 ) ? ( VREG_15_3 ) : ( n28182 ) ;
assign n28184 =  ( n27695 ) ? ( VREG_15_4 ) : ( n28183 ) ;
assign n28185 =  ( n27694 ) ? ( VREG_15_5 ) : ( n28184 ) ;
assign n28186 =  ( n27693 ) ? ( VREG_15_6 ) : ( n28185 ) ;
assign n28187 =  ( n27692 ) ? ( VREG_15_7 ) : ( n28186 ) ;
assign n28188 =  ( n27691 ) ? ( VREG_15_8 ) : ( n28187 ) ;
assign n28189 =  ( n27690 ) ? ( VREG_15_9 ) : ( n28188 ) ;
assign n28190 =  ( n27689 ) ? ( VREG_15_10 ) : ( n28189 ) ;
assign n28191 =  ( n27688 ) ? ( VREG_15_11 ) : ( n28190 ) ;
assign n28192 =  ( n27687 ) ? ( VREG_15_12 ) : ( n28191 ) ;
assign n28193 =  ( n27686 ) ? ( VREG_15_13 ) : ( n28192 ) ;
assign n28194 =  ( n27685 ) ? ( VREG_15_14 ) : ( n28193 ) ;
assign n28195 =  ( n27684 ) ? ( VREG_15_15 ) : ( n28194 ) ;
assign n28196 =  ( n27683 ) ? ( VREG_16_0 ) : ( n28195 ) ;
assign n28197 =  ( n27682 ) ? ( VREG_16_1 ) : ( n28196 ) ;
assign n28198 =  ( n27681 ) ? ( VREG_16_2 ) : ( n28197 ) ;
assign n28199 =  ( n27680 ) ? ( VREG_16_3 ) : ( n28198 ) ;
assign n28200 =  ( n27679 ) ? ( VREG_16_4 ) : ( n28199 ) ;
assign n28201 =  ( n27678 ) ? ( VREG_16_5 ) : ( n28200 ) ;
assign n28202 =  ( n27677 ) ? ( VREG_16_6 ) : ( n28201 ) ;
assign n28203 =  ( n27676 ) ? ( VREG_16_7 ) : ( n28202 ) ;
assign n28204 =  ( n27675 ) ? ( VREG_16_8 ) : ( n28203 ) ;
assign n28205 =  ( n27674 ) ? ( VREG_16_9 ) : ( n28204 ) ;
assign n28206 =  ( n27673 ) ? ( VREG_16_10 ) : ( n28205 ) ;
assign n28207 =  ( n27672 ) ? ( VREG_16_11 ) : ( n28206 ) ;
assign n28208 =  ( n27671 ) ? ( VREG_16_12 ) : ( n28207 ) ;
assign n28209 =  ( n27670 ) ? ( VREG_16_13 ) : ( n28208 ) ;
assign n28210 =  ( n27669 ) ? ( VREG_16_14 ) : ( n28209 ) ;
assign n28211 =  ( n27668 ) ? ( VREG_16_15 ) : ( n28210 ) ;
assign n28212 =  ( n27667 ) ? ( VREG_17_0 ) : ( n28211 ) ;
assign n28213 =  ( n27666 ) ? ( VREG_17_1 ) : ( n28212 ) ;
assign n28214 =  ( n27665 ) ? ( VREG_17_2 ) : ( n28213 ) ;
assign n28215 =  ( n27664 ) ? ( VREG_17_3 ) : ( n28214 ) ;
assign n28216 =  ( n27663 ) ? ( VREG_17_4 ) : ( n28215 ) ;
assign n28217 =  ( n27662 ) ? ( VREG_17_5 ) : ( n28216 ) ;
assign n28218 =  ( n27661 ) ? ( VREG_17_6 ) : ( n28217 ) ;
assign n28219 =  ( n27660 ) ? ( VREG_17_7 ) : ( n28218 ) ;
assign n28220 =  ( n27659 ) ? ( VREG_17_8 ) : ( n28219 ) ;
assign n28221 =  ( n27658 ) ? ( VREG_17_9 ) : ( n28220 ) ;
assign n28222 =  ( n27657 ) ? ( VREG_17_10 ) : ( n28221 ) ;
assign n28223 =  ( n27656 ) ? ( VREG_17_11 ) : ( n28222 ) ;
assign n28224 =  ( n27655 ) ? ( VREG_17_12 ) : ( n28223 ) ;
assign n28225 =  ( n27654 ) ? ( VREG_17_13 ) : ( n28224 ) ;
assign n28226 =  ( n27653 ) ? ( VREG_17_14 ) : ( n28225 ) ;
assign n28227 =  ( n27652 ) ? ( VREG_17_15 ) : ( n28226 ) ;
assign n28228 =  ( n27651 ) ? ( VREG_18_0 ) : ( n28227 ) ;
assign n28229 =  ( n27650 ) ? ( VREG_18_1 ) : ( n28228 ) ;
assign n28230 =  ( n27649 ) ? ( VREG_18_2 ) : ( n28229 ) ;
assign n28231 =  ( n27648 ) ? ( VREG_18_3 ) : ( n28230 ) ;
assign n28232 =  ( n27647 ) ? ( VREG_18_4 ) : ( n28231 ) ;
assign n28233 =  ( n27646 ) ? ( VREG_18_5 ) : ( n28232 ) ;
assign n28234 =  ( n27645 ) ? ( VREG_18_6 ) : ( n28233 ) ;
assign n28235 =  ( n27644 ) ? ( VREG_18_7 ) : ( n28234 ) ;
assign n28236 =  ( n27643 ) ? ( VREG_18_8 ) : ( n28235 ) ;
assign n28237 =  ( n27642 ) ? ( VREG_18_9 ) : ( n28236 ) ;
assign n28238 =  ( n27641 ) ? ( VREG_18_10 ) : ( n28237 ) ;
assign n28239 =  ( n27640 ) ? ( VREG_18_11 ) : ( n28238 ) ;
assign n28240 =  ( n27639 ) ? ( VREG_18_12 ) : ( n28239 ) ;
assign n28241 =  ( n27638 ) ? ( VREG_18_13 ) : ( n28240 ) ;
assign n28242 =  ( n27637 ) ? ( VREG_18_14 ) : ( n28241 ) ;
assign n28243 =  ( n27636 ) ? ( VREG_18_15 ) : ( n28242 ) ;
assign n28244 =  ( n27635 ) ? ( VREG_19_0 ) : ( n28243 ) ;
assign n28245 =  ( n27634 ) ? ( VREG_19_1 ) : ( n28244 ) ;
assign n28246 =  ( n27633 ) ? ( VREG_19_2 ) : ( n28245 ) ;
assign n28247 =  ( n27632 ) ? ( VREG_19_3 ) : ( n28246 ) ;
assign n28248 =  ( n27631 ) ? ( VREG_19_4 ) : ( n28247 ) ;
assign n28249 =  ( n27630 ) ? ( VREG_19_5 ) : ( n28248 ) ;
assign n28250 =  ( n27629 ) ? ( VREG_19_6 ) : ( n28249 ) ;
assign n28251 =  ( n27628 ) ? ( VREG_19_7 ) : ( n28250 ) ;
assign n28252 =  ( n27627 ) ? ( VREG_19_8 ) : ( n28251 ) ;
assign n28253 =  ( n27626 ) ? ( VREG_19_9 ) : ( n28252 ) ;
assign n28254 =  ( n27625 ) ? ( VREG_19_10 ) : ( n28253 ) ;
assign n28255 =  ( n27624 ) ? ( VREG_19_11 ) : ( n28254 ) ;
assign n28256 =  ( n27623 ) ? ( VREG_19_12 ) : ( n28255 ) ;
assign n28257 =  ( n27622 ) ? ( VREG_19_13 ) : ( n28256 ) ;
assign n28258 =  ( n27621 ) ? ( VREG_19_14 ) : ( n28257 ) ;
assign n28259 =  ( n27620 ) ? ( VREG_19_15 ) : ( n28258 ) ;
assign n28260 =  ( n27619 ) ? ( VREG_20_0 ) : ( n28259 ) ;
assign n28261 =  ( n27618 ) ? ( VREG_20_1 ) : ( n28260 ) ;
assign n28262 =  ( n27617 ) ? ( VREG_20_2 ) : ( n28261 ) ;
assign n28263 =  ( n27616 ) ? ( VREG_20_3 ) : ( n28262 ) ;
assign n28264 =  ( n27615 ) ? ( VREG_20_4 ) : ( n28263 ) ;
assign n28265 =  ( n27614 ) ? ( VREG_20_5 ) : ( n28264 ) ;
assign n28266 =  ( n27613 ) ? ( VREG_20_6 ) : ( n28265 ) ;
assign n28267 =  ( n27612 ) ? ( VREG_20_7 ) : ( n28266 ) ;
assign n28268 =  ( n27611 ) ? ( VREG_20_8 ) : ( n28267 ) ;
assign n28269 =  ( n27610 ) ? ( VREG_20_9 ) : ( n28268 ) ;
assign n28270 =  ( n27609 ) ? ( VREG_20_10 ) : ( n28269 ) ;
assign n28271 =  ( n27608 ) ? ( VREG_20_11 ) : ( n28270 ) ;
assign n28272 =  ( n27607 ) ? ( VREG_20_12 ) : ( n28271 ) ;
assign n28273 =  ( n27606 ) ? ( VREG_20_13 ) : ( n28272 ) ;
assign n28274 =  ( n27605 ) ? ( VREG_20_14 ) : ( n28273 ) ;
assign n28275 =  ( n27604 ) ? ( VREG_20_15 ) : ( n28274 ) ;
assign n28276 =  ( n27603 ) ? ( VREG_21_0 ) : ( n28275 ) ;
assign n28277 =  ( n27602 ) ? ( VREG_21_1 ) : ( n28276 ) ;
assign n28278 =  ( n27601 ) ? ( VREG_21_2 ) : ( n28277 ) ;
assign n28279 =  ( n27600 ) ? ( VREG_21_3 ) : ( n28278 ) ;
assign n28280 =  ( n27599 ) ? ( VREG_21_4 ) : ( n28279 ) ;
assign n28281 =  ( n27598 ) ? ( VREG_21_5 ) : ( n28280 ) ;
assign n28282 =  ( n27597 ) ? ( VREG_21_6 ) : ( n28281 ) ;
assign n28283 =  ( n27596 ) ? ( VREG_21_7 ) : ( n28282 ) ;
assign n28284 =  ( n27595 ) ? ( VREG_21_8 ) : ( n28283 ) ;
assign n28285 =  ( n27594 ) ? ( VREG_21_9 ) : ( n28284 ) ;
assign n28286 =  ( n27593 ) ? ( VREG_21_10 ) : ( n28285 ) ;
assign n28287 =  ( n27592 ) ? ( VREG_21_11 ) : ( n28286 ) ;
assign n28288 =  ( n27591 ) ? ( VREG_21_12 ) : ( n28287 ) ;
assign n28289 =  ( n27590 ) ? ( VREG_21_13 ) : ( n28288 ) ;
assign n28290 =  ( n27589 ) ? ( VREG_21_14 ) : ( n28289 ) ;
assign n28291 =  ( n27588 ) ? ( VREG_21_15 ) : ( n28290 ) ;
assign n28292 =  ( n27587 ) ? ( VREG_22_0 ) : ( n28291 ) ;
assign n28293 =  ( n27586 ) ? ( VREG_22_1 ) : ( n28292 ) ;
assign n28294 =  ( n27585 ) ? ( VREG_22_2 ) : ( n28293 ) ;
assign n28295 =  ( n27584 ) ? ( VREG_22_3 ) : ( n28294 ) ;
assign n28296 =  ( n27583 ) ? ( VREG_22_4 ) : ( n28295 ) ;
assign n28297 =  ( n27582 ) ? ( VREG_22_5 ) : ( n28296 ) ;
assign n28298 =  ( n27581 ) ? ( VREG_22_6 ) : ( n28297 ) ;
assign n28299 =  ( n27580 ) ? ( VREG_22_7 ) : ( n28298 ) ;
assign n28300 =  ( n27579 ) ? ( VREG_22_8 ) : ( n28299 ) ;
assign n28301 =  ( n27578 ) ? ( VREG_22_9 ) : ( n28300 ) ;
assign n28302 =  ( n27577 ) ? ( VREG_22_10 ) : ( n28301 ) ;
assign n28303 =  ( n27576 ) ? ( VREG_22_11 ) : ( n28302 ) ;
assign n28304 =  ( n27575 ) ? ( VREG_22_12 ) : ( n28303 ) ;
assign n28305 =  ( n27574 ) ? ( VREG_22_13 ) : ( n28304 ) ;
assign n28306 =  ( n27573 ) ? ( VREG_22_14 ) : ( n28305 ) ;
assign n28307 =  ( n27572 ) ? ( VREG_22_15 ) : ( n28306 ) ;
assign n28308 =  ( n27571 ) ? ( VREG_23_0 ) : ( n28307 ) ;
assign n28309 =  ( n27570 ) ? ( VREG_23_1 ) : ( n28308 ) ;
assign n28310 =  ( n27569 ) ? ( VREG_23_2 ) : ( n28309 ) ;
assign n28311 =  ( n27568 ) ? ( VREG_23_3 ) : ( n28310 ) ;
assign n28312 =  ( n27567 ) ? ( VREG_23_4 ) : ( n28311 ) ;
assign n28313 =  ( n27566 ) ? ( VREG_23_5 ) : ( n28312 ) ;
assign n28314 =  ( n27565 ) ? ( VREG_23_6 ) : ( n28313 ) ;
assign n28315 =  ( n27564 ) ? ( VREG_23_7 ) : ( n28314 ) ;
assign n28316 =  ( n27563 ) ? ( VREG_23_8 ) : ( n28315 ) ;
assign n28317 =  ( n27562 ) ? ( VREG_23_9 ) : ( n28316 ) ;
assign n28318 =  ( n27561 ) ? ( VREG_23_10 ) : ( n28317 ) ;
assign n28319 =  ( n27560 ) ? ( VREG_23_11 ) : ( n28318 ) ;
assign n28320 =  ( n27559 ) ? ( VREG_23_12 ) : ( n28319 ) ;
assign n28321 =  ( n27558 ) ? ( VREG_23_13 ) : ( n28320 ) ;
assign n28322 =  ( n27557 ) ? ( VREG_23_14 ) : ( n28321 ) ;
assign n28323 =  ( n27556 ) ? ( VREG_23_15 ) : ( n28322 ) ;
assign n28324 =  ( n27555 ) ? ( VREG_24_0 ) : ( n28323 ) ;
assign n28325 =  ( n27554 ) ? ( VREG_24_1 ) : ( n28324 ) ;
assign n28326 =  ( n27553 ) ? ( VREG_24_2 ) : ( n28325 ) ;
assign n28327 =  ( n27552 ) ? ( VREG_24_3 ) : ( n28326 ) ;
assign n28328 =  ( n27551 ) ? ( VREG_24_4 ) : ( n28327 ) ;
assign n28329 =  ( n27550 ) ? ( VREG_24_5 ) : ( n28328 ) ;
assign n28330 =  ( n27549 ) ? ( VREG_24_6 ) : ( n28329 ) ;
assign n28331 =  ( n27548 ) ? ( VREG_24_7 ) : ( n28330 ) ;
assign n28332 =  ( n27547 ) ? ( VREG_24_8 ) : ( n28331 ) ;
assign n28333 =  ( n27546 ) ? ( VREG_24_9 ) : ( n28332 ) ;
assign n28334 =  ( n27545 ) ? ( VREG_24_10 ) : ( n28333 ) ;
assign n28335 =  ( n27544 ) ? ( VREG_24_11 ) : ( n28334 ) ;
assign n28336 =  ( n27543 ) ? ( VREG_24_12 ) : ( n28335 ) ;
assign n28337 =  ( n27542 ) ? ( VREG_24_13 ) : ( n28336 ) ;
assign n28338 =  ( n27541 ) ? ( VREG_24_14 ) : ( n28337 ) ;
assign n28339 =  ( n27540 ) ? ( VREG_24_15 ) : ( n28338 ) ;
assign n28340 =  ( n27539 ) ? ( VREG_25_0 ) : ( n28339 ) ;
assign n28341 =  ( n27538 ) ? ( VREG_25_1 ) : ( n28340 ) ;
assign n28342 =  ( n27537 ) ? ( VREG_25_2 ) : ( n28341 ) ;
assign n28343 =  ( n27536 ) ? ( VREG_25_3 ) : ( n28342 ) ;
assign n28344 =  ( n27535 ) ? ( VREG_25_4 ) : ( n28343 ) ;
assign n28345 =  ( n27534 ) ? ( VREG_25_5 ) : ( n28344 ) ;
assign n28346 =  ( n27533 ) ? ( VREG_25_6 ) : ( n28345 ) ;
assign n28347 =  ( n27532 ) ? ( VREG_25_7 ) : ( n28346 ) ;
assign n28348 =  ( n27531 ) ? ( VREG_25_8 ) : ( n28347 ) ;
assign n28349 =  ( n27530 ) ? ( VREG_25_9 ) : ( n28348 ) ;
assign n28350 =  ( n27529 ) ? ( VREG_25_10 ) : ( n28349 ) ;
assign n28351 =  ( n27528 ) ? ( VREG_25_11 ) : ( n28350 ) ;
assign n28352 =  ( n27527 ) ? ( VREG_25_12 ) : ( n28351 ) ;
assign n28353 =  ( n27526 ) ? ( VREG_25_13 ) : ( n28352 ) ;
assign n28354 =  ( n27525 ) ? ( VREG_25_14 ) : ( n28353 ) ;
assign n28355 =  ( n27524 ) ? ( VREG_25_15 ) : ( n28354 ) ;
assign n28356 =  ( n27523 ) ? ( VREG_26_0 ) : ( n28355 ) ;
assign n28357 =  ( n27522 ) ? ( VREG_26_1 ) : ( n28356 ) ;
assign n28358 =  ( n27521 ) ? ( VREG_26_2 ) : ( n28357 ) ;
assign n28359 =  ( n27520 ) ? ( VREG_26_3 ) : ( n28358 ) ;
assign n28360 =  ( n27519 ) ? ( VREG_26_4 ) : ( n28359 ) ;
assign n28361 =  ( n27518 ) ? ( VREG_26_5 ) : ( n28360 ) ;
assign n28362 =  ( n27517 ) ? ( VREG_26_6 ) : ( n28361 ) ;
assign n28363 =  ( n27516 ) ? ( VREG_26_7 ) : ( n28362 ) ;
assign n28364 =  ( n27515 ) ? ( VREG_26_8 ) : ( n28363 ) ;
assign n28365 =  ( n27514 ) ? ( VREG_26_9 ) : ( n28364 ) ;
assign n28366 =  ( n27513 ) ? ( VREG_26_10 ) : ( n28365 ) ;
assign n28367 =  ( n27512 ) ? ( VREG_26_11 ) : ( n28366 ) ;
assign n28368 =  ( n27511 ) ? ( VREG_26_12 ) : ( n28367 ) ;
assign n28369 =  ( n27510 ) ? ( VREG_26_13 ) : ( n28368 ) ;
assign n28370 =  ( n27509 ) ? ( VREG_26_14 ) : ( n28369 ) ;
assign n28371 =  ( n27508 ) ? ( VREG_26_15 ) : ( n28370 ) ;
assign n28372 =  ( n27507 ) ? ( VREG_27_0 ) : ( n28371 ) ;
assign n28373 =  ( n27506 ) ? ( VREG_27_1 ) : ( n28372 ) ;
assign n28374 =  ( n27505 ) ? ( VREG_27_2 ) : ( n28373 ) ;
assign n28375 =  ( n27504 ) ? ( VREG_27_3 ) : ( n28374 ) ;
assign n28376 =  ( n27503 ) ? ( VREG_27_4 ) : ( n28375 ) ;
assign n28377 =  ( n27502 ) ? ( VREG_27_5 ) : ( n28376 ) ;
assign n28378 =  ( n27501 ) ? ( VREG_27_6 ) : ( n28377 ) ;
assign n28379 =  ( n27500 ) ? ( VREG_27_7 ) : ( n28378 ) ;
assign n28380 =  ( n27499 ) ? ( VREG_27_8 ) : ( n28379 ) ;
assign n28381 =  ( n27498 ) ? ( VREG_27_9 ) : ( n28380 ) ;
assign n28382 =  ( n27497 ) ? ( VREG_27_10 ) : ( n28381 ) ;
assign n28383 =  ( n27496 ) ? ( VREG_27_11 ) : ( n28382 ) ;
assign n28384 =  ( n27495 ) ? ( VREG_27_12 ) : ( n28383 ) ;
assign n28385 =  ( n27494 ) ? ( VREG_27_13 ) : ( n28384 ) ;
assign n28386 =  ( n27493 ) ? ( VREG_27_14 ) : ( n28385 ) ;
assign n28387 =  ( n27492 ) ? ( VREG_27_15 ) : ( n28386 ) ;
assign n28388 =  ( n27491 ) ? ( VREG_28_0 ) : ( n28387 ) ;
assign n28389 =  ( n27490 ) ? ( VREG_28_1 ) : ( n28388 ) ;
assign n28390 =  ( n27489 ) ? ( VREG_28_2 ) : ( n28389 ) ;
assign n28391 =  ( n27488 ) ? ( VREG_28_3 ) : ( n28390 ) ;
assign n28392 =  ( n27487 ) ? ( VREG_28_4 ) : ( n28391 ) ;
assign n28393 =  ( n27486 ) ? ( VREG_28_5 ) : ( n28392 ) ;
assign n28394 =  ( n27485 ) ? ( VREG_28_6 ) : ( n28393 ) ;
assign n28395 =  ( n27484 ) ? ( VREG_28_7 ) : ( n28394 ) ;
assign n28396 =  ( n27483 ) ? ( VREG_28_8 ) : ( n28395 ) ;
assign n28397 =  ( n27482 ) ? ( VREG_28_9 ) : ( n28396 ) ;
assign n28398 =  ( n27481 ) ? ( VREG_28_10 ) : ( n28397 ) ;
assign n28399 =  ( n27480 ) ? ( VREG_28_11 ) : ( n28398 ) ;
assign n28400 =  ( n27479 ) ? ( VREG_28_12 ) : ( n28399 ) ;
assign n28401 =  ( n27478 ) ? ( VREG_28_13 ) : ( n28400 ) ;
assign n28402 =  ( n27477 ) ? ( VREG_28_14 ) : ( n28401 ) ;
assign n28403 =  ( n27476 ) ? ( VREG_28_15 ) : ( n28402 ) ;
assign n28404 =  ( n27475 ) ? ( VREG_29_0 ) : ( n28403 ) ;
assign n28405 =  ( n27474 ) ? ( VREG_29_1 ) : ( n28404 ) ;
assign n28406 =  ( n27473 ) ? ( VREG_29_2 ) : ( n28405 ) ;
assign n28407 =  ( n27472 ) ? ( VREG_29_3 ) : ( n28406 ) ;
assign n28408 =  ( n27471 ) ? ( VREG_29_4 ) : ( n28407 ) ;
assign n28409 =  ( n27470 ) ? ( VREG_29_5 ) : ( n28408 ) ;
assign n28410 =  ( n27469 ) ? ( VREG_29_6 ) : ( n28409 ) ;
assign n28411 =  ( n27468 ) ? ( VREG_29_7 ) : ( n28410 ) ;
assign n28412 =  ( n27467 ) ? ( VREG_29_8 ) : ( n28411 ) ;
assign n28413 =  ( n27466 ) ? ( VREG_29_9 ) : ( n28412 ) ;
assign n28414 =  ( n27465 ) ? ( VREG_29_10 ) : ( n28413 ) ;
assign n28415 =  ( n27464 ) ? ( VREG_29_11 ) : ( n28414 ) ;
assign n28416 =  ( n27463 ) ? ( VREG_29_12 ) : ( n28415 ) ;
assign n28417 =  ( n27462 ) ? ( VREG_29_13 ) : ( n28416 ) ;
assign n28418 =  ( n27461 ) ? ( VREG_29_14 ) : ( n28417 ) ;
assign n28419 =  ( n27460 ) ? ( VREG_29_15 ) : ( n28418 ) ;
assign n28420 =  ( n27459 ) ? ( VREG_30_0 ) : ( n28419 ) ;
assign n28421 =  ( n27458 ) ? ( VREG_30_1 ) : ( n28420 ) ;
assign n28422 =  ( n27457 ) ? ( VREG_30_2 ) : ( n28421 ) ;
assign n28423 =  ( n27456 ) ? ( VREG_30_3 ) : ( n28422 ) ;
assign n28424 =  ( n27455 ) ? ( VREG_30_4 ) : ( n28423 ) ;
assign n28425 =  ( n27454 ) ? ( VREG_30_5 ) : ( n28424 ) ;
assign n28426 =  ( n27453 ) ? ( VREG_30_6 ) : ( n28425 ) ;
assign n28427 =  ( n27452 ) ? ( VREG_30_7 ) : ( n28426 ) ;
assign n28428 =  ( n27451 ) ? ( VREG_30_8 ) : ( n28427 ) ;
assign n28429 =  ( n27450 ) ? ( VREG_30_9 ) : ( n28428 ) ;
assign n28430 =  ( n27449 ) ? ( VREG_30_10 ) : ( n28429 ) ;
assign n28431 =  ( n27448 ) ? ( VREG_30_11 ) : ( n28430 ) ;
assign n28432 =  ( n27447 ) ? ( VREG_30_12 ) : ( n28431 ) ;
assign n28433 =  ( n27446 ) ? ( VREG_30_13 ) : ( n28432 ) ;
assign n28434 =  ( n27445 ) ? ( VREG_30_14 ) : ( n28433 ) ;
assign n28435 =  ( n27444 ) ? ( VREG_30_15 ) : ( n28434 ) ;
assign n28436 =  ( n27443 ) ? ( VREG_31_0 ) : ( n28435 ) ;
assign n28437 =  ( n27442 ) ? ( VREG_31_1 ) : ( n28436 ) ;
assign n28438 =  ( n27441 ) ? ( VREG_31_2 ) : ( n28437 ) ;
assign n28439 =  ( n27440 ) ? ( VREG_31_3 ) : ( n28438 ) ;
assign n28440 =  ( n27439 ) ? ( VREG_31_4 ) : ( n28439 ) ;
assign n28441 =  ( n27438 ) ? ( VREG_31_5 ) : ( n28440 ) ;
assign n28442 =  ( n27437 ) ? ( VREG_31_6 ) : ( n28441 ) ;
assign n28443 =  ( n27436 ) ? ( VREG_31_7 ) : ( n28442 ) ;
assign n28444 =  ( n27435 ) ? ( VREG_31_8 ) : ( n28443 ) ;
assign n28445 =  ( n27434 ) ? ( VREG_31_9 ) : ( n28444 ) ;
assign n28446 =  ( n27433 ) ? ( VREG_31_10 ) : ( n28445 ) ;
assign n28447 =  ( n27432 ) ? ( VREG_31_11 ) : ( n28446 ) ;
assign n28448 =  ( n27431 ) ? ( VREG_31_12 ) : ( n28447 ) ;
assign n28449 =  ( n27430 ) ? ( VREG_31_13 ) : ( n28448 ) ;
assign n28450 =  ( n27429 ) ? ( VREG_31_14 ) : ( n28449 ) ;
assign n28451 =  ( n27428 ) ? ( VREG_31_15 ) : ( n28450 ) ;
assign n28452 =  ( n27417 ) + ( n28451 )  ;
assign n28453 =  ( n27417 ) - ( n28451 )  ;
assign n28454 =  ( n27417 ) & ( n28451 )  ;
assign n28455 =  ( n27417 ) | ( n28451 )  ;
assign n28456 =  ( ( n27417 ) * ( n28451 ))  ;
assign n28457 =  ( n148 ) ? ( n28456 ) : ( VREG_0_6 ) ;
assign n28458 =  ( n146 ) ? ( n28455 ) : ( n28457 ) ;
assign n28459 =  ( n144 ) ? ( n28454 ) : ( n28458 ) ;
assign n28460 =  ( n142 ) ? ( n28453 ) : ( n28459 ) ;
assign n28461 =  ( n10 ) ? ( n28452 ) : ( n28460 ) ;
assign n28462 = n3030[6:6] ;
assign n28463 =  ( n28462 ) == ( 1'd0 )  ;
assign n28464 =  ( n28463 ) ? ( VREG_0_6 ) : ( n27427 ) ;
assign n28465 =  ( n28463 ) ? ( VREG_0_6 ) : ( n28461 ) ;
assign n28466 =  ( n3034 ) ? ( n28465 ) : ( VREG_0_6 ) ;
assign n28467 =  ( n2965 ) ? ( n28464 ) : ( n28466 ) ;
assign n28468 =  ( n1930 ) ? ( n28461 ) : ( n28467 ) ;
assign n28469 =  ( n879 ) ? ( n27427 ) : ( n28468 ) ;
assign n28470 =  ( n27417 ) + ( n164 )  ;
assign n28471 =  ( n27417 ) - ( n164 )  ;
assign n28472 =  ( n27417 ) & ( n164 )  ;
assign n28473 =  ( n27417 ) | ( n164 )  ;
assign n28474 =  ( ( n27417 ) * ( n164 ))  ;
assign n28475 =  ( n172 ) ? ( n28474 ) : ( VREG_0_6 ) ;
assign n28476 =  ( n170 ) ? ( n28473 ) : ( n28475 ) ;
assign n28477 =  ( n168 ) ? ( n28472 ) : ( n28476 ) ;
assign n28478 =  ( n166 ) ? ( n28471 ) : ( n28477 ) ;
assign n28479 =  ( n162 ) ? ( n28470 ) : ( n28478 ) ;
assign n28480 =  ( n27417 ) + ( n180 )  ;
assign n28481 =  ( n27417 ) - ( n180 )  ;
assign n28482 =  ( n27417 ) & ( n180 )  ;
assign n28483 =  ( n27417 ) | ( n180 )  ;
assign n28484 =  ( ( n27417 ) * ( n180 ))  ;
assign n28485 =  ( n172 ) ? ( n28484 ) : ( VREG_0_6 ) ;
assign n28486 =  ( n170 ) ? ( n28483 ) : ( n28485 ) ;
assign n28487 =  ( n168 ) ? ( n28482 ) : ( n28486 ) ;
assign n28488 =  ( n166 ) ? ( n28481 ) : ( n28487 ) ;
assign n28489 =  ( n162 ) ? ( n28480 ) : ( n28488 ) ;
assign n28490 =  ( n28463 ) ? ( VREG_0_6 ) : ( n28489 ) ;
assign n28491 =  ( n3051 ) ? ( n28490 ) : ( VREG_0_6 ) ;
assign n28492 =  ( n3040 ) ? ( n28479 ) : ( n28491 ) ;
assign n28493 =  ( n192 ) ? ( VREG_0_6 ) : ( VREG_0_6 ) ;
assign n28494 =  ( n157 ) ? ( n28492 ) : ( n28493 ) ;
assign n28495 =  ( n6 ) ? ( n28469 ) : ( n28494 ) ;
assign n28496 =  ( n4 ) ? ( n28495 ) : ( VREG_0_6 ) ;
assign n28497 =  ( 32'd7 ) == ( 32'd15 )  ;
assign n28498 =  ( n12 ) & ( n28497 )  ;
assign n28499 =  ( 32'd7 ) == ( 32'd14 )  ;
assign n28500 =  ( n12 ) & ( n28499 )  ;
assign n28501 =  ( 32'd7 ) == ( 32'd13 )  ;
assign n28502 =  ( n12 ) & ( n28501 )  ;
assign n28503 =  ( 32'd7 ) == ( 32'd12 )  ;
assign n28504 =  ( n12 ) & ( n28503 )  ;
assign n28505 =  ( 32'd7 ) == ( 32'd11 )  ;
assign n28506 =  ( n12 ) & ( n28505 )  ;
assign n28507 =  ( 32'd7 ) == ( 32'd10 )  ;
assign n28508 =  ( n12 ) & ( n28507 )  ;
assign n28509 =  ( 32'd7 ) == ( 32'd9 )  ;
assign n28510 =  ( n12 ) & ( n28509 )  ;
assign n28511 =  ( 32'd7 ) == ( 32'd8 )  ;
assign n28512 =  ( n12 ) & ( n28511 )  ;
assign n28513 =  ( 32'd7 ) == ( 32'd7 )  ;
assign n28514 =  ( n12 ) & ( n28513 )  ;
assign n28515 =  ( 32'd7 ) == ( 32'd6 )  ;
assign n28516 =  ( n12 ) & ( n28515 )  ;
assign n28517 =  ( 32'd7 ) == ( 32'd5 )  ;
assign n28518 =  ( n12 ) & ( n28517 )  ;
assign n28519 =  ( 32'd7 ) == ( 32'd4 )  ;
assign n28520 =  ( n12 ) & ( n28519 )  ;
assign n28521 =  ( 32'd7 ) == ( 32'd3 )  ;
assign n28522 =  ( n12 ) & ( n28521 )  ;
assign n28523 =  ( 32'd7 ) == ( 32'd2 )  ;
assign n28524 =  ( n12 ) & ( n28523 )  ;
assign n28525 =  ( 32'd7 ) == ( 32'd1 )  ;
assign n28526 =  ( n12 ) & ( n28525 )  ;
assign n28527 =  ( 32'd7 ) == ( 32'd0 )  ;
assign n28528 =  ( n12 ) & ( n28527 )  ;
assign n28529 =  ( n13 ) & ( n28497 )  ;
assign n28530 =  ( n13 ) & ( n28499 )  ;
assign n28531 =  ( n13 ) & ( n28501 )  ;
assign n28532 =  ( n13 ) & ( n28503 )  ;
assign n28533 =  ( n13 ) & ( n28505 )  ;
assign n28534 =  ( n13 ) & ( n28507 )  ;
assign n28535 =  ( n13 ) & ( n28509 )  ;
assign n28536 =  ( n13 ) & ( n28511 )  ;
assign n28537 =  ( n13 ) & ( n28513 )  ;
assign n28538 =  ( n13 ) & ( n28515 )  ;
assign n28539 =  ( n13 ) & ( n28517 )  ;
assign n28540 =  ( n13 ) & ( n28519 )  ;
assign n28541 =  ( n13 ) & ( n28521 )  ;
assign n28542 =  ( n13 ) & ( n28523 )  ;
assign n28543 =  ( n13 ) & ( n28525 )  ;
assign n28544 =  ( n13 ) & ( n28527 )  ;
assign n28545 =  ( n14 ) & ( n28497 )  ;
assign n28546 =  ( n14 ) & ( n28499 )  ;
assign n28547 =  ( n14 ) & ( n28501 )  ;
assign n28548 =  ( n14 ) & ( n28503 )  ;
assign n28549 =  ( n14 ) & ( n28505 )  ;
assign n28550 =  ( n14 ) & ( n28507 )  ;
assign n28551 =  ( n14 ) & ( n28509 )  ;
assign n28552 =  ( n14 ) & ( n28511 )  ;
assign n28553 =  ( n14 ) & ( n28513 )  ;
assign n28554 =  ( n14 ) & ( n28515 )  ;
assign n28555 =  ( n14 ) & ( n28517 )  ;
assign n28556 =  ( n14 ) & ( n28519 )  ;
assign n28557 =  ( n14 ) & ( n28521 )  ;
assign n28558 =  ( n14 ) & ( n28523 )  ;
assign n28559 =  ( n14 ) & ( n28525 )  ;
assign n28560 =  ( n14 ) & ( n28527 )  ;
assign n28561 =  ( n15 ) & ( n28497 )  ;
assign n28562 =  ( n15 ) & ( n28499 )  ;
assign n28563 =  ( n15 ) & ( n28501 )  ;
assign n28564 =  ( n15 ) & ( n28503 )  ;
assign n28565 =  ( n15 ) & ( n28505 )  ;
assign n28566 =  ( n15 ) & ( n28507 )  ;
assign n28567 =  ( n15 ) & ( n28509 )  ;
assign n28568 =  ( n15 ) & ( n28511 )  ;
assign n28569 =  ( n15 ) & ( n28513 )  ;
assign n28570 =  ( n15 ) & ( n28515 )  ;
assign n28571 =  ( n15 ) & ( n28517 )  ;
assign n28572 =  ( n15 ) & ( n28519 )  ;
assign n28573 =  ( n15 ) & ( n28521 )  ;
assign n28574 =  ( n15 ) & ( n28523 )  ;
assign n28575 =  ( n15 ) & ( n28525 )  ;
assign n28576 =  ( n15 ) & ( n28527 )  ;
assign n28577 =  ( n16 ) & ( n28497 )  ;
assign n28578 =  ( n16 ) & ( n28499 )  ;
assign n28579 =  ( n16 ) & ( n28501 )  ;
assign n28580 =  ( n16 ) & ( n28503 )  ;
assign n28581 =  ( n16 ) & ( n28505 )  ;
assign n28582 =  ( n16 ) & ( n28507 )  ;
assign n28583 =  ( n16 ) & ( n28509 )  ;
assign n28584 =  ( n16 ) & ( n28511 )  ;
assign n28585 =  ( n16 ) & ( n28513 )  ;
assign n28586 =  ( n16 ) & ( n28515 )  ;
assign n28587 =  ( n16 ) & ( n28517 )  ;
assign n28588 =  ( n16 ) & ( n28519 )  ;
assign n28589 =  ( n16 ) & ( n28521 )  ;
assign n28590 =  ( n16 ) & ( n28523 )  ;
assign n28591 =  ( n16 ) & ( n28525 )  ;
assign n28592 =  ( n16 ) & ( n28527 )  ;
assign n28593 =  ( n17 ) & ( n28497 )  ;
assign n28594 =  ( n17 ) & ( n28499 )  ;
assign n28595 =  ( n17 ) & ( n28501 )  ;
assign n28596 =  ( n17 ) & ( n28503 )  ;
assign n28597 =  ( n17 ) & ( n28505 )  ;
assign n28598 =  ( n17 ) & ( n28507 )  ;
assign n28599 =  ( n17 ) & ( n28509 )  ;
assign n28600 =  ( n17 ) & ( n28511 )  ;
assign n28601 =  ( n17 ) & ( n28513 )  ;
assign n28602 =  ( n17 ) & ( n28515 )  ;
assign n28603 =  ( n17 ) & ( n28517 )  ;
assign n28604 =  ( n17 ) & ( n28519 )  ;
assign n28605 =  ( n17 ) & ( n28521 )  ;
assign n28606 =  ( n17 ) & ( n28523 )  ;
assign n28607 =  ( n17 ) & ( n28525 )  ;
assign n28608 =  ( n17 ) & ( n28527 )  ;
assign n28609 =  ( n18 ) & ( n28497 )  ;
assign n28610 =  ( n18 ) & ( n28499 )  ;
assign n28611 =  ( n18 ) & ( n28501 )  ;
assign n28612 =  ( n18 ) & ( n28503 )  ;
assign n28613 =  ( n18 ) & ( n28505 )  ;
assign n28614 =  ( n18 ) & ( n28507 )  ;
assign n28615 =  ( n18 ) & ( n28509 )  ;
assign n28616 =  ( n18 ) & ( n28511 )  ;
assign n28617 =  ( n18 ) & ( n28513 )  ;
assign n28618 =  ( n18 ) & ( n28515 )  ;
assign n28619 =  ( n18 ) & ( n28517 )  ;
assign n28620 =  ( n18 ) & ( n28519 )  ;
assign n28621 =  ( n18 ) & ( n28521 )  ;
assign n28622 =  ( n18 ) & ( n28523 )  ;
assign n28623 =  ( n18 ) & ( n28525 )  ;
assign n28624 =  ( n18 ) & ( n28527 )  ;
assign n28625 =  ( n19 ) & ( n28497 )  ;
assign n28626 =  ( n19 ) & ( n28499 )  ;
assign n28627 =  ( n19 ) & ( n28501 )  ;
assign n28628 =  ( n19 ) & ( n28503 )  ;
assign n28629 =  ( n19 ) & ( n28505 )  ;
assign n28630 =  ( n19 ) & ( n28507 )  ;
assign n28631 =  ( n19 ) & ( n28509 )  ;
assign n28632 =  ( n19 ) & ( n28511 )  ;
assign n28633 =  ( n19 ) & ( n28513 )  ;
assign n28634 =  ( n19 ) & ( n28515 )  ;
assign n28635 =  ( n19 ) & ( n28517 )  ;
assign n28636 =  ( n19 ) & ( n28519 )  ;
assign n28637 =  ( n19 ) & ( n28521 )  ;
assign n28638 =  ( n19 ) & ( n28523 )  ;
assign n28639 =  ( n19 ) & ( n28525 )  ;
assign n28640 =  ( n19 ) & ( n28527 )  ;
assign n28641 =  ( n20 ) & ( n28497 )  ;
assign n28642 =  ( n20 ) & ( n28499 )  ;
assign n28643 =  ( n20 ) & ( n28501 )  ;
assign n28644 =  ( n20 ) & ( n28503 )  ;
assign n28645 =  ( n20 ) & ( n28505 )  ;
assign n28646 =  ( n20 ) & ( n28507 )  ;
assign n28647 =  ( n20 ) & ( n28509 )  ;
assign n28648 =  ( n20 ) & ( n28511 )  ;
assign n28649 =  ( n20 ) & ( n28513 )  ;
assign n28650 =  ( n20 ) & ( n28515 )  ;
assign n28651 =  ( n20 ) & ( n28517 )  ;
assign n28652 =  ( n20 ) & ( n28519 )  ;
assign n28653 =  ( n20 ) & ( n28521 )  ;
assign n28654 =  ( n20 ) & ( n28523 )  ;
assign n28655 =  ( n20 ) & ( n28525 )  ;
assign n28656 =  ( n20 ) & ( n28527 )  ;
assign n28657 =  ( n21 ) & ( n28497 )  ;
assign n28658 =  ( n21 ) & ( n28499 )  ;
assign n28659 =  ( n21 ) & ( n28501 )  ;
assign n28660 =  ( n21 ) & ( n28503 )  ;
assign n28661 =  ( n21 ) & ( n28505 )  ;
assign n28662 =  ( n21 ) & ( n28507 )  ;
assign n28663 =  ( n21 ) & ( n28509 )  ;
assign n28664 =  ( n21 ) & ( n28511 )  ;
assign n28665 =  ( n21 ) & ( n28513 )  ;
assign n28666 =  ( n21 ) & ( n28515 )  ;
assign n28667 =  ( n21 ) & ( n28517 )  ;
assign n28668 =  ( n21 ) & ( n28519 )  ;
assign n28669 =  ( n21 ) & ( n28521 )  ;
assign n28670 =  ( n21 ) & ( n28523 )  ;
assign n28671 =  ( n21 ) & ( n28525 )  ;
assign n28672 =  ( n21 ) & ( n28527 )  ;
assign n28673 =  ( n22 ) & ( n28497 )  ;
assign n28674 =  ( n22 ) & ( n28499 )  ;
assign n28675 =  ( n22 ) & ( n28501 )  ;
assign n28676 =  ( n22 ) & ( n28503 )  ;
assign n28677 =  ( n22 ) & ( n28505 )  ;
assign n28678 =  ( n22 ) & ( n28507 )  ;
assign n28679 =  ( n22 ) & ( n28509 )  ;
assign n28680 =  ( n22 ) & ( n28511 )  ;
assign n28681 =  ( n22 ) & ( n28513 )  ;
assign n28682 =  ( n22 ) & ( n28515 )  ;
assign n28683 =  ( n22 ) & ( n28517 )  ;
assign n28684 =  ( n22 ) & ( n28519 )  ;
assign n28685 =  ( n22 ) & ( n28521 )  ;
assign n28686 =  ( n22 ) & ( n28523 )  ;
assign n28687 =  ( n22 ) & ( n28525 )  ;
assign n28688 =  ( n22 ) & ( n28527 )  ;
assign n28689 =  ( n23 ) & ( n28497 )  ;
assign n28690 =  ( n23 ) & ( n28499 )  ;
assign n28691 =  ( n23 ) & ( n28501 )  ;
assign n28692 =  ( n23 ) & ( n28503 )  ;
assign n28693 =  ( n23 ) & ( n28505 )  ;
assign n28694 =  ( n23 ) & ( n28507 )  ;
assign n28695 =  ( n23 ) & ( n28509 )  ;
assign n28696 =  ( n23 ) & ( n28511 )  ;
assign n28697 =  ( n23 ) & ( n28513 )  ;
assign n28698 =  ( n23 ) & ( n28515 )  ;
assign n28699 =  ( n23 ) & ( n28517 )  ;
assign n28700 =  ( n23 ) & ( n28519 )  ;
assign n28701 =  ( n23 ) & ( n28521 )  ;
assign n28702 =  ( n23 ) & ( n28523 )  ;
assign n28703 =  ( n23 ) & ( n28525 )  ;
assign n28704 =  ( n23 ) & ( n28527 )  ;
assign n28705 =  ( n24 ) & ( n28497 )  ;
assign n28706 =  ( n24 ) & ( n28499 )  ;
assign n28707 =  ( n24 ) & ( n28501 )  ;
assign n28708 =  ( n24 ) & ( n28503 )  ;
assign n28709 =  ( n24 ) & ( n28505 )  ;
assign n28710 =  ( n24 ) & ( n28507 )  ;
assign n28711 =  ( n24 ) & ( n28509 )  ;
assign n28712 =  ( n24 ) & ( n28511 )  ;
assign n28713 =  ( n24 ) & ( n28513 )  ;
assign n28714 =  ( n24 ) & ( n28515 )  ;
assign n28715 =  ( n24 ) & ( n28517 )  ;
assign n28716 =  ( n24 ) & ( n28519 )  ;
assign n28717 =  ( n24 ) & ( n28521 )  ;
assign n28718 =  ( n24 ) & ( n28523 )  ;
assign n28719 =  ( n24 ) & ( n28525 )  ;
assign n28720 =  ( n24 ) & ( n28527 )  ;
assign n28721 =  ( n25 ) & ( n28497 )  ;
assign n28722 =  ( n25 ) & ( n28499 )  ;
assign n28723 =  ( n25 ) & ( n28501 )  ;
assign n28724 =  ( n25 ) & ( n28503 )  ;
assign n28725 =  ( n25 ) & ( n28505 )  ;
assign n28726 =  ( n25 ) & ( n28507 )  ;
assign n28727 =  ( n25 ) & ( n28509 )  ;
assign n28728 =  ( n25 ) & ( n28511 )  ;
assign n28729 =  ( n25 ) & ( n28513 )  ;
assign n28730 =  ( n25 ) & ( n28515 )  ;
assign n28731 =  ( n25 ) & ( n28517 )  ;
assign n28732 =  ( n25 ) & ( n28519 )  ;
assign n28733 =  ( n25 ) & ( n28521 )  ;
assign n28734 =  ( n25 ) & ( n28523 )  ;
assign n28735 =  ( n25 ) & ( n28525 )  ;
assign n28736 =  ( n25 ) & ( n28527 )  ;
assign n28737 =  ( n26 ) & ( n28497 )  ;
assign n28738 =  ( n26 ) & ( n28499 )  ;
assign n28739 =  ( n26 ) & ( n28501 )  ;
assign n28740 =  ( n26 ) & ( n28503 )  ;
assign n28741 =  ( n26 ) & ( n28505 )  ;
assign n28742 =  ( n26 ) & ( n28507 )  ;
assign n28743 =  ( n26 ) & ( n28509 )  ;
assign n28744 =  ( n26 ) & ( n28511 )  ;
assign n28745 =  ( n26 ) & ( n28513 )  ;
assign n28746 =  ( n26 ) & ( n28515 )  ;
assign n28747 =  ( n26 ) & ( n28517 )  ;
assign n28748 =  ( n26 ) & ( n28519 )  ;
assign n28749 =  ( n26 ) & ( n28521 )  ;
assign n28750 =  ( n26 ) & ( n28523 )  ;
assign n28751 =  ( n26 ) & ( n28525 )  ;
assign n28752 =  ( n26 ) & ( n28527 )  ;
assign n28753 =  ( n27 ) & ( n28497 )  ;
assign n28754 =  ( n27 ) & ( n28499 )  ;
assign n28755 =  ( n27 ) & ( n28501 )  ;
assign n28756 =  ( n27 ) & ( n28503 )  ;
assign n28757 =  ( n27 ) & ( n28505 )  ;
assign n28758 =  ( n27 ) & ( n28507 )  ;
assign n28759 =  ( n27 ) & ( n28509 )  ;
assign n28760 =  ( n27 ) & ( n28511 )  ;
assign n28761 =  ( n27 ) & ( n28513 )  ;
assign n28762 =  ( n27 ) & ( n28515 )  ;
assign n28763 =  ( n27 ) & ( n28517 )  ;
assign n28764 =  ( n27 ) & ( n28519 )  ;
assign n28765 =  ( n27 ) & ( n28521 )  ;
assign n28766 =  ( n27 ) & ( n28523 )  ;
assign n28767 =  ( n27 ) & ( n28525 )  ;
assign n28768 =  ( n27 ) & ( n28527 )  ;
assign n28769 =  ( n28 ) & ( n28497 )  ;
assign n28770 =  ( n28 ) & ( n28499 )  ;
assign n28771 =  ( n28 ) & ( n28501 )  ;
assign n28772 =  ( n28 ) & ( n28503 )  ;
assign n28773 =  ( n28 ) & ( n28505 )  ;
assign n28774 =  ( n28 ) & ( n28507 )  ;
assign n28775 =  ( n28 ) & ( n28509 )  ;
assign n28776 =  ( n28 ) & ( n28511 )  ;
assign n28777 =  ( n28 ) & ( n28513 )  ;
assign n28778 =  ( n28 ) & ( n28515 )  ;
assign n28779 =  ( n28 ) & ( n28517 )  ;
assign n28780 =  ( n28 ) & ( n28519 )  ;
assign n28781 =  ( n28 ) & ( n28521 )  ;
assign n28782 =  ( n28 ) & ( n28523 )  ;
assign n28783 =  ( n28 ) & ( n28525 )  ;
assign n28784 =  ( n28 ) & ( n28527 )  ;
assign n28785 =  ( n29 ) & ( n28497 )  ;
assign n28786 =  ( n29 ) & ( n28499 )  ;
assign n28787 =  ( n29 ) & ( n28501 )  ;
assign n28788 =  ( n29 ) & ( n28503 )  ;
assign n28789 =  ( n29 ) & ( n28505 )  ;
assign n28790 =  ( n29 ) & ( n28507 )  ;
assign n28791 =  ( n29 ) & ( n28509 )  ;
assign n28792 =  ( n29 ) & ( n28511 )  ;
assign n28793 =  ( n29 ) & ( n28513 )  ;
assign n28794 =  ( n29 ) & ( n28515 )  ;
assign n28795 =  ( n29 ) & ( n28517 )  ;
assign n28796 =  ( n29 ) & ( n28519 )  ;
assign n28797 =  ( n29 ) & ( n28521 )  ;
assign n28798 =  ( n29 ) & ( n28523 )  ;
assign n28799 =  ( n29 ) & ( n28525 )  ;
assign n28800 =  ( n29 ) & ( n28527 )  ;
assign n28801 =  ( n30 ) & ( n28497 )  ;
assign n28802 =  ( n30 ) & ( n28499 )  ;
assign n28803 =  ( n30 ) & ( n28501 )  ;
assign n28804 =  ( n30 ) & ( n28503 )  ;
assign n28805 =  ( n30 ) & ( n28505 )  ;
assign n28806 =  ( n30 ) & ( n28507 )  ;
assign n28807 =  ( n30 ) & ( n28509 )  ;
assign n28808 =  ( n30 ) & ( n28511 )  ;
assign n28809 =  ( n30 ) & ( n28513 )  ;
assign n28810 =  ( n30 ) & ( n28515 )  ;
assign n28811 =  ( n30 ) & ( n28517 )  ;
assign n28812 =  ( n30 ) & ( n28519 )  ;
assign n28813 =  ( n30 ) & ( n28521 )  ;
assign n28814 =  ( n30 ) & ( n28523 )  ;
assign n28815 =  ( n30 ) & ( n28525 )  ;
assign n28816 =  ( n30 ) & ( n28527 )  ;
assign n28817 =  ( n31 ) & ( n28497 )  ;
assign n28818 =  ( n31 ) & ( n28499 )  ;
assign n28819 =  ( n31 ) & ( n28501 )  ;
assign n28820 =  ( n31 ) & ( n28503 )  ;
assign n28821 =  ( n31 ) & ( n28505 )  ;
assign n28822 =  ( n31 ) & ( n28507 )  ;
assign n28823 =  ( n31 ) & ( n28509 )  ;
assign n28824 =  ( n31 ) & ( n28511 )  ;
assign n28825 =  ( n31 ) & ( n28513 )  ;
assign n28826 =  ( n31 ) & ( n28515 )  ;
assign n28827 =  ( n31 ) & ( n28517 )  ;
assign n28828 =  ( n31 ) & ( n28519 )  ;
assign n28829 =  ( n31 ) & ( n28521 )  ;
assign n28830 =  ( n31 ) & ( n28523 )  ;
assign n28831 =  ( n31 ) & ( n28525 )  ;
assign n28832 =  ( n31 ) & ( n28527 )  ;
assign n28833 =  ( n32 ) & ( n28497 )  ;
assign n28834 =  ( n32 ) & ( n28499 )  ;
assign n28835 =  ( n32 ) & ( n28501 )  ;
assign n28836 =  ( n32 ) & ( n28503 )  ;
assign n28837 =  ( n32 ) & ( n28505 )  ;
assign n28838 =  ( n32 ) & ( n28507 )  ;
assign n28839 =  ( n32 ) & ( n28509 )  ;
assign n28840 =  ( n32 ) & ( n28511 )  ;
assign n28841 =  ( n32 ) & ( n28513 )  ;
assign n28842 =  ( n32 ) & ( n28515 )  ;
assign n28843 =  ( n32 ) & ( n28517 )  ;
assign n28844 =  ( n32 ) & ( n28519 )  ;
assign n28845 =  ( n32 ) & ( n28521 )  ;
assign n28846 =  ( n32 ) & ( n28523 )  ;
assign n28847 =  ( n32 ) & ( n28525 )  ;
assign n28848 =  ( n32 ) & ( n28527 )  ;
assign n28849 =  ( n33 ) & ( n28497 )  ;
assign n28850 =  ( n33 ) & ( n28499 )  ;
assign n28851 =  ( n33 ) & ( n28501 )  ;
assign n28852 =  ( n33 ) & ( n28503 )  ;
assign n28853 =  ( n33 ) & ( n28505 )  ;
assign n28854 =  ( n33 ) & ( n28507 )  ;
assign n28855 =  ( n33 ) & ( n28509 )  ;
assign n28856 =  ( n33 ) & ( n28511 )  ;
assign n28857 =  ( n33 ) & ( n28513 )  ;
assign n28858 =  ( n33 ) & ( n28515 )  ;
assign n28859 =  ( n33 ) & ( n28517 )  ;
assign n28860 =  ( n33 ) & ( n28519 )  ;
assign n28861 =  ( n33 ) & ( n28521 )  ;
assign n28862 =  ( n33 ) & ( n28523 )  ;
assign n28863 =  ( n33 ) & ( n28525 )  ;
assign n28864 =  ( n33 ) & ( n28527 )  ;
assign n28865 =  ( n34 ) & ( n28497 )  ;
assign n28866 =  ( n34 ) & ( n28499 )  ;
assign n28867 =  ( n34 ) & ( n28501 )  ;
assign n28868 =  ( n34 ) & ( n28503 )  ;
assign n28869 =  ( n34 ) & ( n28505 )  ;
assign n28870 =  ( n34 ) & ( n28507 )  ;
assign n28871 =  ( n34 ) & ( n28509 )  ;
assign n28872 =  ( n34 ) & ( n28511 )  ;
assign n28873 =  ( n34 ) & ( n28513 )  ;
assign n28874 =  ( n34 ) & ( n28515 )  ;
assign n28875 =  ( n34 ) & ( n28517 )  ;
assign n28876 =  ( n34 ) & ( n28519 )  ;
assign n28877 =  ( n34 ) & ( n28521 )  ;
assign n28878 =  ( n34 ) & ( n28523 )  ;
assign n28879 =  ( n34 ) & ( n28525 )  ;
assign n28880 =  ( n34 ) & ( n28527 )  ;
assign n28881 =  ( n35 ) & ( n28497 )  ;
assign n28882 =  ( n35 ) & ( n28499 )  ;
assign n28883 =  ( n35 ) & ( n28501 )  ;
assign n28884 =  ( n35 ) & ( n28503 )  ;
assign n28885 =  ( n35 ) & ( n28505 )  ;
assign n28886 =  ( n35 ) & ( n28507 )  ;
assign n28887 =  ( n35 ) & ( n28509 )  ;
assign n28888 =  ( n35 ) & ( n28511 )  ;
assign n28889 =  ( n35 ) & ( n28513 )  ;
assign n28890 =  ( n35 ) & ( n28515 )  ;
assign n28891 =  ( n35 ) & ( n28517 )  ;
assign n28892 =  ( n35 ) & ( n28519 )  ;
assign n28893 =  ( n35 ) & ( n28521 )  ;
assign n28894 =  ( n35 ) & ( n28523 )  ;
assign n28895 =  ( n35 ) & ( n28525 )  ;
assign n28896 =  ( n35 ) & ( n28527 )  ;
assign n28897 =  ( n36 ) & ( n28497 )  ;
assign n28898 =  ( n36 ) & ( n28499 )  ;
assign n28899 =  ( n36 ) & ( n28501 )  ;
assign n28900 =  ( n36 ) & ( n28503 )  ;
assign n28901 =  ( n36 ) & ( n28505 )  ;
assign n28902 =  ( n36 ) & ( n28507 )  ;
assign n28903 =  ( n36 ) & ( n28509 )  ;
assign n28904 =  ( n36 ) & ( n28511 )  ;
assign n28905 =  ( n36 ) & ( n28513 )  ;
assign n28906 =  ( n36 ) & ( n28515 )  ;
assign n28907 =  ( n36 ) & ( n28517 )  ;
assign n28908 =  ( n36 ) & ( n28519 )  ;
assign n28909 =  ( n36 ) & ( n28521 )  ;
assign n28910 =  ( n36 ) & ( n28523 )  ;
assign n28911 =  ( n36 ) & ( n28525 )  ;
assign n28912 =  ( n36 ) & ( n28527 )  ;
assign n28913 =  ( n37 ) & ( n28497 )  ;
assign n28914 =  ( n37 ) & ( n28499 )  ;
assign n28915 =  ( n37 ) & ( n28501 )  ;
assign n28916 =  ( n37 ) & ( n28503 )  ;
assign n28917 =  ( n37 ) & ( n28505 )  ;
assign n28918 =  ( n37 ) & ( n28507 )  ;
assign n28919 =  ( n37 ) & ( n28509 )  ;
assign n28920 =  ( n37 ) & ( n28511 )  ;
assign n28921 =  ( n37 ) & ( n28513 )  ;
assign n28922 =  ( n37 ) & ( n28515 )  ;
assign n28923 =  ( n37 ) & ( n28517 )  ;
assign n28924 =  ( n37 ) & ( n28519 )  ;
assign n28925 =  ( n37 ) & ( n28521 )  ;
assign n28926 =  ( n37 ) & ( n28523 )  ;
assign n28927 =  ( n37 ) & ( n28525 )  ;
assign n28928 =  ( n37 ) & ( n28527 )  ;
assign n28929 =  ( n38 ) & ( n28497 )  ;
assign n28930 =  ( n38 ) & ( n28499 )  ;
assign n28931 =  ( n38 ) & ( n28501 )  ;
assign n28932 =  ( n38 ) & ( n28503 )  ;
assign n28933 =  ( n38 ) & ( n28505 )  ;
assign n28934 =  ( n38 ) & ( n28507 )  ;
assign n28935 =  ( n38 ) & ( n28509 )  ;
assign n28936 =  ( n38 ) & ( n28511 )  ;
assign n28937 =  ( n38 ) & ( n28513 )  ;
assign n28938 =  ( n38 ) & ( n28515 )  ;
assign n28939 =  ( n38 ) & ( n28517 )  ;
assign n28940 =  ( n38 ) & ( n28519 )  ;
assign n28941 =  ( n38 ) & ( n28521 )  ;
assign n28942 =  ( n38 ) & ( n28523 )  ;
assign n28943 =  ( n38 ) & ( n28525 )  ;
assign n28944 =  ( n38 ) & ( n28527 )  ;
assign n28945 =  ( n39 ) & ( n28497 )  ;
assign n28946 =  ( n39 ) & ( n28499 )  ;
assign n28947 =  ( n39 ) & ( n28501 )  ;
assign n28948 =  ( n39 ) & ( n28503 )  ;
assign n28949 =  ( n39 ) & ( n28505 )  ;
assign n28950 =  ( n39 ) & ( n28507 )  ;
assign n28951 =  ( n39 ) & ( n28509 )  ;
assign n28952 =  ( n39 ) & ( n28511 )  ;
assign n28953 =  ( n39 ) & ( n28513 )  ;
assign n28954 =  ( n39 ) & ( n28515 )  ;
assign n28955 =  ( n39 ) & ( n28517 )  ;
assign n28956 =  ( n39 ) & ( n28519 )  ;
assign n28957 =  ( n39 ) & ( n28521 )  ;
assign n28958 =  ( n39 ) & ( n28523 )  ;
assign n28959 =  ( n39 ) & ( n28525 )  ;
assign n28960 =  ( n39 ) & ( n28527 )  ;
assign n28961 =  ( n40 ) & ( n28497 )  ;
assign n28962 =  ( n40 ) & ( n28499 )  ;
assign n28963 =  ( n40 ) & ( n28501 )  ;
assign n28964 =  ( n40 ) & ( n28503 )  ;
assign n28965 =  ( n40 ) & ( n28505 )  ;
assign n28966 =  ( n40 ) & ( n28507 )  ;
assign n28967 =  ( n40 ) & ( n28509 )  ;
assign n28968 =  ( n40 ) & ( n28511 )  ;
assign n28969 =  ( n40 ) & ( n28513 )  ;
assign n28970 =  ( n40 ) & ( n28515 )  ;
assign n28971 =  ( n40 ) & ( n28517 )  ;
assign n28972 =  ( n40 ) & ( n28519 )  ;
assign n28973 =  ( n40 ) & ( n28521 )  ;
assign n28974 =  ( n40 ) & ( n28523 )  ;
assign n28975 =  ( n40 ) & ( n28525 )  ;
assign n28976 =  ( n40 ) & ( n28527 )  ;
assign n28977 =  ( n41 ) & ( n28497 )  ;
assign n28978 =  ( n41 ) & ( n28499 )  ;
assign n28979 =  ( n41 ) & ( n28501 )  ;
assign n28980 =  ( n41 ) & ( n28503 )  ;
assign n28981 =  ( n41 ) & ( n28505 )  ;
assign n28982 =  ( n41 ) & ( n28507 )  ;
assign n28983 =  ( n41 ) & ( n28509 )  ;
assign n28984 =  ( n41 ) & ( n28511 )  ;
assign n28985 =  ( n41 ) & ( n28513 )  ;
assign n28986 =  ( n41 ) & ( n28515 )  ;
assign n28987 =  ( n41 ) & ( n28517 )  ;
assign n28988 =  ( n41 ) & ( n28519 )  ;
assign n28989 =  ( n41 ) & ( n28521 )  ;
assign n28990 =  ( n41 ) & ( n28523 )  ;
assign n28991 =  ( n41 ) & ( n28525 )  ;
assign n28992 =  ( n41 ) & ( n28527 )  ;
assign n28993 =  ( n42 ) & ( n28497 )  ;
assign n28994 =  ( n42 ) & ( n28499 )  ;
assign n28995 =  ( n42 ) & ( n28501 )  ;
assign n28996 =  ( n42 ) & ( n28503 )  ;
assign n28997 =  ( n42 ) & ( n28505 )  ;
assign n28998 =  ( n42 ) & ( n28507 )  ;
assign n28999 =  ( n42 ) & ( n28509 )  ;
assign n29000 =  ( n42 ) & ( n28511 )  ;
assign n29001 =  ( n42 ) & ( n28513 )  ;
assign n29002 =  ( n42 ) & ( n28515 )  ;
assign n29003 =  ( n42 ) & ( n28517 )  ;
assign n29004 =  ( n42 ) & ( n28519 )  ;
assign n29005 =  ( n42 ) & ( n28521 )  ;
assign n29006 =  ( n42 ) & ( n28523 )  ;
assign n29007 =  ( n42 ) & ( n28525 )  ;
assign n29008 =  ( n42 ) & ( n28527 )  ;
assign n29009 =  ( n43 ) & ( n28497 )  ;
assign n29010 =  ( n43 ) & ( n28499 )  ;
assign n29011 =  ( n43 ) & ( n28501 )  ;
assign n29012 =  ( n43 ) & ( n28503 )  ;
assign n29013 =  ( n43 ) & ( n28505 )  ;
assign n29014 =  ( n43 ) & ( n28507 )  ;
assign n29015 =  ( n43 ) & ( n28509 )  ;
assign n29016 =  ( n43 ) & ( n28511 )  ;
assign n29017 =  ( n43 ) & ( n28513 )  ;
assign n29018 =  ( n43 ) & ( n28515 )  ;
assign n29019 =  ( n43 ) & ( n28517 )  ;
assign n29020 =  ( n43 ) & ( n28519 )  ;
assign n29021 =  ( n43 ) & ( n28521 )  ;
assign n29022 =  ( n43 ) & ( n28523 )  ;
assign n29023 =  ( n43 ) & ( n28525 )  ;
assign n29024 =  ( n43 ) & ( n28527 )  ;
assign n29025 =  ( n29024 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n29026 =  ( n29023 ) ? ( VREG_0_1 ) : ( n29025 ) ;
assign n29027 =  ( n29022 ) ? ( VREG_0_2 ) : ( n29026 ) ;
assign n29028 =  ( n29021 ) ? ( VREG_0_3 ) : ( n29027 ) ;
assign n29029 =  ( n29020 ) ? ( VREG_0_4 ) : ( n29028 ) ;
assign n29030 =  ( n29019 ) ? ( VREG_0_5 ) : ( n29029 ) ;
assign n29031 =  ( n29018 ) ? ( VREG_0_6 ) : ( n29030 ) ;
assign n29032 =  ( n29017 ) ? ( VREG_0_7 ) : ( n29031 ) ;
assign n29033 =  ( n29016 ) ? ( VREG_0_8 ) : ( n29032 ) ;
assign n29034 =  ( n29015 ) ? ( VREG_0_9 ) : ( n29033 ) ;
assign n29035 =  ( n29014 ) ? ( VREG_0_10 ) : ( n29034 ) ;
assign n29036 =  ( n29013 ) ? ( VREG_0_11 ) : ( n29035 ) ;
assign n29037 =  ( n29012 ) ? ( VREG_0_12 ) : ( n29036 ) ;
assign n29038 =  ( n29011 ) ? ( VREG_0_13 ) : ( n29037 ) ;
assign n29039 =  ( n29010 ) ? ( VREG_0_14 ) : ( n29038 ) ;
assign n29040 =  ( n29009 ) ? ( VREG_0_15 ) : ( n29039 ) ;
assign n29041 =  ( n29008 ) ? ( VREG_1_0 ) : ( n29040 ) ;
assign n29042 =  ( n29007 ) ? ( VREG_1_1 ) : ( n29041 ) ;
assign n29043 =  ( n29006 ) ? ( VREG_1_2 ) : ( n29042 ) ;
assign n29044 =  ( n29005 ) ? ( VREG_1_3 ) : ( n29043 ) ;
assign n29045 =  ( n29004 ) ? ( VREG_1_4 ) : ( n29044 ) ;
assign n29046 =  ( n29003 ) ? ( VREG_1_5 ) : ( n29045 ) ;
assign n29047 =  ( n29002 ) ? ( VREG_1_6 ) : ( n29046 ) ;
assign n29048 =  ( n29001 ) ? ( VREG_1_7 ) : ( n29047 ) ;
assign n29049 =  ( n29000 ) ? ( VREG_1_8 ) : ( n29048 ) ;
assign n29050 =  ( n28999 ) ? ( VREG_1_9 ) : ( n29049 ) ;
assign n29051 =  ( n28998 ) ? ( VREG_1_10 ) : ( n29050 ) ;
assign n29052 =  ( n28997 ) ? ( VREG_1_11 ) : ( n29051 ) ;
assign n29053 =  ( n28996 ) ? ( VREG_1_12 ) : ( n29052 ) ;
assign n29054 =  ( n28995 ) ? ( VREG_1_13 ) : ( n29053 ) ;
assign n29055 =  ( n28994 ) ? ( VREG_1_14 ) : ( n29054 ) ;
assign n29056 =  ( n28993 ) ? ( VREG_1_15 ) : ( n29055 ) ;
assign n29057 =  ( n28992 ) ? ( VREG_2_0 ) : ( n29056 ) ;
assign n29058 =  ( n28991 ) ? ( VREG_2_1 ) : ( n29057 ) ;
assign n29059 =  ( n28990 ) ? ( VREG_2_2 ) : ( n29058 ) ;
assign n29060 =  ( n28989 ) ? ( VREG_2_3 ) : ( n29059 ) ;
assign n29061 =  ( n28988 ) ? ( VREG_2_4 ) : ( n29060 ) ;
assign n29062 =  ( n28987 ) ? ( VREG_2_5 ) : ( n29061 ) ;
assign n29063 =  ( n28986 ) ? ( VREG_2_6 ) : ( n29062 ) ;
assign n29064 =  ( n28985 ) ? ( VREG_2_7 ) : ( n29063 ) ;
assign n29065 =  ( n28984 ) ? ( VREG_2_8 ) : ( n29064 ) ;
assign n29066 =  ( n28983 ) ? ( VREG_2_9 ) : ( n29065 ) ;
assign n29067 =  ( n28982 ) ? ( VREG_2_10 ) : ( n29066 ) ;
assign n29068 =  ( n28981 ) ? ( VREG_2_11 ) : ( n29067 ) ;
assign n29069 =  ( n28980 ) ? ( VREG_2_12 ) : ( n29068 ) ;
assign n29070 =  ( n28979 ) ? ( VREG_2_13 ) : ( n29069 ) ;
assign n29071 =  ( n28978 ) ? ( VREG_2_14 ) : ( n29070 ) ;
assign n29072 =  ( n28977 ) ? ( VREG_2_15 ) : ( n29071 ) ;
assign n29073 =  ( n28976 ) ? ( VREG_3_0 ) : ( n29072 ) ;
assign n29074 =  ( n28975 ) ? ( VREG_3_1 ) : ( n29073 ) ;
assign n29075 =  ( n28974 ) ? ( VREG_3_2 ) : ( n29074 ) ;
assign n29076 =  ( n28973 ) ? ( VREG_3_3 ) : ( n29075 ) ;
assign n29077 =  ( n28972 ) ? ( VREG_3_4 ) : ( n29076 ) ;
assign n29078 =  ( n28971 ) ? ( VREG_3_5 ) : ( n29077 ) ;
assign n29079 =  ( n28970 ) ? ( VREG_3_6 ) : ( n29078 ) ;
assign n29080 =  ( n28969 ) ? ( VREG_3_7 ) : ( n29079 ) ;
assign n29081 =  ( n28968 ) ? ( VREG_3_8 ) : ( n29080 ) ;
assign n29082 =  ( n28967 ) ? ( VREG_3_9 ) : ( n29081 ) ;
assign n29083 =  ( n28966 ) ? ( VREG_3_10 ) : ( n29082 ) ;
assign n29084 =  ( n28965 ) ? ( VREG_3_11 ) : ( n29083 ) ;
assign n29085 =  ( n28964 ) ? ( VREG_3_12 ) : ( n29084 ) ;
assign n29086 =  ( n28963 ) ? ( VREG_3_13 ) : ( n29085 ) ;
assign n29087 =  ( n28962 ) ? ( VREG_3_14 ) : ( n29086 ) ;
assign n29088 =  ( n28961 ) ? ( VREG_3_15 ) : ( n29087 ) ;
assign n29089 =  ( n28960 ) ? ( VREG_4_0 ) : ( n29088 ) ;
assign n29090 =  ( n28959 ) ? ( VREG_4_1 ) : ( n29089 ) ;
assign n29091 =  ( n28958 ) ? ( VREG_4_2 ) : ( n29090 ) ;
assign n29092 =  ( n28957 ) ? ( VREG_4_3 ) : ( n29091 ) ;
assign n29093 =  ( n28956 ) ? ( VREG_4_4 ) : ( n29092 ) ;
assign n29094 =  ( n28955 ) ? ( VREG_4_5 ) : ( n29093 ) ;
assign n29095 =  ( n28954 ) ? ( VREG_4_6 ) : ( n29094 ) ;
assign n29096 =  ( n28953 ) ? ( VREG_4_7 ) : ( n29095 ) ;
assign n29097 =  ( n28952 ) ? ( VREG_4_8 ) : ( n29096 ) ;
assign n29098 =  ( n28951 ) ? ( VREG_4_9 ) : ( n29097 ) ;
assign n29099 =  ( n28950 ) ? ( VREG_4_10 ) : ( n29098 ) ;
assign n29100 =  ( n28949 ) ? ( VREG_4_11 ) : ( n29099 ) ;
assign n29101 =  ( n28948 ) ? ( VREG_4_12 ) : ( n29100 ) ;
assign n29102 =  ( n28947 ) ? ( VREG_4_13 ) : ( n29101 ) ;
assign n29103 =  ( n28946 ) ? ( VREG_4_14 ) : ( n29102 ) ;
assign n29104 =  ( n28945 ) ? ( VREG_4_15 ) : ( n29103 ) ;
assign n29105 =  ( n28944 ) ? ( VREG_5_0 ) : ( n29104 ) ;
assign n29106 =  ( n28943 ) ? ( VREG_5_1 ) : ( n29105 ) ;
assign n29107 =  ( n28942 ) ? ( VREG_5_2 ) : ( n29106 ) ;
assign n29108 =  ( n28941 ) ? ( VREG_5_3 ) : ( n29107 ) ;
assign n29109 =  ( n28940 ) ? ( VREG_5_4 ) : ( n29108 ) ;
assign n29110 =  ( n28939 ) ? ( VREG_5_5 ) : ( n29109 ) ;
assign n29111 =  ( n28938 ) ? ( VREG_5_6 ) : ( n29110 ) ;
assign n29112 =  ( n28937 ) ? ( VREG_5_7 ) : ( n29111 ) ;
assign n29113 =  ( n28936 ) ? ( VREG_5_8 ) : ( n29112 ) ;
assign n29114 =  ( n28935 ) ? ( VREG_5_9 ) : ( n29113 ) ;
assign n29115 =  ( n28934 ) ? ( VREG_5_10 ) : ( n29114 ) ;
assign n29116 =  ( n28933 ) ? ( VREG_5_11 ) : ( n29115 ) ;
assign n29117 =  ( n28932 ) ? ( VREG_5_12 ) : ( n29116 ) ;
assign n29118 =  ( n28931 ) ? ( VREG_5_13 ) : ( n29117 ) ;
assign n29119 =  ( n28930 ) ? ( VREG_5_14 ) : ( n29118 ) ;
assign n29120 =  ( n28929 ) ? ( VREG_5_15 ) : ( n29119 ) ;
assign n29121 =  ( n28928 ) ? ( VREG_6_0 ) : ( n29120 ) ;
assign n29122 =  ( n28927 ) ? ( VREG_6_1 ) : ( n29121 ) ;
assign n29123 =  ( n28926 ) ? ( VREG_6_2 ) : ( n29122 ) ;
assign n29124 =  ( n28925 ) ? ( VREG_6_3 ) : ( n29123 ) ;
assign n29125 =  ( n28924 ) ? ( VREG_6_4 ) : ( n29124 ) ;
assign n29126 =  ( n28923 ) ? ( VREG_6_5 ) : ( n29125 ) ;
assign n29127 =  ( n28922 ) ? ( VREG_6_6 ) : ( n29126 ) ;
assign n29128 =  ( n28921 ) ? ( VREG_6_7 ) : ( n29127 ) ;
assign n29129 =  ( n28920 ) ? ( VREG_6_8 ) : ( n29128 ) ;
assign n29130 =  ( n28919 ) ? ( VREG_6_9 ) : ( n29129 ) ;
assign n29131 =  ( n28918 ) ? ( VREG_6_10 ) : ( n29130 ) ;
assign n29132 =  ( n28917 ) ? ( VREG_6_11 ) : ( n29131 ) ;
assign n29133 =  ( n28916 ) ? ( VREG_6_12 ) : ( n29132 ) ;
assign n29134 =  ( n28915 ) ? ( VREG_6_13 ) : ( n29133 ) ;
assign n29135 =  ( n28914 ) ? ( VREG_6_14 ) : ( n29134 ) ;
assign n29136 =  ( n28913 ) ? ( VREG_6_15 ) : ( n29135 ) ;
assign n29137 =  ( n28912 ) ? ( VREG_7_0 ) : ( n29136 ) ;
assign n29138 =  ( n28911 ) ? ( VREG_7_1 ) : ( n29137 ) ;
assign n29139 =  ( n28910 ) ? ( VREG_7_2 ) : ( n29138 ) ;
assign n29140 =  ( n28909 ) ? ( VREG_7_3 ) : ( n29139 ) ;
assign n29141 =  ( n28908 ) ? ( VREG_7_4 ) : ( n29140 ) ;
assign n29142 =  ( n28907 ) ? ( VREG_7_5 ) : ( n29141 ) ;
assign n29143 =  ( n28906 ) ? ( VREG_7_6 ) : ( n29142 ) ;
assign n29144 =  ( n28905 ) ? ( VREG_7_7 ) : ( n29143 ) ;
assign n29145 =  ( n28904 ) ? ( VREG_7_8 ) : ( n29144 ) ;
assign n29146 =  ( n28903 ) ? ( VREG_7_9 ) : ( n29145 ) ;
assign n29147 =  ( n28902 ) ? ( VREG_7_10 ) : ( n29146 ) ;
assign n29148 =  ( n28901 ) ? ( VREG_7_11 ) : ( n29147 ) ;
assign n29149 =  ( n28900 ) ? ( VREG_7_12 ) : ( n29148 ) ;
assign n29150 =  ( n28899 ) ? ( VREG_7_13 ) : ( n29149 ) ;
assign n29151 =  ( n28898 ) ? ( VREG_7_14 ) : ( n29150 ) ;
assign n29152 =  ( n28897 ) ? ( VREG_7_15 ) : ( n29151 ) ;
assign n29153 =  ( n28896 ) ? ( VREG_8_0 ) : ( n29152 ) ;
assign n29154 =  ( n28895 ) ? ( VREG_8_1 ) : ( n29153 ) ;
assign n29155 =  ( n28894 ) ? ( VREG_8_2 ) : ( n29154 ) ;
assign n29156 =  ( n28893 ) ? ( VREG_8_3 ) : ( n29155 ) ;
assign n29157 =  ( n28892 ) ? ( VREG_8_4 ) : ( n29156 ) ;
assign n29158 =  ( n28891 ) ? ( VREG_8_5 ) : ( n29157 ) ;
assign n29159 =  ( n28890 ) ? ( VREG_8_6 ) : ( n29158 ) ;
assign n29160 =  ( n28889 ) ? ( VREG_8_7 ) : ( n29159 ) ;
assign n29161 =  ( n28888 ) ? ( VREG_8_8 ) : ( n29160 ) ;
assign n29162 =  ( n28887 ) ? ( VREG_8_9 ) : ( n29161 ) ;
assign n29163 =  ( n28886 ) ? ( VREG_8_10 ) : ( n29162 ) ;
assign n29164 =  ( n28885 ) ? ( VREG_8_11 ) : ( n29163 ) ;
assign n29165 =  ( n28884 ) ? ( VREG_8_12 ) : ( n29164 ) ;
assign n29166 =  ( n28883 ) ? ( VREG_8_13 ) : ( n29165 ) ;
assign n29167 =  ( n28882 ) ? ( VREG_8_14 ) : ( n29166 ) ;
assign n29168 =  ( n28881 ) ? ( VREG_8_15 ) : ( n29167 ) ;
assign n29169 =  ( n28880 ) ? ( VREG_9_0 ) : ( n29168 ) ;
assign n29170 =  ( n28879 ) ? ( VREG_9_1 ) : ( n29169 ) ;
assign n29171 =  ( n28878 ) ? ( VREG_9_2 ) : ( n29170 ) ;
assign n29172 =  ( n28877 ) ? ( VREG_9_3 ) : ( n29171 ) ;
assign n29173 =  ( n28876 ) ? ( VREG_9_4 ) : ( n29172 ) ;
assign n29174 =  ( n28875 ) ? ( VREG_9_5 ) : ( n29173 ) ;
assign n29175 =  ( n28874 ) ? ( VREG_9_6 ) : ( n29174 ) ;
assign n29176 =  ( n28873 ) ? ( VREG_9_7 ) : ( n29175 ) ;
assign n29177 =  ( n28872 ) ? ( VREG_9_8 ) : ( n29176 ) ;
assign n29178 =  ( n28871 ) ? ( VREG_9_9 ) : ( n29177 ) ;
assign n29179 =  ( n28870 ) ? ( VREG_9_10 ) : ( n29178 ) ;
assign n29180 =  ( n28869 ) ? ( VREG_9_11 ) : ( n29179 ) ;
assign n29181 =  ( n28868 ) ? ( VREG_9_12 ) : ( n29180 ) ;
assign n29182 =  ( n28867 ) ? ( VREG_9_13 ) : ( n29181 ) ;
assign n29183 =  ( n28866 ) ? ( VREG_9_14 ) : ( n29182 ) ;
assign n29184 =  ( n28865 ) ? ( VREG_9_15 ) : ( n29183 ) ;
assign n29185 =  ( n28864 ) ? ( VREG_10_0 ) : ( n29184 ) ;
assign n29186 =  ( n28863 ) ? ( VREG_10_1 ) : ( n29185 ) ;
assign n29187 =  ( n28862 ) ? ( VREG_10_2 ) : ( n29186 ) ;
assign n29188 =  ( n28861 ) ? ( VREG_10_3 ) : ( n29187 ) ;
assign n29189 =  ( n28860 ) ? ( VREG_10_4 ) : ( n29188 ) ;
assign n29190 =  ( n28859 ) ? ( VREG_10_5 ) : ( n29189 ) ;
assign n29191 =  ( n28858 ) ? ( VREG_10_6 ) : ( n29190 ) ;
assign n29192 =  ( n28857 ) ? ( VREG_10_7 ) : ( n29191 ) ;
assign n29193 =  ( n28856 ) ? ( VREG_10_8 ) : ( n29192 ) ;
assign n29194 =  ( n28855 ) ? ( VREG_10_9 ) : ( n29193 ) ;
assign n29195 =  ( n28854 ) ? ( VREG_10_10 ) : ( n29194 ) ;
assign n29196 =  ( n28853 ) ? ( VREG_10_11 ) : ( n29195 ) ;
assign n29197 =  ( n28852 ) ? ( VREG_10_12 ) : ( n29196 ) ;
assign n29198 =  ( n28851 ) ? ( VREG_10_13 ) : ( n29197 ) ;
assign n29199 =  ( n28850 ) ? ( VREG_10_14 ) : ( n29198 ) ;
assign n29200 =  ( n28849 ) ? ( VREG_10_15 ) : ( n29199 ) ;
assign n29201 =  ( n28848 ) ? ( VREG_11_0 ) : ( n29200 ) ;
assign n29202 =  ( n28847 ) ? ( VREG_11_1 ) : ( n29201 ) ;
assign n29203 =  ( n28846 ) ? ( VREG_11_2 ) : ( n29202 ) ;
assign n29204 =  ( n28845 ) ? ( VREG_11_3 ) : ( n29203 ) ;
assign n29205 =  ( n28844 ) ? ( VREG_11_4 ) : ( n29204 ) ;
assign n29206 =  ( n28843 ) ? ( VREG_11_5 ) : ( n29205 ) ;
assign n29207 =  ( n28842 ) ? ( VREG_11_6 ) : ( n29206 ) ;
assign n29208 =  ( n28841 ) ? ( VREG_11_7 ) : ( n29207 ) ;
assign n29209 =  ( n28840 ) ? ( VREG_11_8 ) : ( n29208 ) ;
assign n29210 =  ( n28839 ) ? ( VREG_11_9 ) : ( n29209 ) ;
assign n29211 =  ( n28838 ) ? ( VREG_11_10 ) : ( n29210 ) ;
assign n29212 =  ( n28837 ) ? ( VREG_11_11 ) : ( n29211 ) ;
assign n29213 =  ( n28836 ) ? ( VREG_11_12 ) : ( n29212 ) ;
assign n29214 =  ( n28835 ) ? ( VREG_11_13 ) : ( n29213 ) ;
assign n29215 =  ( n28834 ) ? ( VREG_11_14 ) : ( n29214 ) ;
assign n29216 =  ( n28833 ) ? ( VREG_11_15 ) : ( n29215 ) ;
assign n29217 =  ( n28832 ) ? ( VREG_12_0 ) : ( n29216 ) ;
assign n29218 =  ( n28831 ) ? ( VREG_12_1 ) : ( n29217 ) ;
assign n29219 =  ( n28830 ) ? ( VREG_12_2 ) : ( n29218 ) ;
assign n29220 =  ( n28829 ) ? ( VREG_12_3 ) : ( n29219 ) ;
assign n29221 =  ( n28828 ) ? ( VREG_12_4 ) : ( n29220 ) ;
assign n29222 =  ( n28827 ) ? ( VREG_12_5 ) : ( n29221 ) ;
assign n29223 =  ( n28826 ) ? ( VREG_12_6 ) : ( n29222 ) ;
assign n29224 =  ( n28825 ) ? ( VREG_12_7 ) : ( n29223 ) ;
assign n29225 =  ( n28824 ) ? ( VREG_12_8 ) : ( n29224 ) ;
assign n29226 =  ( n28823 ) ? ( VREG_12_9 ) : ( n29225 ) ;
assign n29227 =  ( n28822 ) ? ( VREG_12_10 ) : ( n29226 ) ;
assign n29228 =  ( n28821 ) ? ( VREG_12_11 ) : ( n29227 ) ;
assign n29229 =  ( n28820 ) ? ( VREG_12_12 ) : ( n29228 ) ;
assign n29230 =  ( n28819 ) ? ( VREG_12_13 ) : ( n29229 ) ;
assign n29231 =  ( n28818 ) ? ( VREG_12_14 ) : ( n29230 ) ;
assign n29232 =  ( n28817 ) ? ( VREG_12_15 ) : ( n29231 ) ;
assign n29233 =  ( n28816 ) ? ( VREG_13_0 ) : ( n29232 ) ;
assign n29234 =  ( n28815 ) ? ( VREG_13_1 ) : ( n29233 ) ;
assign n29235 =  ( n28814 ) ? ( VREG_13_2 ) : ( n29234 ) ;
assign n29236 =  ( n28813 ) ? ( VREG_13_3 ) : ( n29235 ) ;
assign n29237 =  ( n28812 ) ? ( VREG_13_4 ) : ( n29236 ) ;
assign n29238 =  ( n28811 ) ? ( VREG_13_5 ) : ( n29237 ) ;
assign n29239 =  ( n28810 ) ? ( VREG_13_6 ) : ( n29238 ) ;
assign n29240 =  ( n28809 ) ? ( VREG_13_7 ) : ( n29239 ) ;
assign n29241 =  ( n28808 ) ? ( VREG_13_8 ) : ( n29240 ) ;
assign n29242 =  ( n28807 ) ? ( VREG_13_9 ) : ( n29241 ) ;
assign n29243 =  ( n28806 ) ? ( VREG_13_10 ) : ( n29242 ) ;
assign n29244 =  ( n28805 ) ? ( VREG_13_11 ) : ( n29243 ) ;
assign n29245 =  ( n28804 ) ? ( VREG_13_12 ) : ( n29244 ) ;
assign n29246 =  ( n28803 ) ? ( VREG_13_13 ) : ( n29245 ) ;
assign n29247 =  ( n28802 ) ? ( VREG_13_14 ) : ( n29246 ) ;
assign n29248 =  ( n28801 ) ? ( VREG_13_15 ) : ( n29247 ) ;
assign n29249 =  ( n28800 ) ? ( VREG_14_0 ) : ( n29248 ) ;
assign n29250 =  ( n28799 ) ? ( VREG_14_1 ) : ( n29249 ) ;
assign n29251 =  ( n28798 ) ? ( VREG_14_2 ) : ( n29250 ) ;
assign n29252 =  ( n28797 ) ? ( VREG_14_3 ) : ( n29251 ) ;
assign n29253 =  ( n28796 ) ? ( VREG_14_4 ) : ( n29252 ) ;
assign n29254 =  ( n28795 ) ? ( VREG_14_5 ) : ( n29253 ) ;
assign n29255 =  ( n28794 ) ? ( VREG_14_6 ) : ( n29254 ) ;
assign n29256 =  ( n28793 ) ? ( VREG_14_7 ) : ( n29255 ) ;
assign n29257 =  ( n28792 ) ? ( VREG_14_8 ) : ( n29256 ) ;
assign n29258 =  ( n28791 ) ? ( VREG_14_9 ) : ( n29257 ) ;
assign n29259 =  ( n28790 ) ? ( VREG_14_10 ) : ( n29258 ) ;
assign n29260 =  ( n28789 ) ? ( VREG_14_11 ) : ( n29259 ) ;
assign n29261 =  ( n28788 ) ? ( VREG_14_12 ) : ( n29260 ) ;
assign n29262 =  ( n28787 ) ? ( VREG_14_13 ) : ( n29261 ) ;
assign n29263 =  ( n28786 ) ? ( VREG_14_14 ) : ( n29262 ) ;
assign n29264 =  ( n28785 ) ? ( VREG_14_15 ) : ( n29263 ) ;
assign n29265 =  ( n28784 ) ? ( VREG_15_0 ) : ( n29264 ) ;
assign n29266 =  ( n28783 ) ? ( VREG_15_1 ) : ( n29265 ) ;
assign n29267 =  ( n28782 ) ? ( VREG_15_2 ) : ( n29266 ) ;
assign n29268 =  ( n28781 ) ? ( VREG_15_3 ) : ( n29267 ) ;
assign n29269 =  ( n28780 ) ? ( VREG_15_4 ) : ( n29268 ) ;
assign n29270 =  ( n28779 ) ? ( VREG_15_5 ) : ( n29269 ) ;
assign n29271 =  ( n28778 ) ? ( VREG_15_6 ) : ( n29270 ) ;
assign n29272 =  ( n28777 ) ? ( VREG_15_7 ) : ( n29271 ) ;
assign n29273 =  ( n28776 ) ? ( VREG_15_8 ) : ( n29272 ) ;
assign n29274 =  ( n28775 ) ? ( VREG_15_9 ) : ( n29273 ) ;
assign n29275 =  ( n28774 ) ? ( VREG_15_10 ) : ( n29274 ) ;
assign n29276 =  ( n28773 ) ? ( VREG_15_11 ) : ( n29275 ) ;
assign n29277 =  ( n28772 ) ? ( VREG_15_12 ) : ( n29276 ) ;
assign n29278 =  ( n28771 ) ? ( VREG_15_13 ) : ( n29277 ) ;
assign n29279 =  ( n28770 ) ? ( VREG_15_14 ) : ( n29278 ) ;
assign n29280 =  ( n28769 ) ? ( VREG_15_15 ) : ( n29279 ) ;
assign n29281 =  ( n28768 ) ? ( VREG_16_0 ) : ( n29280 ) ;
assign n29282 =  ( n28767 ) ? ( VREG_16_1 ) : ( n29281 ) ;
assign n29283 =  ( n28766 ) ? ( VREG_16_2 ) : ( n29282 ) ;
assign n29284 =  ( n28765 ) ? ( VREG_16_3 ) : ( n29283 ) ;
assign n29285 =  ( n28764 ) ? ( VREG_16_4 ) : ( n29284 ) ;
assign n29286 =  ( n28763 ) ? ( VREG_16_5 ) : ( n29285 ) ;
assign n29287 =  ( n28762 ) ? ( VREG_16_6 ) : ( n29286 ) ;
assign n29288 =  ( n28761 ) ? ( VREG_16_7 ) : ( n29287 ) ;
assign n29289 =  ( n28760 ) ? ( VREG_16_8 ) : ( n29288 ) ;
assign n29290 =  ( n28759 ) ? ( VREG_16_9 ) : ( n29289 ) ;
assign n29291 =  ( n28758 ) ? ( VREG_16_10 ) : ( n29290 ) ;
assign n29292 =  ( n28757 ) ? ( VREG_16_11 ) : ( n29291 ) ;
assign n29293 =  ( n28756 ) ? ( VREG_16_12 ) : ( n29292 ) ;
assign n29294 =  ( n28755 ) ? ( VREG_16_13 ) : ( n29293 ) ;
assign n29295 =  ( n28754 ) ? ( VREG_16_14 ) : ( n29294 ) ;
assign n29296 =  ( n28753 ) ? ( VREG_16_15 ) : ( n29295 ) ;
assign n29297 =  ( n28752 ) ? ( VREG_17_0 ) : ( n29296 ) ;
assign n29298 =  ( n28751 ) ? ( VREG_17_1 ) : ( n29297 ) ;
assign n29299 =  ( n28750 ) ? ( VREG_17_2 ) : ( n29298 ) ;
assign n29300 =  ( n28749 ) ? ( VREG_17_3 ) : ( n29299 ) ;
assign n29301 =  ( n28748 ) ? ( VREG_17_4 ) : ( n29300 ) ;
assign n29302 =  ( n28747 ) ? ( VREG_17_5 ) : ( n29301 ) ;
assign n29303 =  ( n28746 ) ? ( VREG_17_6 ) : ( n29302 ) ;
assign n29304 =  ( n28745 ) ? ( VREG_17_7 ) : ( n29303 ) ;
assign n29305 =  ( n28744 ) ? ( VREG_17_8 ) : ( n29304 ) ;
assign n29306 =  ( n28743 ) ? ( VREG_17_9 ) : ( n29305 ) ;
assign n29307 =  ( n28742 ) ? ( VREG_17_10 ) : ( n29306 ) ;
assign n29308 =  ( n28741 ) ? ( VREG_17_11 ) : ( n29307 ) ;
assign n29309 =  ( n28740 ) ? ( VREG_17_12 ) : ( n29308 ) ;
assign n29310 =  ( n28739 ) ? ( VREG_17_13 ) : ( n29309 ) ;
assign n29311 =  ( n28738 ) ? ( VREG_17_14 ) : ( n29310 ) ;
assign n29312 =  ( n28737 ) ? ( VREG_17_15 ) : ( n29311 ) ;
assign n29313 =  ( n28736 ) ? ( VREG_18_0 ) : ( n29312 ) ;
assign n29314 =  ( n28735 ) ? ( VREG_18_1 ) : ( n29313 ) ;
assign n29315 =  ( n28734 ) ? ( VREG_18_2 ) : ( n29314 ) ;
assign n29316 =  ( n28733 ) ? ( VREG_18_3 ) : ( n29315 ) ;
assign n29317 =  ( n28732 ) ? ( VREG_18_4 ) : ( n29316 ) ;
assign n29318 =  ( n28731 ) ? ( VREG_18_5 ) : ( n29317 ) ;
assign n29319 =  ( n28730 ) ? ( VREG_18_6 ) : ( n29318 ) ;
assign n29320 =  ( n28729 ) ? ( VREG_18_7 ) : ( n29319 ) ;
assign n29321 =  ( n28728 ) ? ( VREG_18_8 ) : ( n29320 ) ;
assign n29322 =  ( n28727 ) ? ( VREG_18_9 ) : ( n29321 ) ;
assign n29323 =  ( n28726 ) ? ( VREG_18_10 ) : ( n29322 ) ;
assign n29324 =  ( n28725 ) ? ( VREG_18_11 ) : ( n29323 ) ;
assign n29325 =  ( n28724 ) ? ( VREG_18_12 ) : ( n29324 ) ;
assign n29326 =  ( n28723 ) ? ( VREG_18_13 ) : ( n29325 ) ;
assign n29327 =  ( n28722 ) ? ( VREG_18_14 ) : ( n29326 ) ;
assign n29328 =  ( n28721 ) ? ( VREG_18_15 ) : ( n29327 ) ;
assign n29329 =  ( n28720 ) ? ( VREG_19_0 ) : ( n29328 ) ;
assign n29330 =  ( n28719 ) ? ( VREG_19_1 ) : ( n29329 ) ;
assign n29331 =  ( n28718 ) ? ( VREG_19_2 ) : ( n29330 ) ;
assign n29332 =  ( n28717 ) ? ( VREG_19_3 ) : ( n29331 ) ;
assign n29333 =  ( n28716 ) ? ( VREG_19_4 ) : ( n29332 ) ;
assign n29334 =  ( n28715 ) ? ( VREG_19_5 ) : ( n29333 ) ;
assign n29335 =  ( n28714 ) ? ( VREG_19_6 ) : ( n29334 ) ;
assign n29336 =  ( n28713 ) ? ( VREG_19_7 ) : ( n29335 ) ;
assign n29337 =  ( n28712 ) ? ( VREG_19_8 ) : ( n29336 ) ;
assign n29338 =  ( n28711 ) ? ( VREG_19_9 ) : ( n29337 ) ;
assign n29339 =  ( n28710 ) ? ( VREG_19_10 ) : ( n29338 ) ;
assign n29340 =  ( n28709 ) ? ( VREG_19_11 ) : ( n29339 ) ;
assign n29341 =  ( n28708 ) ? ( VREG_19_12 ) : ( n29340 ) ;
assign n29342 =  ( n28707 ) ? ( VREG_19_13 ) : ( n29341 ) ;
assign n29343 =  ( n28706 ) ? ( VREG_19_14 ) : ( n29342 ) ;
assign n29344 =  ( n28705 ) ? ( VREG_19_15 ) : ( n29343 ) ;
assign n29345 =  ( n28704 ) ? ( VREG_20_0 ) : ( n29344 ) ;
assign n29346 =  ( n28703 ) ? ( VREG_20_1 ) : ( n29345 ) ;
assign n29347 =  ( n28702 ) ? ( VREG_20_2 ) : ( n29346 ) ;
assign n29348 =  ( n28701 ) ? ( VREG_20_3 ) : ( n29347 ) ;
assign n29349 =  ( n28700 ) ? ( VREG_20_4 ) : ( n29348 ) ;
assign n29350 =  ( n28699 ) ? ( VREG_20_5 ) : ( n29349 ) ;
assign n29351 =  ( n28698 ) ? ( VREG_20_6 ) : ( n29350 ) ;
assign n29352 =  ( n28697 ) ? ( VREG_20_7 ) : ( n29351 ) ;
assign n29353 =  ( n28696 ) ? ( VREG_20_8 ) : ( n29352 ) ;
assign n29354 =  ( n28695 ) ? ( VREG_20_9 ) : ( n29353 ) ;
assign n29355 =  ( n28694 ) ? ( VREG_20_10 ) : ( n29354 ) ;
assign n29356 =  ( n28693 ) ? ( VREG_20_11 ) : ( n29355 ) ;
assign n29357 =  ( n28692 ) ? ( VREG_20_12 ) : ( n29356 ) ;
assign n29358 =  ( n28691 ) ? ( VREG_20_13 ) : ( n29357 ) ;
assign n29359 =  ( n28690 ) ? ( VREG_20_14 ) : ( n29358 ) ;
assign n29360 =  ( n28689 ) ? ( VREG_20_15 ) : ( n29359 ) ;
assign n29361 =  ( n28688 ) ? ( VREG_21_0 ) : ( n29360 ) ;
assign n29362 =  ( n28687 ) ? ( VREG_21_1 ) : ( n29361 ) ;
assign n29363 =  ( n28686 ) ? ( VREG_21_2 ) : ( n29362 ) ;
assign n29364 =  ( n28685 ) ? ( VREG_21_3 ) : ( n29363 ) ;
assign n29365 =  ( n28684 ) ? ( VREG_21_4 ) : ( n29364 ) ;
assign n29366 =  ( n28683 ) ? ( VREG_21_5 ) : ( n29365 ) ;
assign n29367 =  ( n28682 ) ? ( VREG_21_6 ) : ( n29366 ) ;
assign n29368 =  ( n28681 ) ? ( VREG_21_7 ) : ( n29367 ) ;
assign n29369 =  ( n28680 ) ? ( VREG_21_8 ) : ( n29368 ) ;
assign n29370 =  ( n28679 ) ? ( VREG_21_9 ) : ( n29369 ) ;
assign n29371 =  ( n28678 ) ? ( VREG_21_10 ) : ( n29370 ) ;
assign n29372 =  ( n28677 ) ? ( VREG_21_11 ) : ( n29371 ) ;
assign n29373 =  ( n28676 ) ? ( VREG_21_12 ) : ( n29372 ) ;
assign n29374 =  ( n28675 ) ? ( VREG_21_13 ) : ( n29373 ) ;
assign n29375 =  ( n28674 ) ? ( VREG_21_14 ) : ( n29374 ) ;
assign n29376 =  ( n28673 ) ? ( VREG_21_15 ) : ( n29375 ) ;
assign n29377 =  ( n28672 ) ? ( VREG_22_0 ) : ( n29376 ) ;
assign n29378 =  ( n28671 ) ? ( VREG_22_1 ) : ( n29377 ) ;
assign n29379 =  ( n28670 ) ? ( VREG_22_2 ) : ( n29378 ) ;
assign n29380 =  ( n28669 ) ? ( VREG_22_3 ) : ( n29379 ) ;
assign n29381 =  ( n28668 ) ? ( VREG_22_4 ) : ( n29380 ) ;
assign n29382 =  ( n28667 ) ? ( VREG_22_5 ) : ( n29381 ) ;
assign n29383 =  ( n28666 ) ? ( VREG_22_6 ) : ( n29382 ) ;
assign n29384 =  ( n28665 ) ? ( VREG_22_7 ) : ( n29383 ) ;
assign n29385 =  ( n28664 ) ? ( VREG_22_8 ) : ( n29384 ) ;
assign n29386 =  ( n28663 ) ? ( VREG_22_9 ) : ( n29385 ) ;
assign n29387 =  ( n28662 ) ? ( VREG_22_10 ) : ( n29386 ) ;
assign n29388 =  ( n28661 ) ? ( VREG_22_11 ) : ( n29387 ) ;
assign n29389 =  ( n28660 ) ? ( VREG_22_12 ) : ( n29388 ) ;
assign n29390 =  ( n28659 ) ? ( VREG_22_13 ) : ( n29389 ) ;
assign n29391 =  ( n28658 ) ? ( VREG_22_14 ) : ( n29390 ) ;
assign n29392 =  ( n28657 ) ? ( VREG_22_15 ) : ( n29391 ) ;
assign n29393 =  ( n28656 ) ? ( VREG_23_0 ) : ( n29392 ) ;
assign n29394 =  ( n28655 ) ? ( VREG_23_1 ) : ( n29393 ) ;
assign n29395 =  ( n28654 ) ? ( VREG_23_2 ) : ( n29394 ) ;
assign n29396 =  ( n28653 ) ? ( VREG_23_3 ) : ( n29395 ) ;
assign n29397 =  ( n28652 ) ? ( VREG_23_4 ) : ( n29396 ) ;
assign n29398 =  ( n28651 ) ? ( VREG_23_5 ) : ( n29397 ) ;
assign n29399 =  ( n28650 ) ? ( VREG_23_6 ) : ( n29398 ) ;
assign n29400 =  ( n28649 ) ? ( VREG_23_7 ) : ( n29399 ) ;
assign n29401 =  ( n28648 ) ? ( VREG_23_8 ) : ( n29400 ) ;
assign n29402 =  ( n28647 ) ? ( VREG_23_9 ) : ( n29401 ) ;
assign n29403 =  ( n28646 ) ? ( VREG_23_10 ) : ( n29402 ) ;
assign n29404 =  ( n28645 ) ? ( VREG_23_11 ) : ( n29403 ) ;
assign n29405 =  ( n28644 ) ? ( VREG_23_12 ) : ( n29404 ) ;
assign n29406 =  ( n28643 ) ? ( VREG_23_13 ) : ( n29405 ) ;
assign n29407 =  ( n28642 ) ? ( VREG_23_14 ) : ( n29406 ) ;
assign n29408 =  ( n28641 ) ? ( VREG_23_15 ) : ( n29407 ) ;
assign n29409 =  ( n28640 ) ? ( VREG_24_0 ) : ( n29408 ) ;
assign n29410 =  ( n28639 ) ? ( VREG_24_1 ) : ( n29409 ) ;
assign n29411 =  ( n28638 ) ? ( VREG_24_2 ) : ( n29410 ) ;
assign n29412 =  ( n28637 ) ? ( VREG_24_3 ) : ( n29411 ) ;
assign n29413 =  ( n28636 ) ? ( VREG_24_4 ) : ( n29412 ) ;
assign n29414 =  ( n28635 ) ? ( VREG_24_5 ) : ( n29413 ) ;
assign n29415 =  ( n28634 ) ? ( VREG_24_6 ) : ( n29414 ) ;
assign n29416 =  ( n28633 ) ? ( VREG_24_7 ) : ( n29415 ) ;
assign n29417 =  ( n28632 ) ? ( VREG_24_8 ) : ( n29416 ) ;
assign n29418 =  ( n28631 ) ? ( VREG_24_9 ) : ( n29417 ) ;
assign n29419 =  ( n28630 ) ? ( VREG_24_10 ) : ( n29418 ) ;
assign n29420 =  ( n28629 ) ? ( VREG_24_11 ) : ( n29419 ) ;
assign n29421 =  ( n28628 ) ? ( VREG_24_12 ) : ( n29420 ) ;
assign n29422 =  ( n28627 ) ? ( VREG_24_13 ) : ( n29421 ) ;
assign n29423 =  ( n28626 ) ? ( VREG_24_14 ) : ( n29422 ) ;
assign n29424 =  ( n28625 ) ? ( VREG_24_15 ) : ( n29423 ) ;
assign n29425 =  ( n28624 ) ? ( VREG_25_0 ) : ( n29424 ) ;
assign n29426 =  ( n28623 ) ? ( VREG_25_1 ) : ( n29425 ) ;
assign n29427 =  ( n28622 ) ? ( VREG_25_2 ) : ( n29426 ) ;
assign n29428 =  ( n28621 ) ? ( VREG_25_3 ) : ( n29427 ) ;
assign n29429 =  ( n28620 ) ? ( VREG_25_4 ) : ( n29428 ) ;
assign n29430 =  ( n28619 ) ? ( VREG_25_5 ) : ( n29429 ) ;
assign n29431 =  ( n28618 ) ? ( VREG_25_6 ) : ( n29430 ) ;
assign n29432 =  ( n28617 ) ? ( VREG_25_7 ) : ( n29431 ) ;
assign n29433 =  ( n28616 ) ? ( VREG_25_8 ) : ( n29432 ) ;
assign n29434 =  ( n28615 ) ? ( VREG_25_9 ) : ( n29433 ) ;
assign n29435 =  ( n28614 ) ? ( VREG_25_10 ) : ( n29434 ) ;
assign n29436 =  ( n28613 ) ? ( VREG_25_11 ) : ( n29435 ) ;
assign n29437 =  ( n28612 ) ? ( VREG_25_12 ) : ( n29436 ) ;
assign n29438 =  ( n28611 ) ? ( VREG_25_13 ) : ( n29437 ) ;
assign n29439 =  ( n28610 ) ? ( VREG_25_14 ) : ( n29438 ) ;
assign n29440 =  ( n28609 ) ? ( VREG_25_15 ) : ( n29439 ) ;
assign n29441 =  ( n28608 ) ? ( VREG_26_0 ) : ( n29440 ) ;
assign n29442 =  ( n28607 ) ? ( VREG_26_1 ) : ( n29441 ) ;
assign n29443 =  ( n28606 ) ? ( VREG_26_2 ) : ( n29442 ) ;
assign n29444 =  ( n28605 ) ? ( VREG_26_3 ) : ( n29443 ) ;
assign n29445 =  ( n28604 ) ? ( VREG_26_4 ) : ( n29444 ) ;
assign n29446 =  ( n28603 ) ? ( VREG_26_5 ) : ( n29445 ) ;
assign n29447 =  ( n28602 ) ? ( VREG_26_6 ) : ( n29446 ) ;
assign n29448 =  ( n28601 ) ? ( VREG_26_7 ) : ( n29447 ) ;
assign n29449 =  ( n28600 ) ? ( VREG_26_8 ) : ( n29448 ) ;
assign n29450 =  ( n28599 ) ? ( VREG_26_9 ) : ( n29449 ) ;
assign n29451 =  ( n28598 ) ? ( VREG_26_10 ) : ( n29450 ) ;
assign n29452 =  ( n28597 ) ? ( VREG_26_11 ) : ( n29451 ) ;
assign n29453 =  ( n28596 ) ? ( VREG_26_12 ) : ( n29452 ) ;
assign n29454 =  ( n28595 ) ? ( VREG_26_13 ) : ( n29453 ) ;
assign n29455 =  ( n28594 ) ? ( VREG_26_14 ) : ( n29454 ) ;
assign n29456 =  ( n28593 ) ? ( VREG_26_15 ) : ( n29455 ) ;
assign n29457 =  ( n28592 ) ? ( VREG_27_0 ) : ( n29456 ) ;
assign n29458 =  ( n28591 ) ? ( VREG_27_1 ) : ( n29457 ) ;
assign n29459 =  ( n28590 ) ? ( VREG_27_2 ) : ( n29458 ) ;
assign n29460 =  ( n28589 ) ? ( VREG_27_3 ) : ( n29459 ) ;
assign n29461 =  ( n28588 ) ? ( VREG_27_4 ) : ( n29460 ) ;
assign n29462 =  ( n28587 ) ? ( VREG_27_5 ) : ( n29461 ) ;
assign n29463 =  ( n28586 ) ? ( VREG_27_6 ) : ( n29462 ) ;
assign n29464 =  ( n28585 ) ? ( VREG_27_7 ) : ( n29463 ) ;
assign n29465 =  ( n28584 ) ? ( VREG_27_8 ) : ( n29464 ) ;
assign n29466 =  ( n28583 ) ? ( VREG_27_9 ) : ( n29465 ) ;
assign n29467 =  ( n28582 ) ? ( VREG_27_10 ) : ( n29466 ) ;
assign n29468 =  ( n28581 ) ? ( VREG_27_11 ) : ( n29467 ) ;
assign n29469 =  ( n28580 ) ? ( VREG_27_12 ) : ( n29468 ) ;
assign n29470 =  ( n28579 ) ? ( VREG_27_13 ) : ( n29469 ) ;
assign n29471 =  ( n28578 ) ? ( VREG_27_14 ) : ( n29470 ) ;
assign n29472 =  ( n28577 ) ? ( VREG_27_15 ) : ( n29471 ) ;
assign n29473 =  ( n28576 ) ? ( VREG_28_0 ) : ( n29472 ) ;
assign n29474 =  ( n28575 ) ? ( VREG_28_1 ) : ( n29473 ) ;
assign n29475 =  ( n28574 ) ? ( VREG_28_2 ) : ( n29474 ) ;
assign n29476 =  ( n28573 ) ? ( VREG_28_3 ) : ( n29475 ) ;
assign n29477 =  ( n28572 ) ? ( VREG_28_4 ) : ( n29476 ) ;
assign n29478 =  ( n28571 ) ? ( VREG_28_5 ) : ( n29477 ) ;
assign n29479 =  ( n28570 ) ? ( VREG_28_6 ) : ( n29478 ) ;
assign n29480 =  ( n28569 ) ? ( VREG_28_7 ) : ( n29479 ) ;
assign n29481 =  ( n28568 ) ? ( VREG_28_8 ) : ( n29480 ) ;
assign n29482 =  ( n28567 ) ? ( VREG_28_9 ) : ( n29481 ) ;
assign n29483 =  ( n28566 ) ? ( VREG_28_10 ) : ( n29482 ) ;
assign n29484 =  ( n28565 ) ? ( VREG_28_11 ) : ( n29483 ) ;
assign n29485 =  ( n28564 ) ? ( VREG_28_12 ) : ( n29484 ) ;
assign n29486 =  ( n28563 ) ? ( VREG_28_13 ) : ( n29485 ) ;
assign n29487 =  ( n28562 ) ? ( VREG_28_14 ) : ( n29486 ) ;
assign n29488 =  ( n28561 ) ? ( VREG_28_15 ) : ( n29487 ) ;
assign n29489 =  ( n28560 ) ? ( VREG_29_0 ) : ( n29488 ) ;
assign n29490 =  ( n28559 ) ? ( VREG_29_1 ) : ( n29489 ) ;
assign n29491 =  ( n28558 ) ? ( VREG_29_2 ) : ( n29490 ) ;
assign n29492 =  ( n28557 ) ? ( VREG_29_3 ) : ( n29491 ) ;
assign n29493 =  ( n28556 ) ? ( VREG_29_4 ) : ( n29492 ) ;
assign n29494 =  ( n28555 ) ? ( VREG_29_5 ) : ( n29493 ) ;
assign n29495 =  ( n28554 ) ? ( VREG_29_6 ) : ( n29494 ) ;
assign n29496 =  ( n28553 ) ? ( VREG_29_7 ) : ( n29495 ) ;
assign n29497 =  ( n28552 ) ? ( VREG_29_8 ) : ( n29496 ) ;
assign n29498 =  ( n28551 ) ? ( VREG_29_9 ) : ( n29497 ) ;
assign n29499 =  ( n28550 ) ? ( VREG_29_10 ) : ( n29498 ) ;
assign n29500 =  ( n28549 ) ? ( VREG_29_11 ) : ( n29499 ) ;
assign n29501 =  ( n28548 ) ? ( VREG_29_12 ) : ( n29500 ) ;
assign n29502 =  ( n28547 ) ? ( VREG_29_13 ) : ( n29501 ) ;
assign n29503 =  ( n28546 ) ? ( VREG_29_14 ) : ( n29502 ) ;
assign n29504 =  ( n28545 ) ? ( VREG_29_15 ) : ( n29503 ) ;
assign n29505 =  ( n28544 ) ? ( VREG_30_0 ) : ( n29504 ) ;
assign n29506 =  ( n28543 ) ? ( VREG_30_1 ) : ( n29505 ) ;
assign n29507 =  ( n28542 ) ? ( VREG_30_2 ) : ( n29506 ) ;
assign n29508 =  ( n28541 ) ? ( VREG_30_3 ) : ( n29507 ) ;
assign n29509 =  ( n28540 ) ? ( VREG_30_4 ) : ( n29508 ) ;
assign n29510 =  ( n28539 ) ? ( VREG_30_5 ) : ( n29509 ) ;
assign n29511 =  ( n28538 ) ? ( VREG_30_6 ) : ( n29510 ) ;
assign n29512 =  ( n28537 ) ? ( VREG_30_7 ) : ( n29511 ) ;
assign n29513 =  ( n28536 ) ? ( VREG_30_8 ) : ( n29512 ) ;
assign n29514 =  ( n28535 ) ? ( VREG_30_9 ) : ( n29513 ) ;
assign n29515 =  ( n28534 ) ? ( VREG_30_10 ) : ( n29514 ) ;
assign n29516 =  ( n28533 ) ? ( VREG_30_11 ) : ( n29515 ) ;
assign n29517 =  ( n28532 ) ? ( VREG_30_12 ) : ( n29516 ) ;
assign n29518 =  ( n28531 ) ? ( VREG_30_13 ) : ( n29517 ) ;
assign n29519 =  ( n28530 ) ? ( VREG_30_14 ) : ( n29518 ) ;
assign n29520 =  ( n28529 ) ? ( VREG_30_15 ) : ( n29519 ) ;
assign n29521 =  ( n28528 ) ? ( VREG_31_0 ) : ( n29520 ) ;
assign n29522 =  ( n28526 ) ? ( VREG_31_1 ) : ( n29521 ) ;
assign n29523 =  ( n28524 ) ? ( VREG_31_2 ) : ( n29522 ) ;
assign n29524 =  ( n28522 ) ? ( VREG_31_3 ) : ( n29523 ) ;
assign n29525 =  ( n28520 ) ? ( VREG_31_4 ) : ( n29524 ) ;
assign n29526 =  ( n28518 ) ? ( VREG_31_5 ) : ( n29525 ) ;
assign n29527 =  ( n28516 ) ? ( VREG_31_6 ) : ( n29526 ) ;
assign n29528 =  ( n28514 ) ? ( VREG_31_7 ) : ( n29527 ) ;
assign n29529 =  ( n28512 ) ? ( VREG_31_8 ) : ( n29528 ) ;
assign n29530 =  ( n28510 ) ? ( VREG_31_9 ) : ( n29529 ) ;
assign n29531 =  ( n28508 ) ? ( VREG_31_10 ) : ( n29530 ) ;
assign n29532 =  ( n28506 ) ? ( VREG_31_11 ) : ( n29531 ) ;
assign n29533 =  ( n28504 ) ? ( VREG_31_12 ) : ( n29532 ) ;
assign n29534 =  ( n28502 ) ? ( VREG_31_13 ) : ( n29533 ) ;
assign n29535 =  ( n28500 ) ? ( VREG_31_14 ) : ( n29534 ) ;
assign n29536 =  ( n28498 ) ? ( VREG_31_15 ) : ( n29535 ) ;
assign n29537 =  ( n29536 ) + ( n140 )  ;
assign n29538 =  ( n29536 ) - ( n140 )  ;
assign n29539 =  ( n29536 ) & ( n140 )  ;
assign n29540 =  ( n29536 ) | ( n140 )  ;
assign n29541 =  ( ( n29536 ) * ( n140 ))  ;
assign n29542 =  ( n148 ) ? ( n29541 ) : ( VREG_0_7 ) ;
assign n29543 =  ( n146 ) ? ( n29540 ) : ( n29542 ) ;
assign n29544 =  ( n144 ) ? ( n29539 ) : ( n29543 ) ;
assign n29545 =  ( n142 ) ? ( n29538 ) : ( n29544 ) ;
assign n29546 =  ( n10 ) ? ( n29537 ) : ( n29545 ) ;
assign n29547 =  ( n77 ) & ( n28497 )  ;
assign n29548 =  ( n77 ) & ( n28499 )  ;
assign n29549 =  ( n77 ) & ( n28501 )  ;
assign n29550 =  ( n77 ) & ( n28503 )  ;
assign n29551 =  ( n77 ) & ( n28505 )  ;
assign n29552 =  ( n77 ) & ( n28507 )  ;
assign n29553 =  ( n77 ) & ( n28509 )  ;
assign n29554 =  ( n77 ) & ( n28511 )  ;
assign n29555 =  ( n77 ) & ( n28513 )  ;
assign n29556 =  ( n77 ) & ( n28515 )  ;
assign n29557 =  ( n77 ) & ( n28517 )  ;
assign n29558 =  ( n77 ) & ( n28519 )  ;
assign n29559 =  ( n77 ) & ( n28521 )  ;
assign n29560 =  ( n77 ) & ( n28523 )  ;
assign n29561 =  ( n77 ) & ( n28525 )  ;
assign n29562 =  ( n77 ) & ( n28527 )  ;
assign n29563 =  ( n78 ) & ( n28497 )  ;
assign n29564 =  ( n78 ) & ( n28499 )  ;
assign n29565 =  ( n78 ) & ( n28501 )  ;
assign n29566 =  ( n78 ) & ( n28503 )  ;
assign n29567 =  ( n78 ) & ( n28505 )  ;
assign n29568 =  ( n78 ) & ( n28507 )  ;
assign n29569 =  ( n78 ) & ( n28509 )  ;
assign n29570 =  ( n78 ) & ( n28511 )  ;
assign n29571 =  ( n78 ) & ( n28513 )  ;
assign n29572 =  ( n78 ) & ( n28515 )  ;
assign n29573 =  ( n78 ) & ( n28517 )  ;
assign n29574 =  ( n78 ) & ( n28519 )  ;
assign n29575 =  ( n78 ) & ( n28521 )  ;
assign n29576 =  ( n78 ) & ( n28523 )  ;
assign n29577 =  ( n78 ) & ( n28525 )  ;
assign n29578 =  ( n78 ) & ( n28527 )  ;
assign n29579 =  ( n79 ) & ( n28497 )  ;
assign n29580 =  ( n79 ) & ( n28499 )  ;
assign n29581 =  ( n79 ) & ( n28501 )  ;
assign n29582 =  ( n79 ) & ( n28503 )  ;
assign n29583 =  ( n79 ) & ( n28505 )  ;
assign n29584 =  ( n79 ) & ( n28507 )  ;
assign n29585 =  ( n79 ) & ( n28509 )  ;
assign n29586 =  ( n79 ) & ( n28511 )  ;
assign n29587 =  ( n79 ) & ( n28513 )  ;
assign n29588 =  ( n79 ) & ( n28515 )  ;
assign n29589 =  ( n79 ) & ( n28517 )  ;
assign n29590 =  ( n79 ) & ( n28519 )  ;
assign n29591 =  ( n79 ) & ( n28521 )  ;
assign n29592 =  ( n79 ) & ( n28523 )  ;
assign n29593 =  ( n79 ) & ( n28525 )  ;
assign n29594 =  ( n79 ) & ( n28527 )  ;
assign n29595 =  ( n80 ) & ( n28497 )  ;
assign n29596 =  ( n80 ) & ( n28499 )  ;
assign n29597 =  ( n80 ) & ( n28501 )  ;
assign n29598 =  ( n80 ) & ( n28503 )  ;
assign n29599 =  ( n80 ) & ( n28505 )  ;
assign n29600 =  ( n80 ) & ( n28507 )  ;
assign n29601 =  ( n80 ) & ( n28509 )  ;
assign n29602 =  ( n80 ) & ( n28511 )  ;
assign n29603 =  ( n80 ) & ( n28513 )  ;
assign n29604 =  ( n80 ) & ( n28515 )  ;
assign n29605 =  ( n80 ) & ( n28517 )  ;
assign n29606 =  ( n80 ) & ( n28519 )  ;
assign n29607 =  ( n80 ) & ( n28521 )  ;
assign n29608 =  ( n80 ) & ( n28523 )  ;
assign n29609 =  ( n80 ) & ( n28525 )  ;
assign n29610 =  ( n80 ) & ( n28527 )  ;
assign n29611 =  ( n81 ) & ( n28497 )  ;
assign n29612 =  ( n81 ) & ( n28499 )  ;
assign n29613 =  ( n81 ) & ( n28501 )  ;
assign n29614 =  ( n81 ) & ( n28503 )  ;
assign n29615 =  ( n81 ) & ( n28505 )  ;
assign n29616 =  ( n81 ) & ( n28507 )  ;
assign n29617 =  ( n81 ) & ( n28509 )  ;
assign n29618 =  ( n81 ) & ( n28511 )  ;
assign n29619 =  ( n81 ) & ( n28513 )  ;
assign n29620 =  ( n81 ) & ( n28515 )  ;
assign n29621 =  ( n81 ) & ( n28517 )  ;
assign n29622 =  ( n81 ) & ( n28519 )  ;
assign n29623 =  ( n81 ) & ( n28521 )  ;
assign n29624 =  ( n81 ) & ( n28523 )  ;
assign n29625 =  ( n81 ) & ( n28525 )  ;
assign n29626 =  ( n81 ) & ( n28527 )  ;
assign n29627 =  ( n82 ) & ( n28497 )  ;
assign n29628 =  ( n82 ) & ( n28499 )  ;
assign n29629 =  ( n82 ) & ( n28501 )  ;
assign n29630 =  ( n82 ) & ( n28503 )  ;
assign n29631 =  ( n82 ) & ( n28505 )  ;
assign n29632 =  ( n82 ) & ( n28507 )  ;
assign n29633 =  ( n82 ) & ( n28509 )  ;
assign n29634 =  ( n82 ) & ( n28511 )  ;
assign n29635 =  ( n82 ) & ( n28513 )  ;
assign n29636 =  ( n82 ) & ( n28515 )  ;
assign n29637 =  ( n82 ) & ( n28517 )  ;
assign n29638 =  ( n82 ) & ( n28519 )  ;
assign n29639 =  ( n82 ) & ( n28521 )  ;
assign n29640 =  ( n82 ) & ( n28523 )  ;
assign n29641 =  ( n82 ) & ( n28525 )  ;
assign n29642 =  ( n82 ) & ( n28527 )  ;
assign n29643 =  ( n83 ) & ( n28497 )  ;
assign n29644 =  ( n83 ) & ( n28499 )  ;
assign n29645 =  ( n83 ) & ( n28501 )  ;
assign n29646 =  ( n83 ) & ( n28503 )  ;
assign n29647 =  ( n83 ) & ( n28505 )  ;
assign n29648 =  ( n83 ) & ( n28507 )  ;
assign n29649 =  ( n83 ) & ( n28509 )  ;
assign n29650 =  ( n83 ) & ( n28511 )  ;
assign n29651 =  ( n83 ) & ( n28513 )  ;
assign n29652 =  ( n83 ) & ( n28515 )  ;
assign n29653 =  ( n83 ) & ( n28517 )  ;
assign n29654 =  ( n83 ) & ( n28519 )  ;
assign n29655 =  ( n83 ) & ( n28521 )  ;
assign n29656 =  ( n83 ) & ( n28523 )  ;
assign n29657 =  ( n83 ) & ( n28525 )  ;
assign n29658 =  ( n83 ) & ( n28527 )  ;
assign n29659 =  ( n84 ) & ( n28497 )  ;
assign n29660 =  ( n84 ) & ( n28499 )  ;
assign n29661 =  ( n84 ) & ( n28501 )  ;
assign n29662 =  ( n84 ) & ( n28503 )  ;
assign n29663 =  ( n84 ) & ( n28505 )  ;
assign n29664 =  ( n84 ) & ( n28507 )  ;
assign n29665 =  ( n84 ) & ( n28509 )  ;
assign n29666 =  ( n84 ) & ( n28511 )  ;
assign n29667 =  ( n84 ) & ( n28513 )  ;
assign n29668 =  ( n84 ) & ( n28515 )  ;
assign n29669 =  ( n84 ) & ( n28517 )  ;
assign n29670 =  ( n84 ) & ( n28519 )  ;
assign n29671 =  ( n84 ) & ( n28521 )  ;
assign n29672 =  ( n84 ) & ( n28523 )  ;
assign n29673 =  ( n84 ) & ( n28525 )  ;
assign n29674 =  ( n84 ) & ( n28527 )  ;
assign n29675 =  ( n85 ) & ( n28497 )  ;
assign n29676 =  ( n85 ) & ( n28499 )  ;
assign n29677 =  ( n85 ) & ( n28501 )  ;
assign n29678 =  ( n85 ) & ( n28503 )  ;
assign n29679 =  ( n85 ) & ( n28505 )  ;
assign n29680 =  ( n85 ) & ( n28507 )  ;
assign n29681 =  ( n85 ) & ( n28509 )  ;
assign n29682 =  ( n85 ) & ( n28511 )  ;
assign n29683 =  ( n85 ) & ( n28513 )  ;
assign n29684 =  ( n85 ) & ( n28515 )  ;
assign n29685 =  ( n85 ) & ( n28517 )  ;
assign n29686 =  ( n85 ) & ( n28519 )  ;
assign n29687 =  ( n85 ) & ( n28521 )  ;
assign n29688 =  ( n85 ) & ( n28523 )  ;
assign n29689 =  ( n85 ) & ( n28525 )  ;
assign n29690 =  ( n85 ) & ( n28527 )  ;
assign n29691 =  ( n86 ) & ( n28497 )  ;
assign n29692 =  ( n86 ) & ( n28499 )  ;
assign n29693 =  ( n86 ) & ( n28501 )  ;
assign n29694 =  ( n86 ) & ( n28503 )  ;
assign n29695 =  ( n86 ) & ( n28505 )  ;
assign n29696 =  ( n86 ) & ( n28507 )  ;
assign n29697 =  ( n86 ) & ( n28509 )  ;
assign n29698 =  ( n86 ) & ( n28511 )  ;
assign n29699 =  ( n86 ) & ( n28513 )  ;
assign n29700 =  ( n86 ) & ( n28515 )  ;
assign n29701 =  ( n86 ) & ( n28517 )  ;
assign n29702 =  ( n86 ) & ( n28519 )  ;
assign n29703 =  ( n86 ) & ( n28521 )  ;
assign n29704 =  ( n86 ) & ( n28523 )  ;
assign n29705 =  ( n86 ) & ( n28525 )  ;
assign n29706 =  ( n86 ) & ( n28527 )  ;
assign n29707 =  ( n87 ) & ( n28497 )  ;
assign n29708 =  ( n87 ) & ( n28499 )  ;
assign n29709 =  ( n87 ) & ( n28501 )  ;
assign n29710 =  ( n87 ) & ( n28503 )  ;
assign n29711 =  ( n87 ) & ( n28505 )  ;
assign n29712 =  ( n87 ) & ( n28507 )  ;
assign n29713 =  ( n87 ) & ( n28509 )  ;
assign n29714 =  ( n87 ) & ( n28511 )  ;
assign n29715 =  ( n87 ) & ( n28513 )  ;
assign n29716 =  ( n87 ) & ( n28515 )  ;
assign n29717 =  ( n87 ) & ( n28517 )  ;
assign n29718 =  ( n87 ) & ( n28519 )  ;
assign n29719 =  ( n87 ) & ( n28521 )  ;
assign n29720 =  ( n87 ) & ( n28523 )  ;
assign n29721 =  ( n87 ) & ( n28525 )  ;
assign n29722 =  ( n87 ) & ( n28527 )  ;
assign n29723 =  ( n88 ) & ( n28497 )  ;
assign n29724 =  ( n88 ) & ( n28499 )  ;
assign n29725 =  ( n88 ) & ( n28501 )  ;
assign n29726 =  ( n88 ) & ( n28503 )  ;
assign n29727 =  ( n88 ) & ( n28505 )  ;
assign n29728 =  ( n88 ) & ( n28507 )  ;
assign n29729 =  ( n88 ) & ( n28509 )  ;
assign n29730 =  ( n88 ) & ( n28511 )  ;
assign n29731 =  ( n88 ) & ( n28513 )  ;
assign n29732 =  ( n88 ) & ( n28515 )  ;
assign n29733 =  ( n88 ) & ( n28517 )  ;
assign n29734 =  ( n88 ) & ( n28519 )  ;
assign n29735 =  ( n88 ) & ( n28521 )  ;
assign n29736 =  ( n88 ) & ( n28523 )  ;
assign n29737 =  ( n88 ) & ( n28525 )  ;
assign n29738 =  ( n88 ) & ( n28527 )  ;
assign n29739 =  ( n89 ) & ( n28497 )  ;
assign n29740 =  ( n89 ) & ( n28499 )  ;
assign n29741 =  ( n89 ) & ( n28501 )  ;
assign n29742 =  ( n89 ) & ( n28503 )  ;
assign n29743 =  ( n89 ) & ( n28505 )  ;
assign n29744 =  ( n89 ) & ( n28507 )  ;
assign n29745 =  ( n89 ) & ( n28509 )  ;
assign n29746 =  ( n89 ) & ( n28511 )  ;
assign n29747 =  ( n89 ) & ( n28513 )  ;
assign n29748 =  ( n89 ) & ( n28515 )  ;
assign n29749 =  ( n89 ) & ( n28517 )  ;
assign n29750 =  ( n89 ) & ( n28519 )  ;
assign n29751 =  ( n89 ) & ( n28521 )  ;
assign n29752 =  ( n89 ) & ( n28523 )  ;
assign n29753 =  ( n89 ) & ( n28525 )  ;
assign n29754 =  ( n89 ) & ( n28527 )  ;
assign n29755 =  ( n90 ) & ( n28497 )  ;
assign n29756 =  ( n90 ) & ( n28499 )  ;
assign n29757 =  ( n90 ) & ( n28501 )  ;
assign n29758 =  ( n90 ) & ( n28503 )  ;
assign n29759 =  ( n90 ) & ( n28505 )  ;
assign n29760 =  ( n90 ) & ( n28507 )  ;
assign n29761 =  ( n90 ) & ( n28509 )  ;
assign n29762 =  ( n90 ) & ( n28511 )  ;
assign n29763 =  ( n90 ) & ( n28513 )  ;
assign n29764 =  ( n90 ) & ( n28515 )  ;
assign n29765 =  ( n90 ) & ( n28517 )  ;
assign n29766 =  ( n90 ) & ( n28519 )  ;
assign n29767 =  ( n90 ) & ( n28521 )  ;
assign n29768 =  ( n90 ) & ( n28523 )  ;
assign n29769 =  ( n90 ) & ( n28525 )  ;
assign n29770 =  ( n90 ) & ( n28527 )  ;
assign n29771 =  ( n91 ) & ( n28497 )  ;
assign n29772 =  ( n91 ) & ( n28499 )  ;
assign n29773 =  ( n91 ) & ( n28501 )  ;
assign n29774 =  ( n91 ) & ( n28503 )  ;
assign n29775 =  ( n91 ) & ( n28505 )  ;
assign n29776 =  ( n91 ) & ( n28507 )  ;
assign n29777 =  ( n91 ) & ( n28509 )  ;
assign n29778 =  ( n91 ) & ( n28511 )  ;
assign n29779 =  ( n91 ) & ( n28513 )  ;
assign n29780 =  ( n91 ) & ( n28515 )  ;
assign n29781 =  ( n91 ) & ( n28517 )  ;
assign n29782 =  ( n91 ) & ( n28519 )  ;
assign n29783 =  ( n91 ) & ( n28521 )  ;
assign n29784 =  ( n91 ) & ( n28523 )  ;
assign n29785 =  ( n91 ) & ( n28525 )  ;
assign n29786 =  ( n91 ) & ( n28527 )  ;
assign n29787 =  ( n92 ) & ( n28497 )  ;
assign n29788 =  ( n92 ) & ( n28499 )  ;
assign n29789 =  ( n92 ) & ( n28501 )  ;
assign n29790 =  ( n92 ) & ( n28503 )  ;
assign n29791 =  ( n92 ) & ( n28505 )  ;
assign n29792 =  ( n92 ) & ( n28507 )  ;
assign n29793 =  ( n92 ) & ( n28509 )  ;
assign n29794 =  ( n92 ) & ( n28511 )  ;
assign n29795 =  ( n92 ) & ( n28513 )  ;
assign n29796 =  ( n92 ) & ( n28515 )  ;
assign n29797 =  ( n92 ) & ( n28517 )  ;
assign n29798 =  ( n92 ) & ( n28519 )  ;
assign n29799 =  ( n92 ) & ( n28521 )  ;
assign n29800 =  ( n92 ) & ( n28523 )  ;
assign n29801 =  ( n92 ) & ( n28525 )  ;
assign n29802 =  ( n92 ) & ( n28527 )  ;
assign n29803 =  ( n93 ) & ( n28497 )  ;
assign n29804 =  ( n93 ) & ( n28499 )  ;
assign n29805 =  ( n93 ) & ( n28501 )  ;
assign n29806 =  ( n93 ) & ( n28503 )  ;
assign n29807 =  ( n93 ) & ( n28505 )  ;
assign n29808 =  ( n93 ) & ( n28507 )  ;
assign n29809 =  ( n93 ) & ( n28509 )  ;
assign n29810 =  ( n93 ) & ( n28511 )  ;
assign n29811 =  ( n93 ) & ( n28513 )  ;
assign n29812 =  ( n93 ) & ( n28515 )  ;
assign n29813 =  ( n93 ) & ( n28517 )  ;
assign n29814 =  ( n93 ) & ( n28519 )  ;
assign n29815 =  ( n93 ) & ( n28521 )  ;
assign n29816 =  ( n93 ) & ( n28523 )  ;
assign n29817 =  ( n93 ) & ( n28525 )  ;
assign n29818 =  ( n93 ) & ( n28527 )  ;
assign n29819 =  ( n94 ) & ( n28497 )  ;
assign n29820 =  ( n94 ) & ( n28499 )  ;
assign n29821 =  ( n94 ) & ( n28501 )  ;
assign n29822 =  ( n94 ) & ( n28503 )  ;
assign n29823 =  ( n94 ) & ( n28505 )  ;
assign n29824 =  ( n94 ) & ( n28507 )  ;
assign n29825 =  ( n94 ) & ( n28509 )  ;
assign n29826 =  ( n94 ) & ( n28511 )  ;
assign n29827 =  ( n94 ) & ( n28513 )  ;
assign n29828 =  ( n94 ) & ( n28515 )  ;
assign n29829 =  ( n94 ) & ( n28517 )  ;
assign n29830 =  ( n94 ) & ( n28519 )  ;
assign n29831 =  ( n94 ) & ( n28521 )  ;
assign n29832 =  ( n94 ) & ( n28523 )  ;
assign n29833 =  ( n94 ) & ( n28525 )  ;
assign n29834 =  ( n94 ) & ( n28527 )  ;
assign n29835 =  ( n95 ) & ( n28497 )  ;
assign n29836 =  ( n95 ) & ( n28499 )  ;
assign n29837 =  ( n95 ) & ( n28501 )  ;
assign n29838 =  ( n95 ) & ( n28503 )  ;
assign n29839 =  ( n95 ) & ( n28505 )  ;
assign n29840 =  ( n95 ) & ( n28507 )  ;
assign n29841 =  ( n95 ) & ( n28509 )  ;
assign n29842 =  ( n95 ) & ( n28511 )  ;
assign n29843 =  ( n95 ) & ( n28513 )  ;
assign n29844 =  ( n95 ) & ( n28515 )  ;
assign n29845 =  ( n95 ) & ( n28517 )  ;
assign n29846 =  ( n95 ) & ( n28519 )  ;
assign n29847 =  ( n95 ) & ( n28521 )  ;
assign n29848 =  ( n95 ) & ( n28523 )  ;
assign n29849 =  ( n95 ) & ( n28525 )  ;
assign n29850 =  ( n95 ) & ( n28527 )  ;
assign n29851 =  ( n96 ) & ( n28497 )  ;
assign n29852 =  ( n96 ) & ( n28499 )  ;
assign n29853 =  ( n96 ) & ( n28501 )  ;
assign n29854 =  ( n96 ) & ( n28503 )  ;
assign n29855 =  ( n96 ) & ( n28505 )  ;
assign n29856 =  ( n96 ) & ( n28507 )  ;
assign n29857 =  ( n96 ) & ( n28509 )  ;
assign n29858 =  ( n96 ) & ( n28511 )  ;
assign n29859 =  ( n96 ) & ( n28513 )  ;
assign n29860 =  ( n96 ) & ( n28515 )  ;
assign n29861 =  ( n96 ) & ( n28517 )  ;
assign n29862 =  ( n96 ) & ( n28519 )  ;
assign n29863 =  ( n96 ) & ( n28521 )  ;
assign n29864 =  ( n96 ) & ( n28523 )  ;
assign n29865 =  ( n96 ) & ( n28525 )  ;
assign n29866 =  ( n96 ) & ( n28527 )  ;
assign n29867 =  ( n97 ) & ( n28497 )  ;
assign n29868 =  ( n97 ) & ( n28499 )  ;
assign n29869 =  ( n97 ) & ( n28501 )  ;
assign n29870 =  ( n97 ) & ( n28503 )  ;
assign n29871 =  ( n97 ) & ( n28505 )  ;
assign n29872 =  ( n97 ) & ( n28507 )  ;
assign n29873 =  ( n97 ) & ( n28509 )  ;
assign n29874 =  ( n97 ) & ( n28511 )  ;
assign n29875 =  ( n97 ) & ( n28513 )  ;
assign n29876 =  ( n97 ) & ( n28515 )  ;
assign n29877 =  ( n97 ) & ( n28517 )  ;
assign n29878 =  ( n97 ) & ( n28519 )  ;
assign n29879 =  ( n97 ) & ( n28521 )  ;
assign n29880 =  ( n97 ) & ( n28523 )  ;
assign n29881 =  ( n97 ) & ( n28525 )  ;
assign n29882 =  ( n97 ) & ( n28527 )  ;
assign n29883 =  ( n98 ) & ( n28497 )  ;
assign n29884 =  ( n98 ) & ( n28499 )  ;
assign n29885 =  ( n98 ) & ( n28501 )  ;
assign n29886 =  ( n98 ) & ( n28503 )  ;
assign n29887 =  ( n98 ) & ( n28505 )  ;
assign n29888 =  ( n98 ) & ( n28507 )  ;
assign n29889 =  ( n98 ) & ( n28509 )  ;
assign n29890 =  ( n98 ) & ( n28511 )  ;
assign n29891 =  ( n98 ) & ( n28513 )  ;
assign n29892 =  ( n98 ) & ( n28515 )  ;
assign n29893 =  ( n98 ) & ( n28517 )  ;
assign n29894 =  ( n98 ) & ( n28519 )  ;
assign n29895 =  ( n98 ) & ( n28521 )  ;
assign n29896 =  ( n98 ) & ( n28523 )  ;
assign n29897 =  ( n98 ) & ( n28525 )  ;
assign n29898 =  ( n98 ) & ( n28527 )  ;
assign n29899 =  ( n99 ) & ( n28497 )  ;
assign n29900 =  ( n99 ) & ( n28499 )  ;
assign n29901 =  ( n99 ) & ( n28501 )  ;
assign n29902 =  ( n99 ) & ( n28503 )  ;
assign n29903 =  ( n99 ) & ( n28505 )  ;
assign n29904 =  ( n99 ) & ( n28507 )  ;
assign n29905 =  ( n99 ) & ( n28509 )  ;
assign n29906 =  ( n99 ) & ( n28511 )  ;
assign n29907 =  ( n99 ) & ( n28513 )  ;
assign n29908 =  ( n99 ) & ( n28515 )  ;
assign n29909 =  ( n99 ) & ( n28517 )  ;
assign n29910 =  ( n99 ) & ( n28519 )  ;
assign n29911 =  ( n99 ) & ( n28521 )  ;
assign n29912 =  ( n99 ) & ( n28523 )  ;
assign n29913 =  ( n99 ) & ( n28525 )  ;
assign n29914 =  ( n99 ) & ( n28527 )  ;
assign n29915 =  ( n100 ) & ( n28497 )  ;
assign n29916 =  ( n100 ) & ( n28499 )  ;
assign n29917 =  ( n100 ) & ( n28501 )  ;
assign n29918 =  ( n100 ) & ( n28503 )  ;
assign n29919 =  ( n100 ) & ( n28505 )  ;
assign n29920 =  ( n100 ) & ( n28507 )  ;
assign n29921 =  ( n100 ) & ( n28509 )  ;
assign n29922 =  ( n100 ) & ( n28511 )  ;
assign n29923 =  ( n100 ) & ( n28513 )  ;
assign n29924 =  ( n100 ) & ( n28515 )  ;
assign n29925 =  ( n100 ) & ( n28517 )  ;
assign n29926 =  ( n100 ) & ( n28519 )  ;
assign n29927 =  ( n100 ) & ( n28521 )  ;
assign n29928 =  ( n100 ) & ( n28523 )  ;
assign n29929 =  ( n100 ) & ( n28525 )  ;
assign n29930 =  ( n100 ) & ( n28527 )  ;
assign n29931 =  ( n101 ) & ( n28497 )  ;
assign n29932 =  ( n101 ) & ( n28499 )  ;
assign n29933 =  ( n101 ) & ( n28501 )  ;
assign n29934 =  ( n101 ) & ( n28503 )  ;
assign n29935 =  ( n101 ) & ( n28505 )  ;
assign n29936 =  ( n101 ) & ( n28507 )  ;
assign n29937 =  ( n101 ) & ( n28509 )  ;
assign n29938 =  ( n101 ) & ( n28511 )  ;
assign n29939 =  ( n101 ) & ( n28513 )  ;
assign n29940 =  ( n101 ) & ( n28515 )  ;
assign n29941 =  ( n101 ) & ( n28517 )  ;
assign n29942 =  ( n101 ) & ( n28519 )  ;
assign n29943 =  ( n101 ) & ( n28521 )  ;
assign n29944 =  ( n101 ) & ( n28523 )  ;
assign n29945 =  ( n101 ) & ( n28525 )  ;
assign n29946 =  ( n101 ) & ( n28527 )  ;
assign n29947 =  ( n102 ) & ( n28497 )  ;
assign n29948 =  ( n102 ) & ( n28499 )  ;
assign n29949 =  ( n102 ) & ( n28501 )  ;
assign n29950 =  ( n102 ) & ( n28503 )  ;
assign n29951 =  ( n102 ) & ( n28505 )  ;
assign n29952 =  ( n102 ) & ( n28507 )  ;
assign n29953 =  ( n102 ) & ( n28509 )  ;
assign n29954 =  ( n102 ) & ( n28511 )  ;
assign n29955 =  ( n102 ) & ( n28513 )  ;
assign n29956 =  ( n102 ) & ( n28515 )  ;
assign n29957 =  ( n102 ) & ( n28517 )  ;
assign n29958 =  ( n102 ) & ( n28519 )  ;
assign n29959 =  ( n102 ) & ( n28521 )  ;
assign n29960 =  ( n102 ) & ( n28523 )  ;
assign n29961 =  ( n102 ) & ( n28525 )  ;
assign n29962 =  ( n102 ) & ( n28527 )  ;
assign n29963 =  ( n103 ) & ( n28497 )  ;
assign n29964 =  ( n103 ) & ( n28499 )  ;
assign n29965 =  ( n103 ) & ( n28501 )  ;
assign n29966 =  ( n103 ) & ( n28503 )  ;
assign n29967 =  ( n103 ) & ( n28505 )  ;
assign n29968 =  ( n103 ) & ( n28507 )  ;
assign n29969 =  ( n103 ) & ( n28509 )  ;
assign n29970 =  ( n103 ) & ( n28511 )  ;
assign n29971 =  ( n103 ) & ( n28513 )  ;
assign n29972 =  ( n103 ) & ( n28515 )  ;
assign n29973 =  ( n103 ) & ( n28517 )  ;
assign n29974 =  ( n103 ) & ( n28519 )  ;
assign n29975 =  ( n103 ) & ( n28521 )  ;
assign n29976 =  ( n103 ) & ( n28523 )  ;
assign n29977 =  ( n103 ) & ( n28525 )  ;
assign n29978 =  ( n103 ) & ( n28527 )  ;
assign n29979 =  ( n104 ) & ( n28497 )  ;
assign n29980 =  ( n104 ) & ( n28499 )  ;
assign n29981 =  ( n104 ) & ( n28501 )  ;
assign n29982 =  ( n104 ) & ( n28503 )  ;
assign n29983 =  ( n104 ) & ( n28505 )  ;
assign n29984 =  ( n104 ) & ( n28507 )  ;
assign n29985 =  ( n104 ) & ( n28509 )  ;
assign n29986 =  ( n104 ) & ( n28511 )  ;
assign n29987 =  ( n104 ) & ( n28513 )  ;
assign n29988 =  ( n104 ) & ( n28515 )  ;
assign n29989 =  ( n104 ) & ( n28517 )  ;
assign n29990 =  ( n104 ) & ( n28519 )  ;
assign n29991 =  ( n104 ) & ( n28521 )  ;
assign n29992 =  ( n104 ) & ( n28523 )  ;
assign n29993 =  ( n104 ) & ( n28525 )  ;
assign n29994 =  ( n104 ) & ( n28527 )  ;
assign n29995 =  ( n105 ) & ( n28497 )  ;
assign n29996 =  ( n105 ) & ( n28499 )  ;
assign n29997 =  ( n105 ) & ( n28501 )  ;
assign n29998 =  ( n105 ) & ( n28503 )  ;
assign n29999 =  ( n105 ) & ( n28505 )  ;
assign n30000 =  ( n105 ) & ( n28507 )  ;
assign n30001 =  ( n105 ) & ( n28509 )  ;
assign n30002 =  ( n105 ) & ( n28511 )  ;
assign n30003 =  ( n105 ) & ( n28513 )  ;
assign n30004 =  ( n105 ) & ( n28515 )  ;
assign n30005 =  ( n105 ) & ( n28517 )  ;
assign n30006 =  ( n105 ) & ( n28519 )  ;
assign n30007 =  ( n105 ) & ( n28521 )  ;
assign n30008 =  ( n105 ) & ( n28523 )  ;
assign n30009 =  ( n105 ) & ( n28525 )  ;
assign n30010 =  ( n105 ) & ( n28527 )  ;
assign n30011 =  ( n106 ) & ( n28497 )  ;
assign n30012 =  ( n106 ) & ( n28499 )  ;
assign n30013 =  ( n106 ) & ( n28501 )  ;
assign n30014 =  ( n106 ) & ( n28503 )  ;
assign n30015 =  ( n106 ) & ( n28505 )  ;
assign n30016 =  ( n106 ) & ( n28507 )  ;
assign n30017 =  ( n106 ) & ( n28509 )  ;
assign n30018 =  ( n106 ) & ( n28511 )  ;
assign n30019 =  ( n106 ) & ( n28513 )  ;
assign n30020 =  ( n106 ) & ( n28515 )  ;
assign n30021 =  ( n106 ) & ( n28517 )  ;
assign n30022 =  ( n106 ) & ( n28519 )  ;
assign n30023 =  ( n106 ) & ( n28521 )  ;
assign n30024 =  ( n106 ) & ( n28523 )  ;
assign n30025 =  ( n106 ) & ( n28525 )  ;
assign n30026 =  ( n106 ) & ( n28527 )  ;
assign n30027 =  ( n107 ) & ( n28497 )  ;
assign n30028 =  ( n107 ) & ( n28499 )  ;
assign n30029 =  ( n107 ) & ( n28501 )  ;
assign n30030 =  ( n107 ) & ( n28503 )  ;
assign n30031 =  ( n107 ) & ( n28505 )  ;
assign n30032 =  ( n107 ) & ( n28507 )  ;
assign n30033 =  ( n107 ) & ( n28509 )  ;
assign n30034 =  ( n107 ) & ( n28511 )  ;
assign n30035 =  ( n107 ) & ( n28513 )  ;
assign n30036 =  ( n107 ) & ( n28515 )  ;
assign n30037 =  ( n107 ) & ( n28517 )  ;
assign n30038 =  ( n107 ) & ( n28519 )  ;
assign n30039 =  ( n107 ) & ( n28521 )  ;
assign n30040 =  ( n107 ) & ( n28523 )  ;
assign n30041 =  ( n107 ) & ( n28525 )  ;
assign n30042 =  ( n107 ) & ( n28527 )  ;
assign n30043 =  ( n108 ) & ( n28497 )  ;
assign n30044 =  ( n108 ) & ( n28499 )  ;
assign n30045 =  ( n108 ) & ( n28501 )  ;
assign n30046 =  ( n108 ) & ( n28503 )  ;
assign n30047 =  ( n108 ) & ( n28505 )  ;
assign n30048 =  ( n108 ) & ( n28507 )  ;
assign n30049 =  ( n108 ) & ( n28509 )  ;
assign n30050 =  ( n108 ) & ( n28511 )  ;
assign n30051 =  ( n108 ) & ( n28513 )  ;
assign n30052 =  ( n108 ) & ( n28515 )  ;
assign n30053 =  ( n108 ) & ( n28517 )  ;
assign n30054 =  ( n108 ) & ( n28519 )  ;
assign n30055 =  ( n108 ) & ( n28521 )  ;
assign n30056 =  ( n108 ) & ( n28523 )  ;
assign n30057 =  ( n108 ) & ( n28525 )  ;
assign n30058 =  ( n108 ) & ( n28527 )  ;
assign n30059 =  ( n30058 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n30060 =  ( n30057 ) ? ( VREG_0_1 ) : ( n30059 ) ;
assign n30061 =  ( n30056 ) ? ( VREG_0_2 ) : ( n30060 ) ;
assign n30062 =  ( n30055 ) ? ( VREG_0_3 ) : ( n30061 ) ;
assign n30063 =  ( n30054 ) ? ( VREG_0_4 ) : ( n30062 ) ;
assign n30064 =  ( n30053 ) ? ( VREG_0_5 ) : ( n30063 ) ;
assign n30065 =  ( n30052 ) ? ( VREG_0_6 ) : ( n30064 ) ;
assign n30066 =  ( n30051 ) ? ( VREG_0_7 ) : ( n30065 ) ;
assign n30067 =  ( n30050 ) ? ( VREG_0_8 ) : ( n30066 ) ;
assign n30068 =  ( n30049 ) ? ( VREG_0_9 ) : ( n30067 ) ;
assign n30069 =  ( n30048 ) ? ( VREG_0_10 ) : ( n30068 ) ;
assign n30070 =  ( n30047 ) ? ( VREG_0_11 ) : ( n30069 ) ;
assign n30071 =  ( n30046 ) ? ( VREG_0_12 ) : ( n30070 ) ;
assign n30072 =  ( n30045 ) ? ( VREG_0_13 ) : ( n30071 ) ;
assign n30073 =  ( n30044 ) ? ( VREG_0_14 ) : ( n30072 ) ;
assign n30074 =  ( n30043 ) ? ( VREG_0_15 ) : ( n30073 ) ;
assign n30075 =  ( n30042 ) ? ( VREG_1_0 ) : ( n30074 ) ;
assign n30076 =  ( n30041 ) ? ( VREG_1_1 ) : ( n30075 ) ;
assign n30077 =  ( n30040 ) ? ( VREG_1_2 ) : ( n30076 ) ;
assign n30078 =  ( n30039 ) ? ( VREG_1_3 ) : ( n30077 ) ;
assign n30079 =  ( n30038 ) ? ( VREG_1_4 ) : ( n30078 ) ;
assign n30080 =  ( n30037 ) ? ( VREG_1_5 ) : ( n30079 ) ;
assign n30081 =  ( n30036 ) ? ( VREG_1_6 ) : ( n30080 ) ;
assign n30082 =  ( n30035 ) ? ( VREG_1_7 ) : ( n30081 ) ;
assign n30083 =  ( n30034 ) ? ( VREG_1_8 ) : ( n30082 ) ;
assign n30084 =  ( n30033 ) ? ( VREG_1_9 ) : ( n30083 ) ;
assign n30085 =  ( n30032 ) ? ( VREG_1_10 ) : ( n30084 ) ;
assign n30086 =  ( n30031 ) ? ( VREG_1_11 ) : ( n30085 ) ;
assign n30087 =  ( n30030 ) ? ( VREG_1_12 ) : ( n30086 ) ;
assign n30088 =  ( n30029 ) ? ( VREG_1_13 ) : ( n30087 ) ;
assign n30089 =  ( n30028 ) ? ( VREG_1_14 ) : ( n30088 ) ;
assign n30090 =  ( n30027 ) ? ( VREG_1_15 ) : ( n30089 ) ;
assign n30091 =  ( n30026 ) ? ( VREG_2_0 ) : ( n30090 ) ;
assign n30092 =  ( n30025 ) ? ( VREG_2_1 ) : ( n30091 ) ;
assign n30093 =  ( n30024 ) ? ( VREG_2_2 ) : ( n30092 ) ;
assign n30094 =  ( n30023 ) ? ( VREG_2_3 ) : ( n30093 ) ;
assign n30095 =  ( n30022 ) ? ( VREG_2_4 ) : ( n30094 ) ;
assign n30096 =  ( n30021 ) ? ( VREG_2_5 ) : ( n30095 ) ;
assign n30097 =  ( n30020 ) ? ( VREG_2_6 ) : ( n30096 ) ;
assign n30098 =  ( n30019 ) ? ( VREG_2_7 ) : ( n30097 ) ;
assign n30099 =  ( n30018 ) ? ( VREG_2_8 ) : ( n30098 ) ;
assign n30100 =  ( n30017 ) ? ( VREG_2_9 ) : ( n30099 ) ;
assign n30101 =  ( n30016 ) ? ( VREG_2_10 ) : ( n30100 ) ;
assign n30102 =  ( n30015 ) ? ( VREG_2_11 ) : ( n30101 ) ;
assign n30103 =  ( n30014 ) ? ( VREG_2_12 ) : ( n30102 ) ;
assign n30104 =  ( n30013 ) ? ( VREG_2_13 ) : ( n30103 ) ;
assign n30105 =  ( n30012 ) ? ( VREG_2_14 ) : ( n30104 ) ;
assign n30106 =  ( n30011 ) ? ( VREG_2_15 ) : ( n30105 ) ;
assign n30107 =  ( n30010 ) ? ( VREG_3_0 ) : ( n30106 ) ;
assign n30108 =  ( n30009 ) ? ( VREG_3_1 ) : ( n30107 ) ;
assign n30109 =  ( n30008 ) ? ( VREG_3_2 ) : ( n30108 ) ;
assign n30110 =  ( n30007 ) ? ( VREG_3_3 ) : ( n30109 ) ;
assign n30111 =  ( n30006 ) ? ( VREG_3_4 ) : ( n30110 ) ;
assign n30112 =  ( n30005 ) ? ( VREG_3_5 ) : ( n30111 ) ;
assign n30113 =  ( n30004 ) ? ( VREG_3_6 ) : ( n30112 ) ;
assign n30114 =  ( n30003 ) ? ( VREG_3_7 ) : ( n30113 ) ;
assign n30115 =  ( n30002 ) ? ( VREG_3_8 ) : ( n30114 ) ;
assign n30116 =  ( n30001 ) ? ( VREG_3_9 ) : ( n30115 ) ;
assign n30117 =  ( n30000 ) ? ( VREG_3_10 ) : ( n30116 ) ;
assign n30118 =  ( n29999 ) ? ( VREG_3_11 ) : ( n30117 ) ;
assign n30119 =  ( n29998 ) ? ( VREG_3_12 ) : ( n30118 ) ;
assign n30120 =  ( n29997 ) ? ( VREG_3_13 ) : ( n30119 ) ;
assign n30121 =  ( n29996 ) ? ( VREG_3_14 ) : ( n30120 ) ;
assign n30122 =  ( n29995 ) ? ( VREG_3_15 ) : ( n30121 ) ;
assign n30123 =  ( n29994 ) ? ( VREG_4_0 ) : ( n30122 ) ;
assign n30124 =  ( n29993 ) ? ( VREG_4_1 ) : ( n30123 ) ;
assign n30125 =  ( n29992 ) ? ( VREG_4_2 ) : ( n30124 ) ;
assign n30126 =  ( n29991 ) ? ( VREG_4_3 ) : ( n30125 ) ;
assign n30127 =  ( n29990 ) ? ( VREG_4_4 ) : ( n30126 ) ;
assign n30128 =  ( n29989 ) ? ( VREG_4_5 ) : ( n30127 ) ;
assign n30129 =  ( n29988 ) ? ( VREG_4_6 ) : ( n30128 ) ;
assign n30130 =  ( n29987 ) ? ( VREG_4_7 ) : ( n30129 ) ;
assign n30131 =  ( n29986 ) ? ( VREG_4_8 ) : ( n30130 ) ;
assign n30132 =  ( n29985 ) ? ( VREG_4_9 ) : ( n30131 ) ;
assign n30133 =  ( n29984 ) ? ( VREG_4_10 ) : ( n30132 ) ;
assign n30134 =  ( n29983 ) ? ( VREG_4_11 ) : ( n30133 ) ;
assign n30135 =  ( n29982 ) ? ( VREG_4_12 ) : ( n30134 ) ;
assign n30136 =  ( n29981 ) ? ( VREG_4_13 ) : ( n30135 ) ;
assign n30137 =  ( n29980 ) ? ( VREG_4_14 ) : ( n30136 ) ;
assign n30138 =  ( n29979 ) ? ( VREG_4_15 ) : ( n30137 ) ;
assign n30139 =  ( n29978 ) ? ( VREG_5_0 ) : ( n30138 ) ;
assign n30140 =  ( n29977 ) ? ( VREG_5_1 ) : ( n30139 ) ;
assign n30141 =  ( n29976 ) ? ( VREG_5_2 ) : ( n30140 ) ;
assign n30142 =  ( n29975 ) ? ( VREG_5_3 ) : ( n30141 ) ;
assign n30143 =  ( n29974 ) ? ( VREG_5_4 ) : ( n30142 ) ;
assign n30144 =  ( n29973 ) ? ( VREG_5_5 ) : ( n30143 ) ;
assign n30145 =  ( n29972 ) ? ( VREG_5_6 ) : ( n30144 ) ;
assign n30146 =  ( n29971 ) ? ( VREG_5_7 ) : ( n30145 ) ;
assign n30147 =  ( n29970 ) ? ( VREG_5_8 ) : ( n30146 ) ;
assign n30148 =  ( n29969 ) ? ( VREG_5_9 ) : ( n30147 ) ;
assign n30149 =  ( n29968 ) ? ( VREG_5_10 ) : ( n30148 ) ;
assign n30150 =  ( n29967 ) ? ( VREG_5_11 ) : ( n30149 ) ;
assign n30151 =  ( n29966 ) ? ( VREG_5_12 ) : ( n30150 ) ;
assign n30152 =  ( n29965 ) ? ( VREG_5_13 ) : ( n30151 ) ;
assign n30153 =  ( n29964 ) ? ( VREG_5_14 ) : ( n30152 ) ;
assign n30154 =  ( n29963 ) ? ( VREG_5_15 ) : ( n30153 ) ;
assign n30155 =  ( n29962 ) ? ( VREG_6_0 ) : ( n30154 ) ;
assign n30156 =  ( n29961 ) ? ( VREG_6_1 ) : ( n30155 ) ;
assign n30157 =  ( n29960 ) ? ( VREG_6_2 ) : ( n30156 ) ;
assign n30158 =  ( n29959 ) ? ( VREG_6_3 ) : ( n30157 ) ;
assign n30159 =  ( n29958 ) ? ( VREG_6_4 ) : ( n30158 ) ;
assign n30160 =  ( n29957 ) ? ( VREG_6_5 ) : ( n30159 ) ;
assign n30161 =  ( n29956 ) ? ( VREG_6_6 ) : ( n30160 ) ;
assign n30162 =  ( n29955 ) ? ( VREG_6_7 ) : ( n30161 ) ;
assign n30163 =  ( n29954 ) ? ( VREG_6_8 ) : ( n30162 ) ;
assign n30164 =  ( n29953 ) ? ( VREG_6_9 ) : ( n30163 ) ;
assign n30165 =  ( n29952 ) ? ( VREG_6_10 ) : ( n30164 ) ;
assign n30166 =  ( n29951 ) ? ( VREG_6_11 ) : ( n30165 ) ;
assign n30167 =  ( n29950 ) ? ( VREG_6_12 ) : ( n30166 ) ;
assign n30168 =  ( n29949 ) ? ( VREG_6_13 ) : ( n30167 ) ;
assign n30169 =  ( n29948 ) ? ( VREG_6_14 ) : ( n30168 ) ;
assign n30170 =  ( n29947 ) ? ( VREG_6_15 ) : ( n30169 ) ;
assign n30171 =  ( n29946 ) ? ( VREG_7_0 ) : ( n30170 ) ;
assign n30172 =  ( n29945 ) ? ( VREG_7_1 ) : ( n30171 ) ;
assign n30173 =  ( n29944 ) ? ( VREG_7_2 ) : ( n30172 ) ;
assign n30174 =  ( n29943 ) ? ( VREG_7_3 ) : ( n30173 ) ;
assign n30175 =  ( n29942 ) ? ( VREG_7_4 ) : ( n30174 ) ;
assign n30176 =  ( n29941 ) ? ( VREG_7_5 ) : ( n30175 ) ;
assign n30177 =  ( n29940 ) ? ( VREG_7_6 ) : ( n30176 ) ;
assign n30178 =  ( n29939 ) ? ( VREG_7_7 ) : ( n30177 ) ;
assign n30179 =  ( n29938 ) ? ( VREG_7_8 ) : ( n30178 ) ;
assign n30180 =  ( n29937 ) ? ( VREG_7_9 ) : ( n30179 ) ;
assign n30181 =  ( n29936 ) ? ( VREG_7_10 ) : ( n30180 ) ;
assign n30182 =  ( n29935 ) ? ( VREG_7_11 ) : ( n30181 ) ;
assign n30183 =  ( n29934 ) ? ( VREG_7_12 ) : ( n30182 ) ;
assign n30184 =  ( n29933 ) ? ( VREG_7_13 ) : ( n30183 ) ;
assign n30185 =  ( n29932 ) ? ( VREG_7_14 ) : ( n30184 ) ;
assign n30186 =  ( n29931 ) ? ( VREG_7_15 ) : ( n30185 ) ;
assign n30187 =  ( n29930 ) ? ( VREG_8_0 ) : ( n30186 ) ;
assign n30188 =  ( n29929 ) ? ( VREG_8_1 ) : ( n30187 ) ;
assign n30189 =  ( n29928 ) ? ( VREG_8_2 ) : ( n30188 ) ;
assign n30190 =  ( n29927 ) ? ( VREG_8_3 ) : ( n30189 ) ;
assign n30191 =  ( n29926 ) ? ( VREG_8_4 ) : ( n30190 ) ;
assign n30192 =  ( n29925 ) ? ( VREG_8_5 ) : ( n30191 ) ;
assign n30193 =  ( n29924 ) ? ( VREG_8_6 ) : ( n30192 ) ;
assign n30194 =  ( n29923 ) ? ( VREG_8_7 ) : ( n30193 ) ;
assign n30195 =  ( n29922 ) ? ( VREG_8_8 ) : ( n30194 ) ;
assign n30196 =  ( n29921 ) ? ( VREG_8_9 ) : ( n30195 ) ;
assign n30197 =  ( n29920 ) ? ( VREG_8_10 ) : ( n30196 ) ;
assign n30198 =  ( n29919 ) ? ( VREG_8_11 ) : ( n30197 ) ;
assign n30199 =  ( n29918 ) ? ( VREG_8_12 ) : ( n30198 ) ;
assign n30200 =  ( n29917 ) ? ( VREG_8_13 ) : ( n30199 ) ;
assign n30201 =  ( n29916 ) ? ( VREG_8_14 ) : ( n30200 ) ;
assign n30202 =  ( n29915 ) ? ( VREG_8_15 ) : ( n30201 ) ;
assign n30203 =  ( n29914 ) ? ( VREG_9_0 ) : ( n30202 ) ;
assign n30204 =  ( n29913 ) ? ( VREG_9_1 ) : ( n30203 ) ;
assign n30205 =  ( n29912 ) ? ( VREG_9_2 ) : ( n30204 ) ;
assign n30206 =  ( n29911 ) ? ( VREG_9_3 ) : ( n30205 ) ;
assign n30207 =  ( n29910 ) ? ( VREG_9_4 ) : ( n30206 ) ;
assign n30208 =  ( n29909 ) ? ( VREG_9_5 ) : ( n30207 ) ;
assign n30209 =  ( n29908 ) ? ( VREG_9_6 ) : ( n30208 ) ;
assign n30210 =  ( n29907 ) ? ( VREG_9_7 ) : ( n30209 ) ;
assign n30211 =  ( n29906 ) ? ( VREG_9_8 ) : ( n30210 ) ;
assign n30212 =  ( n29905 ) ? ( VREG_9_9 ) : ( n30211 ) ;
assign n30213 =  ( n29904 ) ? ( VREG_9_10 ) : ( n30212 ) ;
assign n30214 =  ( n29903 ) ? ( VREG_9_11 ) : ( n30213 ) ;
assign n30215 =  ( n29902 ) ? ( VREG_9_12 ) : ( n30214 ) ;
assign n30216 =  ( n29901 ) ? ( VREG_9_13 ) : ( n30215 ) ;
assign n30217 =  ( n29900 ) ? ( VREG_9_14 ) : ( n30216 ) ;
assign n30218 =  ( n29899 ) ? ( VREG_9_15 ) : ( n30217 ) ;
assign n30219 =  ( n29898 ) ? ( VREG_10_0 ) : ( n30218 ) ;
assign n30220 =  ( n29897 ) ? ( VREG_10_1 ) : ( n30219 ) ;
assign n30221 =  ( n29896 ) ? ( VREG_10_2 ) : ( n30220 ) ;
assign n30222 =  ( n29895 ) ? ( VREG_10_3 ) : ( n30221 ) ;
assign n30223 =  ( n29894 ) ? ( VREG_10_4 ) : ( n30222 ) ;
assign n30224 =  ( n29893 ) ? ( VREG_10_5 ) : ( n30223 ) ;
assign n30225 =  ( n29892 ) ? ( VREG_10_6 ) : ( n30224 ) ;
assign n30226 =  ( n29891 ) ? ( VREG_10_7 ) : ( n30225 ) ;
assign n30227 =  ( n29890 ) ? ( VREG_10_8 ) : ( n30226 ) ;
assign n30228 =  ( n29889 ) ? ( VREG_10_9 ) : ( n30227 ) ;
assign n30229 =  ( n29888 ) ? ( VREG_10_10 ) : ( n30228 ) ;
assign n30230 =  ( n29887 ) ? ( VREG_10_11 ) : ( n30229 ) ;
assign n30231 =  ( n29886 ) ? ( VREG_10_12 ) : ( n30230 ) ;
assign n30232 =  ( n29885 ) ? ( VREG_10_13 ) : ( n30231 ) ;
assign n30233 =  ( n29884 ) ? ( VREG_10_14 ) : ( n30232 ) ;
assign n30234 =  ( n29883 ) ? ( VREG_10_15 ) : ( n30233 ) ;
assign n30235 =  ( n29882 ) ? ( VREG_11_0 ) : ( n30234 ) ;
assign n30236 =  ( n29881 ) ? ( VREG_11_1 ) : ( n30235 ) ;
assign n30237 =  ( n29880 ) ? ( VREG_11_2 ) : ( n30236 ) ;
assign n30238 =  ( n29879 ) ? ( VREG_11_3 ) : ( n30237 ) ;
assign n30239 =  ( n29878 ) ? ( VREG_11_4 ) : ( n30238 ) ;
assign n30240 =  ( n29877 ) ? ( VREG_11_5 ) : ( n30239 ) ;
assign n30241 =  ( n29876 ) ? ( VREG_11_6 ) : ( n30240 ) ;
assign n30242 =  ( n29875 ) ? ( VREG_11_7 ) : ( n30241 ) ;
assign n30243 =  ( n29874 ) ? ( VREG_11_8 ) : ( n30242 ) ;
assign n30244 =  ( n29873 ) ? ( VREG_11_9 ) : ( n30243 ) ;
assign n30245 =  ( n29872 ) ? ( VREG_11_10 ) : ( n30244 ) ;
assign n30246 =  ( n29871 ) ? ( VREG_11_11 ) : ( n30245 ) ;
assign n30247 =  ( n29870 ) ? ( VREG_11_12 ) : ( n30246 ) ;
assign n30248 =  ( n29869 ) ? ( VREG_11_13 ) : ( n30247 ) ;
assign n30249 =  ( n29868 ) ? ( VREG_11_14 ) : ( n30248 ) ;
assign n30250 =  ( n29867 ) ? ( VREG_11_15 ) : ( n30249 ) ;
assign n30251 =  ( n29866 ) ? ( VREG_12_0 ) : ( n30250 ) ;
assign n30252 =  ( n29865 ) ? ( VREG_12_1 ) : ( n30251 ) ;
assign n30253 =  ( n29864 ) ? ( VREG_12_2 ) : ( n30252 ) ;
assign n30254 =  ( n29863 ) ? ( VREG_12_3 ) : ( n30253 ) ;
assign n30255 =  ( n29862 ) ? ( VREG_12_4 ) : ( n30254 ) ;
assign n30256 =  ( n29861 ) ? ( VREG_12_5 ) : ( n30255 ) ;
assign n30257 =  ( n29860 ) ? ( VREG_12_6 ) : ( n30256 ) ;
assign n30258 =  ( n29859 ) ? ( VREG_12_7 ) : ( n30257 ) ;
assign n30259 =  ( n29858 ) ? ( VREG_12_8 ) : ( n30258 ) ;
assign n30260 =  ( n29857 ) ? ( VREG_12_9 ) : ( n30259 ) ;
assign n30261 =  ( n29856 ) ? ( VREG_12_10 ) : ( n30260 ) ;
assign n30262 =  ( n29855 ) ? ( VREG_12_11 ) : ( n30261 ) ;
assign n30263 =  ( n29854 ) ? ( VREG_12_12 ) : ( n30262 ) ;
assign n30264 =  ( n29853 ) ? ( VREG_12_13 ) : ( n30263 ) ;
assign n30265 =  ( n29852 ) ? ( VREG_12_14 ) : ( n30264 ) ;
assign n30266 =  ( n29851 ) ? ( VREG_12_15 ) : ( n30265 ) ;
assign n30267 =  ( n29850 ) ? ( VREG_13_0 ) : ( n30266 ) ;
assign n30268 =  ( n29849 ) ? ( VREG_13_1 ) : ( n30267 ) ;
assign n30269 =  ( n29848 ) ? ( VREG_13_2 ) : ( n30268 ) ;
assign n30270 =  ( n29847 ) ? ( VREG_13_3 ) : ( n30269 ) ;
assign n30271 =  ( n29846 ) ? ( VREG_13_4 ) : ( n30270 ) ;
assign n30272 =  ( n29845 ) ? ( VREG_13_5 ) : ( n30271 ) ;
assign n30273 =  ( n29844 ) ? ( VREG_13_6 ) : ( n30272 ) ;
assign n30274 =  ( n29843 ) ? ( VREG_13_7 ) : ( n30273 ) ;
assign n30275 =  ( n29842 ) ? ( VREG_13_8 ) : ( n30274 ) ;
assign n30276 =  ( n29841 ) ? ( VREG_13_9 ) : ( n30275 ) ;
assign n30277 =  ( n29840 ) ? ( VREG_13_10 ) : ( n30276 ) ;
assign n30278 =  ( n29839 ) ? ( VREG_13_11 ) : ( n30277 ) ;
assign n30279 =  ( n29838 ) ? ( VREG_13_12 ) : ( n30278 ) ;
assign n30280 =  ( n29837 ) ? ( VREG_13_13 ) : ( n30279 ) ;
assign n30281 =  ( n29836 ) ? ( VREG_13_14 ) : ( n30280 ) ;
assign n30282 =  ( n29835 ) ? ( VREG_13_15 ) : ( n30281 ) ;
assign n30283 =  ( n29834 ) ? ( VREG_14_0 ) : ( n30282 ) ;
assign n30284 =  ( n29833 ) ? ( VREG_14_1 ) : ( n30283 ) ;
assign n30285 =  ( n29832 ) ? ( VREG_14_2 ) : ( n30284 ) ;
assign n30286 =  ( n29831 ) ? ( VREG_14_3 ) : ( n30285 ) ;
assign n30287 =  ( n29830 ) ? ( VREG_14_4 ) : ( n30286 ) ;
assign n30288 =  ( n29829 ) ? ( VREG_14_5 ) : ( n30287 ) ;
assign n30289 =  ( n29828 ) ? ( VREG_14_6 ) : ( n30288 ) ;
assign n30290 =  ( n29827 ) ? ( VREG_14_7 ) : ( n30289 ) ;
assign n30291 =  ( n29826 ) ? ( VREG_14_8 ) : ( n30290 ) ;
assign n30292 =  ( n29825 ) ? ( VREG_14_9 ) : ( n30291 ) ;
assign n30293 =  ( n29824 ) ? ( VREG_14_10 ) : ( n30292 ) ;
assign n30294 =  ( n29823 ) ? ( VREG_14_11 ) : ( n30293 ) ;
assign n30295 =  ( n29822 ) ? ( VREG_14_12 ) : ( n30294 ) ;
assign n30296 =  ( n29821 ) ? ( VREG_14_13 ) : ( n30295 ) ;
assign n30297 =  ( n29820 ) ? ( VREG_14_14 ) : ( n30296 ) ;
assign n30298 =  ( n29819 ) ? ( VREG_14_15 ) : ( n30297 ) ;
assign n30299 =  ( n29818 ) ? ( VREG_15_0 ) : ( n30298 ) ;
assign n30300 =  ( n29817 ) ? ( VREG_15_1 ) : ( n30299 ) ;
assign n30301 =  ( n29816 ) ? ( VREG_15_2 ) : ( n30300 ) ;
assign n30302 =  ( n29815 ) ? ( VREG_15_3 ) : ( n30301 ) ;
assign n30303 =  ( n29814 ) ? ( VREG_15_4 ) : ( n30302 ) ;
assign n30304 =  ( n29813 ) ? ( VREG_15_5 ) : ( n30303 ) ;
assign n30305 =  ( n29812 ) ? ( VREG_15_6 ) : ( n30304 ) ;
assign n30306 =  ( n29811 ) ? ( VREG_15_7 ) : ( n30305 ) ;
assign n30307 =  ( n29810 ) ? ( VREG_15_8 ) : ( n30306 ) ;
assign n30308 =  ( n29809 ) ? ( VREG_15_9 ) : ( n30307 ) ;
assign n30309 =  ( n29808 ) ? ( VREG_15_10 ) : ( n30308 ) ;
assign n30310 =  ( n29807 ) ? ( VREG_15_11 ) : ( n30309 ) ;
assign n30311 =  ( n29806 ) ? ( VREG_15_12 ) : ( n30310 ) ;
assign n30312 =  ( n29805 ) ? ( VREG_15_13 ) : ( n30311 ) ;
assign n30313 =  ( n29804 ) ? ( VREG_15_14 ) : ( n30312 ) ;
assign n30314 =  ( n29803 ) ? ( VREG_15_15 ) : ( n30313 ) ;
assign n30315 =  ( n29802 ) ? ( VREG_16_0 ) : ( n30314 ) ;
assign n30316 =  ( n29801 ) ? ( VREG_16_1 ) : ( n30315 ) ;
assign n30317 =  ( n29800 ) ? ( VREG_16_2 ) : ( n30316 ) ;
assign n30318 =  ( n29799 ) ? ( VREG_16_3 ) : ( n30317 ) ;
assign n30319 =  ( n29798 ) ? ( VREG_16_4 ) : ( n30318 ) ;
assign n30320 =  ( n29797 ) ? ( VREG_16_5 ) : ( n30319 ) ;
assign n30321 =  ( n29796 ) ? ( VREG_16_6 ) : ( n30320 ) ;
assign n30322 =  ( n29795 ) ? ( VREG_16_7 ) : ( n30321 ) ;
assign n30323 =  ( n29794 ) ? ( VREG_16_8 ) : ( n30322 ) ;
assign n30324 =  ( n29793 ) ? ( VREG_16_9 ) : ( n30323 ) ;
assign n30325 =  ( n29792 ) ? ( VREG_16_10 ) : ( n30324 ) ;
assign n30326 =  ( n29791 ) ? ( VREG_16_11 ) : ( n30325 ) ;
assign n30327 =  ( n29790 ) ? ( VREG_16_12 ) : ( n30326 ) ;
assign n30328 =  ( n29789 ) ? ( VREG_16_13 ) : ( n30327 ) ;
assign n30329 =  ( n29788 ) ? ( VREG_16_14 ) : ( n30328 ) ;
assign n30330 =  ( n29787 ) ? ( VREG_16_15 ) : ( n30329 ) ;
assign n30331 =  ( n29786 ) ? ( VREG_17_0 ) : ( n30330 ) ;
assign n30332 =  ( n29785 ) ? ( VREG_17_1 ) : ( n30331 ) ;
assign n30333 =  ( n29784 ) ? ( VREG_17_2 ) : ( n30332 ) ;
assign n30334 =  ( n29783 ) ? ( VREG_17_3 ) : ( n30333 ) ;
assign n30335 =  ( n29782 ) ? ( VREG_17_4 ) : ( n30334 ) ;
assign n30336 =  ( n29781 ) ? ( VREG_17_5 ) : ( n30335 ) ;
assign n30337 =  ( n29780 ) ? ( VREG_17_6 ) : ( n30336 ) ;
assign n30338 =  ( n29779 ) ? ( VREG_17_7 ) : ( n30337 ) ;
assign n30339 =  ( n29778 ) ? ( VREG_17_8 ) : ( n30338 ) ;
assign n30340 =  ( n29777 ) ? ( VREG_17_9 ) : ( n30339 ) ;
assign n30341 =  ( n29776 ) ? ( VREG_17_10 ) : ( n30340 ) ;
assign n30342 =  ( n29775 ) ? ( VREG_17_11 ) : ( n30341 ) ;
assign n30343 =  ( n29774 ) ? ( VREG_17_12 ) : ( n30342 ) ;
assign n30344 =  ( n29773 ) ? ( VREG_17_13 ) : ( n30343 ) ;
assign n30345 =  ( n29772 ) ? ( VREG_17_14 ) : ( n30344 ) ;
assign n30346 =  ( n29771 ) ? ( VREG_17_15 ) : ( n30345 ) ;
assign n30347 =  ( n29770 ) ? ( VREG_18_0 ) : ( n30346 ) ;
assign n30348 =  ( n29769 ) ? ( VREG_18_1 ) : ( n30347 ) ;
assign n30349 =  ( n29768 ) ? ( VREG_18_2 ) : ( n30348 ) ;
assign n30350 =  ( n29767 ) ? ( VREG_18_3 ) : ( n30349 ) ;
assign n30351 =  ( n29766 ) ? ( VREG_18_4 ) : ( n30350 ) ;
assign n30352 =  ( n29765 ) ? ( VREG_18_5 ) : ( n30351 ) ;
assign n30353 =  ( n29764 ) ? ( VREG_18_6 ) : ( n30352 ) ;
assign n30354 =  ( n29763 ) ? ( VREG_18_7 ) : ( n30353 ) ;
assign n30355 =  ( n29762 ) ? ( VREG_18_8 ) : ( n30354 ) ;
assign n30356 =  ( n29761 ) ? ( VREG_18_9 ) : ( n30355 ) ;
assign n30357 =  ( n29760 ) ? ( VREG_18_10 ) : ( n30356 ) ;
assign n30358 =  ( n29759 ) ? ( VREG_18_11 ) : ( n30357 ) ;
assign n30359 =  ( n29758 ) ? ( VREG_18_12 ) : ( n30358 ) ;
assign n30360 =  ( n29757 ) ? ( VREG_18_13 ) : ( n30359 ) ;
assign n30361 =  ( n29756 ) ? ( VREG_18_14 ) : ( n30360 ) ;
assign n30362 =  ( n29755 ) ? ( VREG_18_15 ) : ( n30361 ) ;
assign n30363 =  ( n29754 ) ? ( VREG_19_0 ) : ( n30362 ) ;
assign n30364 =  ( n29753 ) ? ( VREG_19_1 ) : ( n30363 ) ;
assign n30365 =  ( n29752 ) ? ( VREG_19_2 ) : ( n30364 ) ;
assign n30366 =  ( n29751 ) ? ( VREG_19_3 ) : ( n30365 ) ;
assign n30367 =  ( n29750 ) ? ( VREG_19_4 ) : ( n30366 ) ;
assign n30368 =  ( n29749 ) ? ( VREG_19_5 ) : ( n30367 ) ;
assign n30369 =  ( n29748 ) ? ( VREG_19_6 ) : ( n30368 ) ;
assign n30370 =  ( n29747 ) ? ( VREG_19_7 ) : ( n30369 ) ;
assign n30371 =  ( n29746 ) ? ( VREG_19_8 ) : ( n30370 ) ;
assign n30372 =  ( n29745 ) ? ( VREG_19_9 ) : ( n30371 ) ;
assign n30373 =  ( n29744 ) ? ( VREG_19_10 ) : ( n30372 ) ;
assign n30374 =  ( n29743 ) ? ( VREG_19_11 ) : ( n30373 ) ;
assign n30375 =  ( n29742 ) ? ( VREG_19_12 ) : ( n30374 ) ;
assign n30376 =  ( n29741 ) ? ( VREG_19_13 ) : ( n30375 ) ;
assign n30377 =  ( n29740 ) ? ( VREG_19_14 ) : ( n30376 ) ;
assign n30378 =  ( n29739 ) ? ( VREG_19_15 ) : ( n30377 ) ;
assign n30379 =  ( n29738 ) ? ( VREG_20_0 ) : ( n30378 ) ;
assign n30380 =  ( n29737 ) ? ( VREG_20_1 ) : ( n30379 ) ;
assign n30381 =  ( n29736 ) ? ( VREG_20_2 ) : ( n30380 ) ;
assign n30382 =  ( n29735 ) ? ( VREG_20_3 ) : ( n30381 ) ;
assign n30383 =  ( n29734 ) ? ( VREG_20_4 ) : ( n30382 ) ;
assign n30384 =  ( n29733 ) ? ( VREG_20_5 ) : ( n30383 ) ;
assign n30385 =  ( n29732 ) ? ( VREG_20_6 ) : ( n30384 ) ;
assign n30386 =  ( n29731 ) ? ( VREG_20_7 ) : ( n30385 ) ;
assign n30387 =  ( n29730 ) ? ( VREG_20_8 ) : ( n30386 ) ;
assign n30388 =  ( n29729 ) ? ( VREG_20_9 ) : ( n30387 ) ;
assign n30389 =  ( n29728 ) ? ( VREG_20_10 ) : ( n30388 ) ;
assign n30390 =  ( n29727 ) ? ( VREG_20_11 ) : ( n30389 ) ;
assign n30391 =  ( n29726 ) ? ( VREG_20_12 ) : ( n30390 ) ;
assign n30392 =  ( n29725 ) ? ( VREG_20_13 ) : ( n30391 ) ;
assign n30393 =  ( n29724 ) ? ( VREG_20_14 ) : ( n30392 ) ;
assign n30394 =  ( n29723 ) ? ( VREG_20_15 ) : ( n30393 ) ;
assign n30395 =  ( n29722 ) ? ( VREG_21_0 ) : ( n30394 ) ;
assign n30396 =  ( n29721 ) ? ( VREG_21_1 ) : ( n30395 ) ;
assign n30397 =  ( n29720 ) ? ( VREG_21_2 ) : ( n30396 ) ;
assign n30398 =  ( n29719 ) ? ( VREG_21_3 ) : ( n30397 ) ;
assign n30399 =  ( n29718 ) ? ( VREG_21_4 ) : ( n30398 ) ;
assign n30400 =  ( n29717 ) ? ( VREG_21_5 ) : ( n30399 ) ;
assign n30401 =  ( n29716 ) ? ( VREG_21_6 ) : ( n30400 ) ;
assign n30402 =  ( n29715 ) ? ( VREG_21_7 ) : ( n30401 ) ;
assign n30403 =  ( n29714 ) ? ( VREG_21_8 ) : ( n30402 ) ;
assign n30404 =  ( n29713 ) ? ( VREG_21_9 ) : ( n30403 ) ;
assign n30405 =  ( n29712 ) ? ( VREG_21_10 ) : ( n30404 ) ;
assign n30406 =  ( n29711 ) ? ( VREG_21_11 ) : ( n30405 ) ;
assign n30407 =  ( n29710 ) ? ( VREG_21_12 ) : ( n30406 ) ;
assign n30408 =  ( n29709 ) ? ( VREG_21_13 ) : ( n30407 ) ;
assign n30409 =  ( n29708 ) ? ( VREG_21_14 ) : ( n30408 ) ;
assign n30410 =  ( n29707 ) ? ( VREG_21_15 ) : ( n30409 ) ;
assign n30411 =  ( n29706 ) ? ( VREG_22_0 ) : ( n30410 ) ;
assign n30412 =  ( n29705 ) ? ( VREG_22_1 ) : ( n30411 ) ;
assign n30413 =  ( n29704 ) ? ( VREG_22_2 ) : ( n30412 ) ;
assign n30414 =  ( n29703 ) ? ( VREG_22_3 ) : ( n30413 ) ;
assign n30415 =  ( n29702 ) ? ( VREG_22_4 ) : ( n30414 ) ;
assign n30416 =  ( n29701 ) ? ( VREG_22_5 ) : ( n30415 ) ;
assign n30417 =  ( n29700 ) ? ( VREG_22_6 ) : ( n30416 ) ;
assign n30418 =  ( n29699 ) ? ( VREG_22_7 ) : ( n30417 ) ;
assign n30419 =  ( n29698 ) ? ( VREG_22_8 ) : ( n30418 ) ;
assign n30420 =  ( n29697 ) ? ( VREG_22_9 ) : ( n30419 ) ;
assign n30421 =  ( n29696 ) ? ( VREG_22_10 ) : ( n30420 ) ;
assign n30422 =  ( n29695 ) ? ( VREG_22_11 ) : ( n30421 ) ;
assign n30423 =  ( n29694 ) ? ( VREG_22_12 ) : ( n30422 ) ;
assign n30424 =  ( n29693 ) ? ( VREG_22_13 ) : ( n30423 ) ;
assign n30425 =  ( n29692 ) ? ( VREG_22_14 ) : ( n30424 ) ;
assign n30426 =  ( n29691 ) ? ( VREG_22_15 ) : ( n30425 ) ;
assign n30427 =  ( n29690 ) ? ( VREG_23_0 ) : ( n30426 ) ;
assign n30428 =  ( n29689 ) ? ( VREG_23_1 ) : ( n30427 ) ;
assign n30429 =  ( n29688 ) ? ( VREG_23_2 ) : ( n30428 ) ;
assign n30430 =  ( n29687 ) ? ( VREG_23_3 ) : ( n30429 ) ;
assign n30431 =  ( n29686 ) ? ( VREG_23_4 ) : ( n30430 ) ;
assign n30432 =  ( n29685 ) ? ( VREG_23_5 ) : ( n30431 ) ;
assign n30433 =  ( n29684 ) ? ( VREG_23_6 ) : ( n30432 ) ;
assign n30434 =  ( n29683 ) ? ( VREG_23_7 ) : ( n30433 ) ;
assign n30435 =  ( n29682 ) ? ( VREG_23_8 ) : ( n30434 ) ;
assign n30436 =  ( n29681 ) ? ( VREG_23_9 ) : ( n30435 ) ;
assign n30437 =  ( n29680 ) ? ( VREG_23_10 ) : ( n30436 ) ;
assign n30438 =  ( n29679 ) ? ( VREG_23_11 ) : ( n30437 ) ;
assign n30439 =  ( n29678 ) ? ( VREG_23_12 ) : ( n30438 ) ;
assign n30440 =  ( n29677 ) ? ( VREG_23_13 ) : ( n30439 ) ;
assign n30441 =  ( n29676 ) ? ( VREG_23_14 ) : ( n30440 ) ;
assign n30442 =  ( n29675 ) ? ( VREG_23_15 ) : ( n30441 ) ;
assign n30443 =  ( n29674 ) ? ( VREG_24_0 ) : ( n30442 ) ;
assign n30444 =  ( n29673 ) ? ( VREG_24_1 ) : ( n30443 ) ;
assign n30445 =  ( n29672 ) ? ( VREG_24_2 ) : ( n30444 ) ;
assign n30446 =  ( n29671 ) ? ( VREG_24_3 ) : ( n30445 ) ;
assign n30447 =  ( n29670 ) ? ( VREG_24_4 ) : ( n30446 ) ;
assign n30448 =  ( n29669 ) ? ( VREG_24_5 ) : ( n30447 ) ;
assign n30449 =  ( n29668 ) ? ( VREG_24_6 ) : ( n30448 ) ;
assign n30450 =  ( n29667 ) ? ( VREG_24_7 ) : ( n30449 ) ;
assign n30451 =  ( n29666 ) ? ( VREG_24_8 ) : ( n30450 ) ;
assign n30452 =  ( n29665 ) ? ( VREG_24_9 ) : ( n30451 ) ;
assign n30453 =  ( n29664 ) ? ( VREG_24_10 ) : ( n30452 ) ;
assign n30454 =  ( n29663 ) ? ( VREG_24_11 ) : ( n30453 ) ;
assign n30455 =  ( n29662 ) ? ( VREG_24_12 ) : ( n30454 ) ;
assign n30456 =  ( n29661 ) ? ( VREG_24_13 ) : ( n30455 ) ;
assign n30457 =  ( n29660 ) ? ( VREG_24_14 ) : ( n30456 ) ;
assign n30458 =  ( n29659 ) ? ( VREG_24_15 ) : ( n30457 ) ;
assign n30459 =  ( n29658 ) ? ( VREG_25_0 ) : ( n30458 ) ;
assign n30460 =  ( n29657 ) ? ( VREG_25_1 ) : ( n30459 ) ;
assign n30461 =  ( n29656 ) ? ( VREG_25_2 ) : ( n30460 ) ;
assign n30462 =  ( n29655 ) ? ( VREG_25_3 ) : ( n30461 ) ;
assign n30463 =  ( n29654 ) ? ( VREG_25_4 ) : ( n30462 ) ;
assign n30464 =  ( n29653 ) ? ( VREG_25_5 ) : ( n30463 ) ;
assign n30465 =  ( n29652 ) ? ( VREG_25_6 ) : ( n30464 ) ;
assign n30466 =  ( n29651 ) ? ( VREG_25_7 ) : ( n30465 ) ;
assign n30467 =  ( n29650 ) ? ( VREG_25_8 ) : ( n30466 ) ;
assign n30468 =  ( n29649 ) ? ( VREG_25_9 ) : ( n30467 ) ;
assign n30469 =  ( n29648 ) ? ( VREG_25_10 ) : ( n30468 ) ;
assign n30470 =  ( n29647 ) ? ( VREG_25_11 ) : ( n30469 ) ;
assign n30471 =  ( n29646 ) ? ( VREG_25_12 ) : ( n30470 ) ;
assign n30472 =  ( n29645 ) ? ( VREG_25_13 ) : ( n30471 ) ;
assign n30473 =  ( n29644 ) ? ( VREG_25_14 ) : ( n30472 ) ;
assign n30474 =  ( n29643 ) ? ( VREG_25_15 ) : ( n30473 ) ;
assign n30475 =  ( n29642 ) ? ( VREG_26_0 ) : ( n30474 ) ;
assign n30476 =  ( n29641 ) ? ( VREG_26_1 ) : ( n30475 ) ;
assign n30477 =  ( n29640 ) ? ( VREG_26_2 ) : ( n30476 ) ;
assign n30478 =  ( n29639 ) ? ( VREG_26_3 ) : ( n30477 ) ;
assign n30479 =  ( n29638 ) ? ( VREG_26_4 ) : ( n30478 ) ;
assign n30480 =  ( n29637 ) ? ( VREG_26_5 ) : ( n30479 ) ;
assign n30481 =  ( n29636 ) ? ( VREG_26_6 ) : ( n30480 ) ;
assign n30482 =  ( n29635 ) ? ( VREG_26_7 ) : ( n30481 ) ;
assign n30483 =  ( n29634 ) ? ( VREG_26_8 ) : ( n30482 ) ;
assign n30484 =  ( n29633 ) ? ( VREG_26_9 ) : ( n30483 ) ;
assign n30485 =  ( n29632 ) ? ( VREG_26_10 ) : ( n30484 ) ;
assign n30486 =  ( n29631 ) ? ( VREG_26_11 ) : ( n30485 ) ;
assign n30487 =  ( n29630 ) ? ( VREG_26_12 ) : ( n30486 ) ;
assign n30488 =  ( n29629 ) ? ( VREG_26_13 ) : ( n30487 ) ;
assign n30489 =  ( n29628 ) ? ( VREG_26_14 ) : ( n30488 ) ;
assign n30490 =  ( n29627 ) ? ( VREG_26_15 ) : ( n30489 ) ;
assign n30491 =  ( n29626 ) ? ( VREG_27_0 ) : ( n30490 ) ;
assign n30492 =  ( n29625 ) ? ( VREG_27_1 ) : ( n30491 ) ;
assign n30493 =  ( n29624 ) ? ( VREG_27_2 ) : ( n30492 ) ;
assign n30494 =  ( n29623 ) ? ( VREG_27_3 ) : ( n30493 ) ;
assign n30495 =  ( n29622 ) ? ( VREG_27_4 ) : ( n30494 ) ;
assign n30496 =  ( n29621 ) ? ( VREG_27_5 ) : ( n30495 ) ;
assign n30497 =  ( n29620 ) ? ( VREG_27_6 ) : ( n30496 ) ;
assign n30498 =  ( n29619 ) ? ( VREG_27_7 ) : ( n30497 ) ;
assign n30499 =  ( n29618 ) ? ( VREG_27_8 ) : ( n30498 ) ;
assign n30500 =  ( n29617 ) ? ( VREG_27_9 ) : ( n30499 ) ;
assign n30501 =  ( n29616 ) ? ( VREG_27_10 ) : ( n30500 ) ;
assign n30502 =  ( n29615 ) ? ( VREG_27_11 ) : ( n30501 ) ;
assign n30503 =  ( n29614 ) ? ( VREG_27_12 ) : ( n30502 ) ;
assign n30504 =  ( n29613 ) ? ( VREG_27_13 ) : ( n30503 ) ;
assign n30505 =  ( n29612 ) ? ( VREG_27_14 ) : ( n30504 ) ;
assign n30506 =  ( n29611 ) ? ( VREG_27_15 ) : ( n30505 ) ;
assign n30507 =  ( n29610 ) ? ( VREG_28_0 ) : ( n30506 ) ;
assign n30508 =  ( n29609 ) ? ( VREG_28_1 ) : ( n30507 ) ;
assign n30509 =  ( n29608 ) ? ( VREG_28_2 ) : ( n30508 ) ;
assign n30510 =  ( n29607 ) ? ( VREG_28_3 ) : ( n30509 ) ;
assign n30511 =  ( n29606 ) ? ( VREG_28_4 ) : ( n30510 ) ;
assign n30512 =  ( n29605 ) ? ( VREG_28_5 ) : ( n30511 ) ;
assign n30513 =  ( n29604 ) ? ( VREG_28_6 ) : ( n30512 ) ;
assign n30514 =  ( n29603 ) ? ( VREG_28_7 ) : ( n30513 ) ;
assign n30515 =  ( n29602 ) ? ( VREG_28_8 ) : ( n30514 ) ;
assign n30516 =  ( n29601 ) ? ( VREG_28_9 ) : ( n30515 ) ;
assign n30517 =  ( n29600 ) ? ( VREG_28_10 ) : ( n30516 ) ;
assign n30518 =  ( n29599 ) ? ( VREG_28_11 ) : ( n30517 ) ;
assign n30519 =  ( n29598 ) ? ( VREG_28_12 ) : ( n30518 ) ;
assign n30520 =  ( n29597 ) ? ( VREG_28_13 ) : ( n30519 ) ;
assign n30521 =  ( n29596 ) ? ( VREG_28_14 ) : ( n30520 ) ;
assign n30522 =  ( n29595 ) ? ( VREG_28_15 ) : ( n30521 ) ;
assign n30523 =  ( n29594 ) ? ( VREG_29_0 ) : ( n30522 ) ;
assign n30524 =  ( n29593 ) ? ( VREG_29_1 ) : ( n30523 ) ;
assign n30525 =  ( n29592 ) ? ( VREG_29_2 ) : ( n30524 ) ;
assign n30526 =  ( n29591 ) ? ( VREG_29_3 ) : ( n30525 ) ;
assign n30527 =  ( n29590 ) ? ( VREG_29_4 ) : ( n30526 ) ;
assign n30528 =  ( n29589 ) ? ( VREG_29_5 ) : ( n30527 ) ;
assign n30529 =  ( n29588 ) ? ( VREG_29_6 ) : ( n30528 ) ;
assign n30530 =  ( n29587 ) ? ( VREG_29_7 ) : ( n30529 ) ;
assign n30531 =  ( n29586 ) ? ( VREG_29_8 ) : ( n30530 ) ;
assign n30532 =  ( n29585 ) ? ( VREG_29_9 ) : ( n30531 ) ;
assign n30533 =  ( n29584 ) ? ( VREG_29_10 ) : ( n30532 ) ;
assign n30534 =  ( n29583 ) ? ( VREG_29_11 ) : ( n30533 ) ;
assign n30535 =  ( n29582 ) ? ( VREG_29_12 ) : ( n30534 ) ;
assign n30536 =  ( n29581 ) ? ( VREG_29_13 ) : ( n30535 ) ;
assign n30537 =  ( n29580 ) ? ( VREG_29_14 ) : ( n30536 ) ;
assign n30538 =  ( n29579 ) ? ( VREG_29_15 ) : ( n30537 ) ;
assign n30539 =  ( n29578 ) ? ( VREG_30_0 ) : ( n30538 ) ;
assign n30540 =  ( n29577 ) ? ( VREG_30_1 ) : ( n30539 ) ;
assign n30541 =  ( n29576 ) ? ( VREG_30_2 ) : ( n30540 ) ;
assign n30542 =  ( n29575 ) ? ( VREG_30_3 ) : ( n30541 ) ;
assign n30543 =  ( n29574 ) ? ( VREG_30_4 ) : ( n30542 ) ;
assign n30544 =  ( n29573 ) ? ( VREG_30_5 ) : ( n30543 ) ;
assign n30545 =  ( n29572 ) ? ( VREG_30_6 ) : ( n30544 ) ;
assign n30546 =  ( n29571 ) ? ( VREG_30_7 ) : ( n30545 ) ;
assign n30547 =  ( n29570 ) ? ( VREG_30_8 ) : ( n30546 ) ;
assign n30548 =  ( n29569 ) ? ( VREG_30_9 ) : ( n30547 ) ;
assign n30549 =  ( n29568 ) ? ( VREG_30_10 ) : ( n30548 ) ;
assign n30550 =  ( n29567 ) ? ( VREG_30_11 ) : ( n30549 ) ;
assign n30551 =  ( n29566 ) ? ( VREG_30_12 ) : ( n30550 ) ;
assign n30552 =  ( n29565 ) ? ( VREG_30_13 ) : ( n30551 ) ;
assign n30553 =  ( n29564 ) ? ( VREG_30_14 ) : ( n30552 ) ;
assign n30554 =  ( n29563 ) ? ( VREG_30_15 ) : ( n30553 ) ;
assign n30555 =  ( n29562 ) ? ( VREG_31_0 ) : ( n30554 ) ;
assign n30556 =  ( n29561 ) ? ( VREG_31_1 ) : ( n30555 ) ;
assign n30557 =  ( n29560 ) ? ( VREG_31_2 ) : ( n30556 ) ;
assign n30558 =  ( n29559 ) ? ( VREG_31_3 ) : ( n30557 ) ;
assign n30559 =  ( n29558 ) ? ( VREG_31_4 ) : ( n30558 ) ;
assign n30560 =  ( n29557 ) ? ( VREG_31_5 ) : ( n30559 ) ;
assign n30561 =  ( n29556 ) ? ( VREG_31_6 ) : ( n30560 ) ;
assign n30562 =  ( n29555 ) ? ( VREG_31_7 ) : ( n30561 ) ;
assign n30563 =  ( n29554 ) ? ( VREG_31_8 ) : ( n30562 ) ;
assign n30564 =  ( n29553 ) ? ( VREG_31_9 ) : ( n30563 ) ;
assign n30565 =  ( n29552 ) ? ( VREG_31_10 ) : ( n30564 ) ;
assign n30566 =  ( n29551 ) ? ( VREG_31_11 ) : ( n30565 ) ;
assign n30567 =  ( n29550 ) ? ( VREG_31_12 ) : ( n30566 ) ;
assign n30568 =  ( n29549 ) ? ( VREG_31_13 ) : ( n30567 ) ;
assign n30569 =  ( n29548 ) ? ( VREG_31_14 ) : ( n30568 ) ;
assign n30570 =  ( n29547 ) ? ( VREG_31_15 ) : ( n30569 ) ;
assign n30571 =  ( n29536 ) + ( n30570 )  ;
assign n30572 =  ( n29536 ) - ( n30570 )  ;
assign n30573 =  ( n29536 ) & ( n30570 )  ;
assign n30574 =  ( n29536 ) | ( n30570 )  ;
assign n30575 =  ( ( n29536 ) * ( n30570 ))  ;
assign n30576 =  ( n148 ) ? ( n30575 ) : ( VREG_0_7 ) ;
assign n30577 =  ( n146 ) ? ( n30574 ) : ( n30576 ) ;
assign n30578 =  ( n144 ) ? ( n30573 ) : ( n30577 ) ;
assign n30579 =  ( n142 ) ? ( n30572 ) : ( n30578 ) ;
assign n30580 =  ( n10 ) ? ( n30571 ) : ( n30579 ) ;
assign n30581 = n3030[7:7] ;
assign n30582 =  ( n30581 ) == ( 1'd0 )  ;
assign n30583 =  ( n30582 ) ? ( VREG_0_7 ) : ( n29546 ) ;
assign n30584 =  ( n30582 ) ? ( VREG_0_7 ) : ( n30580 ) ;
assign n30585 =  ( n3034 ) ? ( n30584 ) : ( VREG_0_7 ) ;
assign n30586 =  ( n2965 ) ? ( n30583 ) : ( n30585 ) ;
assign n30587 =  ( n1930 ) ? ( n30580 ) : ( n30586 ) ;
assign n30588 =  ( n879 ) ? ( n29546 ) : ( n30587 ) ;
assign n30589 =  ( n29536 ) + ( n164 )  ;
assign n30590 =  ( n29536 ) - ( n164 )  ;
assign n30591 =  ( n29536 ) & ( n164 )  ;
assign n30592 =  ( n29536 ) | ( n164 )  ;
assign n30593 =  ( ( n29536 ) * ( n164 ))  ;
assign n30594 =  ( n172 ) ? ( n30593 ) : ( VREG_0_7 ) ;
assign n30595 =  ( n170 ) ? ( n30592 ) : ( n30594 ) ;
assign n30596 =  ( n168 ) ? ( n30591 ) : ( n30595 ) ;
assign n30597 =  ( n166 ) ? ( n30590 ) : ( n30596 ) ;
assign n30598 =  ( n162 ) ? ( n30589 ) : ( n30597 ) ;
assign n30599 =  ( n29536 ) + ( n180 )  ;
assign n30600 =  ( n29536 ) - ( n180 )  ;
assign n30601 =  ( n29536 ) & ( n180 )  ;
assign n30602 =  ( n29536 ) | ( n180 )  ;
assign n30603 =  ( ( n29536 ) * ( n180 ))  ;
assign n30604 =  ( n172 ) ? ( n30603 ) : ( VREG_0_7 ) ;
assign n30605 =  ( n170 ) ? ( n30602 ) : ( n30604 ) ;
assign n30606 =  ( n168 ) ? ( n30601 ) : ( n30605 ) ;
assign n30607 =  ( n166 ) ? ( n30600 ) : ( n30606 ) ;
assign n30608 =  ( n162 ) ? ( n30599 ) : ( n30607 ) ;
assign n30609 =  ( n30582 ) ? ( VREG_0_7 ) : ( n30608 ) ;
assign n30610 =  ( n3051 ) ? ( n30609 ) : ( VREG_0_7 ) ;
assign n30611 =  ( n3040 ) ? ( n30598 ) : ( n30610 ) ;
assign n30612 =  ( n192 ) ? ( VREG_0_7 ) : ( VREG_0_7 ) ;
assign n30613 =  ( n157 ) ? ( n30611 ) : ( n30612 ) ;
assign n30614 =  ( n6 ) ? ( n30588 ) : ( n30613 ) ;
assign n30615 =  ( n4 ) ? ( n30614 ) : ( VREG_0_7 ) ;
assign n30616 =  ( 32'd8 ) == ( 32'd15 )  ;
assign n30617 =  ( n12 ) & ( n30616 )  ;
assign n30618 =  ( 32'd8 ) == ( 32'd14 )  ;
assign n30619 =  ( n12 ) & ( n30618 )  ;
assign n30620 =  ( 32'd8 ) == ( 32'd13 )  ;
assign n30621 =  ( n12 ) & ( n30620 )  ;
assign n30622 =  ( 32'd8 ) == ( 32'd12 )  ;
assign n30623 =  ( n12 ) & ( n30622 )  ;
assign n30624 =  ( 32'd8 ) == ( 32'd11 )  ;
assign n30625 =  ( n12 ) & ( n30624 )  ;
assign n30626 =  ( 32'd8 ) == ( 32'd10 )  ;
assign n30627 =  ( n12 ) & ( n30626 )  ;
assign n30628 =  ( 32'd8 ) == ( 32'd9 )  ;
assign n30629 =  ( n12 ) & ( n30628 )  ;
assign n30630 =  ( 32'd8 ) == ( 32'd8 )  ;
assign n30631 =  ( n12 ) & ( n30630 )  ;
assign n30632 =  ( 32'd8 ) == ( 32'd7 )  ;
assign n30633 =  ( n12 ) & ( n30632 )  ;
assign n30634 =  ( 32'd8 ) == ( 32'd6 )  ;
assign n30635 =  ( n12 ) & ( n30634 )  ;
assign n30636 =  ( 32'd8 ) == ( 32'd5 )  ;
assign n30637 =  ( n12 ) & ( n30636 )  ;
assign n30638 =  ( 32'd8 ) == ( 32'd4 )  ;
assign n30639 =  ( n12 ) & ( n30638 )  ;
assign n30640 =  ( 32'd8 ) == ( 32'd3 )  ;
assign n30641 =  ( n12 ) & ( n30640 )  ;
assign n30642 =  ( 32'd8 ) == ( 32'd2 )  ;
assign n30643 =  ( n12 ) & ( n30642 )  ;
assign n30644 =  ( 32'd8 ) == ( 32'd1 )  ;
assign n30645 =  ( n12 ) & ( n30644 )  ;
assign n30646 =  ( 32'd8 ) == ( 32'd0 )  ;
assign n30647 =  ( n12 ) & ( n30646 )  ;
assign n30648 =  ( n13 ) & ( n30616 )  ;
assign n30649 =  ( n13 ) & ( n30618 )  ;
assign n30650 =  ( n13 ) & ( n30620 )  ;
assign n30651 =  ( n13 ) & ( n30622 )  ;
assign n30652 =  ( n13 ) & ( n30624 )  ;
assign n30653 =  ( n13 ) & ( n30626 )  ;
assign n30654 =  ( n13 ) & ( n30628 )  ;
assign n30655 =  ( n13 ) & ( n30630 )  ;
assign n30656 =  ( n13 ) & ( n30632 )  ;
assign n30657 =  ( n13 ) & ( n30634 )  ;
assign n30658 =  ( n13 ) & ( n30636 )  ;
assign n30659 =  ( n13 ) & ( n30638 )  ;
assign n30660 =  ( n13 ) & ( n30640 )  ;
assign n30661 =  ( n13 ) & ( n30642 )  ;
assign n30662 =  ( n13 ) & ( n30644 )  ;
assign n30663 =  ( n13 ) & ( n30646 )  ;
assign n30664 =  ( n14 ) & ( n30616 )  ;
assign n30665 =  ( n14 ) & ( n30618 )  ;
assign n30666 =  ( n14 ) & ( n30620 )  ;
assign n30667 =  ( n14 ) & ( n30622 )  ;
assign n30668 =  ( n14 ) & ( n30624 )  ;
assign n30669 =  ( n14 ) & ( n30626 )  ;
assign n30670 =  ( n14 ) & ( n30628 )  ;
assign n30671 =  ( n14 ) & ( n30630 )  ;
assign n30672 =  ( n14 ) & ( n30632 )  ;
assign n30673 =  ( n14 ) & ( n30634 )  ;
assign n30674 =  ( n14 ) & ( n30636 )  ;
assign n30675 =  ( n14 ) & ( n30638 )  ;
assign n30676 =  ( n14 ) & ( n30640 )  ;
assign n30677 =  ( n14 ) & ( n30642 )  ;
assign n30678 =  ( n14 ) & ( n30644 )  ;
assign n30679 =  ( n14 ) & ( n30646 )  ;
assign n30680 =  ( n15 ) & ( n30616 )  ;
assign n30681 =  ( n15 ) & ( n30618 )  ;
assign n30682 =  ( n15 ) & ( n30620 )  ;
assign n30683 =  ( n15 ) & ( n30622 )  ;
assign n30684 =  ( n15 ) & ( n30624 )  ;
assign n30685 =  ( n15 ) & ( n30626 )  ;
assign n30686 =  ( n15 ) & ( n30628 )  ;
assign n30687 =  ( n15 ) & ( n30630 )  ;
assign n30688 =  ( n15 ) & ( n30632 )  ;
assign n30689 =  ( n15 ) & ( n30634 )  ;
assign n30690 =  ( n15 ) & ( n30636 )  ;
assign n30691 =  ( n15 ) & ( n30638 )  ;
assign n30692 =  ( n15 ) & ( n30640 )  ;
assign n30693 =  ( n15 ) & ( n30642 )  ;
assign n30694 =  ( n15 ) & ( n30644 )  ;
assign n30695 =  ( n15 ) & ( n30646 )  ;
assign n30696 =  ( n16 ) & ( n30616 )  ;
assign n30697 =  ( n16 ) & ( n30618 )  ;
assign n30698 =  ( n16 ) & ( n30620 )  ;
assign n30699 =  ( n16 ) & ( n30622 )  ;
assign n30700 =  ( n16 ) & ( n30624 )  ;
assign n30701 =  ( n16 ) & ( n30626 )  ;
assign n30702 =  ( n16 ) & ( n30628 )  ;
assign n30703 =  ( n16 ) & ( n30630 )  ;
assign n30704 =  ( n16 ) & ( n30632 )  ;
assign n30705 =  ( n16 ) & ( n30634 )  ;
assign n30706 =  ( n16 ) & ( n30636 )  ;
assign n30707 =  ( n16 ) & ( n30638 )  ;
assign n30708 =  ( n16 ) & ( n30640 )  ;
assign n30709 =  ( n16 ) & ( n30642 )  ;
assign n30710 =  ( n16 ) & ( n30644 )  ;
assign n30711 =  ( n16 ) & ( n30646 )  ;
assign n30712 =  ( n17 ) & ( n30616 )  ;
assign n30713 =  ( n17 ) & ( n30618 )  ;
assign n30714 =  ( n17 ) & ( n30620 )  ;
assign n30715 =  ( n17 ) & ( n30622 )  ;
assign n30716 =  ( n17 ) & ( n30624 )  ;
assign n30717 =  ( n17 ) & ( n30626 )  ;
assign n30718 =  ( n17 ) & ( n30628 )  ;
assign n30719 =  ( n17 ) & ( n30630 )  ;
assign n30720 =  ( n17 ) & ( n30632 )  ;
assign n30721 =  ( n17 ) & ( n30634 )  ;
assign n30722 =  ( n17 ) & ( n30636 )  ;
assign n30723 =  ( n17 ) & ( n30638 )  ;
assign n30724 =  ( n17 ) & ( n30640 )  ;
assign n30725 =  ( n17 ) & ( n30642 )  ;
assign n30726 =  ( n17 ) & ( n30644 )  ;
assign n30727 =  ( n17 ) & ( n30646 )  ;
assign n30728 =  ( n18 ) & ( n30616 )  ;
assign n30729 =  ( n18 ) & ( n30618 )  ;
assign n30730 =  ( n18 ) & ( n30620 )  ;
assign n30731 =  ( n18 ) & ( n30622 )  ;
assign n30732 =  ( n18 ) & ( n30624 )  ;
assign n30733 =  ( n18 ) & ( n30626 )  ;
assign n30734 =  ( n18 ) & ( n30628 )  ;
assign n30735 =  ( n18 ) & ( n30630 )  ;
assign n30736 =  ( n18 ) & ( n30632 )  ;
assign n30737 =  ( n18 ) & ( n30634 )  ;
assign n30738 =  ( n18 ) & ( n30636 )  ;
assign n30739 =  ( n18 ) & ( n30638 )  ;
assign n30740 =  ( n18 ) & ( n30640 )  ;
assign n30741 =  ( n18 ) & ( n30642 )  ;
assign n30742 =  ( n18 ) & ( n30644 )  ;
assign n30743 =  ( n18 ) & ( n30646 )  ;
assign n30744 =  ( n19 ) & ( n30616 )  ;
assign n30745 =  ( n19 ) & ( n30618 )  ;
assign n30746 =  ( n19 ) & ( n30620 )  ;
assign n30747 =  ( n19 ) & ( n30622 )  ;
assign n30748 =  ( n19 ) & ( n30624 )  ;
assign n30749 =  ( n19 ) & ( n30626 )  ;
assign n30750 =  ( n19 ) & ( n30628 )  ;
assign n30751 =  ( n19 ) & ( n30630 )  ;
assign n30752 =  ( n19 ) & ( n30632 )  ;
assign n30753 =  ( n19 ) & ( n30634 )  ;
assign n30754 =  ( n19 ) & ( n30636 )  ;
assign n30755 =  ( n19 ) & ( n30638 )  ;
assign n30756 =  ( n19 ) & ( n30640 )  ;
assign n30757 =  ( n19 ) & ( n30642 )  ;
assign n30758 =  ( n19 ) & ( n30644 )  ;
assign n30759 =  ( n19 ) & ( n30646 )  ;
assign n30760 =  ( n20 ) & ( n30616 )  ;
assign n30761 =  ( n20 ) & ( n30618 )  ;
assign n30762 =  ( n20 ) & ( n30620 )  ;
assign n30763 =  ( n20 ) & ( n30622 )  ;
assign n30764 =  ( n20 ) & ( n30624 )  ;
assign n30765 =  ( n20 ) & ( n30626 )  ;
assign n30766 =  ( n20 ) & ( n30628 )  ;
assign n30767 =  ( n20 ) & ( n30630 )  ;
assign n30768 =  ( n20 ) & ( n30632 )  ;
assign n30769 =  ( n20 ) & ( n30634 )  ;
assign n30770 =  ( n20 ) & ( n30636 )  ;
assign n30771 =  ( n20 ) & ( n30638 )  ;
assign n30772 =  ( n20 ) & ( n30640 )  ;
assign n30773 =  ( n20 ) & ( n30642 )  ;
assign n30774 =  ( n20 ) & ( n30644 )  ;
assign n30775 =  ( n20 ) & ( n30646 )  ;
assign n30776 =  ( n21 ) & ( n30616 )  ;
assign n30777 =  ( n21 ) & ( n30618 )  ;
assign n30778 =  ( n21 ) & ( n30620 )  ;
assign n30779 =  ( n21 ) & ( n30622 )  ;
assign n30780 =  ( n21 ) & ( n30624 )  ;
assign n30781 =  ( n21 ) & ( n30626 )  ;
assign n30782 =  ( n21 ) & ( n30628 )  ;
assign n30783 =  ( n21 ) & ( n30630 )  ;
assign n30784 =  ( n21 ) & ( n30632 )  ;
assign n30785 =  ( n21 ) & ( n30634 )  ;
assign n30786 =  ( n21 ) & ( n30636 )  ;
assign n30787 =  ( n21 ) & ( n30638 )  ;
assign n30788 =  ( n21 ) & ( n30640 )  ;
assign n30789 =  ( n21 ) & ( n30642 )  ;
assign n30790 =  ( n21 ) & ( n30644 )  ;
assign n30791 =  ( n21 ) & ( n30646 )  ;
assign n30792 =  ( n22 ) & ( n30616 )  ;
assign n30793 =  ( n22 ) & ( n30618 )  ;
assign n30794 =  ( n22 ) & ( n30620 )  ;
assign n30795 =  ( n22 ) & ( n30622 )  ;
assign n30796 =  ( n22 ) & ( n30624 )  ;
assign n30797 =  ( n22 ) & ( n30626 )  ;
assign n30798 =  ( n22 ) & ( n30628 )  ;
assign n30799 =  ( n22 ) & ( n30630 )  ;
assign n30800 =  ( n22 ) & ( n30632 )  ;
assign n30801 =  ( n22 ) & ( n30634 )  ;
assign n30802 =  ( n22 ) & ( n30636 )  ;
assign n30803 =  ( n22 ) & ( n30638 )  ;
assign n30804 =  ( n22 ) & ( n30640 )  ;
assign n30805 =  ( n22 ) & ( n30642 )  ;
assign n30806 =  ( n22 ) & ( n30644 )  ;
assign n30807 =  ( n22 ) & ( n30646 )  ;
assign n30808 =  ( n23 ) & ( n30616 )  ;
assign n30809 =  ( n23 ) & ( n30618 )  ;
assign n30810 =  ( n23 ) & ( n30620 )  ;
assign n30811 =  ( n23 ) & ( n30622 )  ;
assign n30812 =  ( n23 ) & ( n30624 )  ;
assign n30813 =  ( n23 ) & ( n30626 )  ;
assign n30814 =  ( n23 ) & ( n30628 )  ;
assign n30815 =  ( n23 ) & ( n30630 )  ;
assign n30816 =  ( n23 ) & ( n30632 )  ;
assign n30817 =  ( n23 ) & ( n30634 )  ;
assign n30818 =  ( n23 ) & ( n30636 )  ;
assign n30819 =  ( n23 ) & ( n30638 )  ;
assign n30820 =  ( n23 ) & ( n30640 )  ;
assign n30821 =  ( n23 ) & ( n30642 )  ;
assign n30822 =  ( n23 ) & ( n30644 )  ;
assign n30823 =  ( n23 ) & ( n30646 )  ;
assign n30824 =  ( n24 ) & ( n30616 )  ;
assign n30825 =  ( n24 ) & ( n30618 )  ;
assign n30826 =  ( n24 ) & ( n30620 )  ;
assign n30827 =  ( n24 ) & ( n30622 )  ;
assign n30828 =  ( n24 ) & ( n30624 )  ;
assign n30829 =  ( n24 ) & ( n30626 )  ;
assign n30830 =  ( n24 ) & ( n30628 )  ;
assign n30831 =  ( n24 ) & ( n30630 )  ;
assign n30832 =  ( n24 ) & ( n30632 )  ;
assign n30833 =  ( n24 ) & ( n30634 )  ;
assign n30834 =  ( n24 ) & ( n30636 )  ;
assign n30835 =  ( n24 ) & ( n30638 )  ;
assign n30836 =  ( n24 ) & ( n30640 )  ;
assign n30837 =  ( n24 ) & ( n30642 )  ;
assign n30838 =  ( n24 ) & ( n30644 )  ;
assign n30839 =  ( n24 ) & ( n30646 )  ;
assign n30840 =  ( n25 ) & ( n30616 )  ;
assign n30841 =  ( n25 ) & ( n30618 )  ;
assign n30842 =  ( n25 ) & ( n30620 )  ;
assign n30843 =  ( n25 ) & ( n30622 )  ;
assign n30844 =  ( n25 ) & ( n30624 )  ;
assign n30845 =  ( n25 ) & ( n30626 )  ;
assign n30846 =  ( n25 ) & ( n30628 )  ;
assign n30847 =  ( n25 ) & ( n30630 )  ;
assign n30848 =  ( n25 ) & ( n30632 )  ;
assign n30849 =  ( n25 ) & ( n30634 )  ;
assign n30850 =  ( n25 ) & ( n30636 )  ;
assign n30851 =  ( n25 ) & ( n30638 )  ;
assign n30852 =  ( n25 ) & ( n30640 )  ;
assign n30853 =  ( n25 ) & ( n30642 )  ;
assign n30854 =  ( n25 ) & ( n30644 )  ;
assign n30855 =  ( n25 ) & ( n30646 )  ;
assign n30856 =  ( n26 ) & ( n30616 )  ;
assign n30857 =  ( n26 ) & ( n30618 )  ;
assign n30858 =  ( n26 ) & ( n30620 )  ;
assign n30859 =  ( n26 ) & ( n30622 )  ;
assign n30860 =  ( n26 ) & ( n30624 )  ;
assign n30861 =  ( n26 ) & ( n30626 )  ;
assign n30862 =  ( n26 ) & ( n30628 )  ;
assign n30863 =  ( n26 ) & ( n30630 )  ;
assign n30864 =  ( n26 ) & ( n30632 )  ;
assign n30865 =  ( n26 ) & ( n30634 )  ;
assign n30866 =  ( n26 ) & ( n30636 )  ;
assign n30867 =  ( n26 ) & ( n30638 )  ;
assign n30868 =  ( n26 ) & ( n30640 )  ;
assign n30869 =  ( n26 ) & ( n30642 )  ;
assign n30870 =  ( n26 ) & ( n30644 )  ;
assign n30871 =  ( n26 ) & ( n30646 )  ;
assign n30872 =  ( n27 ) & ( n30616 )  ;
assign n30873 =  ( n27 ) & ( n30618 )  ;
assign n30874 =  ( n27 ) & ( n30620 )  ;
assign n30875 =  ( n27 ) & ( n30622 )  ;
assign n30876 =  ( n27 ) & ( n30624 )  ;
assign n30877 =  ( n27 ) & ( n30626 )  ;
assign n30878 =  ( n27 ) & ( n30628 )  ;
assign n30879 =  ( n27 ) & ( n30630 )  ;
assign n30880 =  ( n27 ) & ( n30632 )  ;
assign n30881 =  ( n27 ) & ( n30634 )  ;
assign n30882 =  ( n27 ) & ( n30636 )  ;
assign n30883 =  ( n27 ) & ( n30638 )  ;
assign n30884 =  ( n27 ) & ( n30640 )  ;
assign n30885 =  ( n27 ) & ( n30642 )  ;
assign n30886 =  ( n27 ) & ( n30644 )  ;
assign n30887 =  ( n27 ) & ( n30646 )  ;
assign n30888 =  ( n28 ) & ( n30616 )  ;
assign n30889 =  ( n28 ) & ( n30618 )  ;
assign n30890 =  ( n28 ) & ( n30620 )  ;
assign n30891 =  ( n28 ) & ( n30622 )  ;
assign n30892 =  ( n28 ) & ( n30624 )  ;
assign n30893 =  ( n28 ) & ( n30626 )  ;
assign n30894 =  ( n28 ) & ( n30628 )  ;
assign n30895 =  ( n28 ) & ( n30630 )  ;
assign n30896 =  ( n28 ) & ( n30632 )  ;
assign n30897 =  ( n28 ) & ( n30634 )  ;
assign n30898 =  ( n28 ) & ( n30636 )  ;
assign n30899 =  ( n28 ) & ( n30638 )  ;
assign n30900 =  ( n28 ) & ( n30640 )  ;
assign n30901 =  ( n28 ) & ( n30642 )  ;
assign n30902 =  ( n28 ) & ( n30644 )  ;
assign n30903 =  ( n28 ) & ( n30646 )  ;
assign n30904 =  ( n29 ) & ( n30616 )  ;
assign n30905 =  ( n29 ) & ( n30618 )  ;
assign n30906 =  ( n29 ) & ( n30620 )  ;
assign n30907 =  ( n29 ) & ( n30622 )  ;
assign n30908 =  ( n29 ) & ( n30624 )  ;
assign n30909 =  ( n29 ) & ( n30626 )  ;
assign n30910 =  ( n29 ) & ( n30628 )  ;
assign n30911 =  ( n29 ) & ( n30630 )  ;
assign n30912 =  ( n29 ) & ( n30632 )  ;
assign n30913 =  ( n29 ) & ( n30634 )  ;
assign n30914 =  ( n29 ) & ( n30636 )  ;
assign n30915 =  ( n29 ) & ( n30638 )  ;
assign n30916 =  ( n29 ) & ( n30640 )  ;
assign n30917 =  ( n29 ) & ( n30642 )  ;
assign n30918 =  ( n29 ) & ( n30644 )  ;
assign n30919 =  ( n29 ) & ( n30646 )  ;
assign n30920 =  ( n30 ) & ( n30616 )  ;
assign n30921 =  ( n30 ) & ( n30618 )  ;
assign n30922 =  ( n30 ) & ( n30620 )  ;
assign n30923 =  ( n30 ) & ( n30622 )  ;
assign n30924 =  ( n30 ) & ( n30624 )  ;
assign n30925 =  ( n30 ) & ( n30626 )  ;
assign n30926 =  ( n30 ) & ( n30628 )  ;
assign n30927 =  ( n30 ) & ( n30630 )  ;
assign n30928 =  ( n30 ) & ( n30632 )  ;
assign n30929 =  ( n30 ) & ( n30634 )  ;
assign n30930 =  ( n30 ) & ( n30636 )  ;
assign n30931 =  ( n30 ) & ( n30638 )  ;
assign n30932 =  ( n30 ) & ( n30640 )  ;
assign n30933 =  ( n30 ) & ( n30642 )  ;
assign n30934 =  ( n30 ) & ( n30644 )  ;
assign n30935 =  ( n30 ) & ( n30646 )  ;
assign n30936 =  ( n31 ) & ( n30616 )  ;
assign n30937 =  ( n31 ) & ( n30618 )  ;
assign n30938 =  ( n31 ) & ( n30620 )  ;
assign n30939 =  ( n31 ) & ( n30622 )  ;
assign n30940 =  ( n31 ) & ( n30624 )  ;
assign n30941 =  ( n31 ) & ( n30626 )  ;
assign n30942 =  ( n31 ) & ( n30628 )  ;
assign n30943 =  ( n31 ) & ( n30630 )  ;
assign n30944 =  ( n31 ) & ( n30632 )  ;
assign n30945 =  ( n31 ) & ( n30634 )  ;
assign n30946 =  ( n31 ) & ( n30636 )  ;
assign n30947 =  ( n31 ) & ( n30638 )  ;
assign n30948 =  ( n31 ) & ( n30640 )  ;
assign n30949 =  ( n31 ) & ( n30642 )  ;
assign n30950 =  ( n31 ) & ( n30644 )  ;
assign n30951 =  ( n31 ) & ( n30646 )  ;
assign n30952 =  ( n32 ) & ( n30616 )  ;
assign n30953 =  ( n32 ) & ( n30618 )  ;
assign n30954 =  ( n32 ) & ( n30620 )  ;
assign n30955 =  ( n32 ) & ( n30622 )  ;
assign n30956 =  ( n32 ) & ( n30624 )  ;
assign n30957 =  ( n32 ) & ( n30626 )  ;
assign n30958 =  ( n32 ) & ( n30628 )  ;
assign n30959 =  ( n32 ) & ( n30630 )  ;
assign n30960 =  ( n32 ) & ( n30632 )  ;
assign n30961 =  ( n32 ) & ( n30634 )  ;
assign n30962 =  ( n32 ) & ( n30636 )  ;
assign n30963 =  ( n32 ) & ( n30638 )  ;
assign n30964 =  ( n32 ) & ( n30640 )  ;
assign n30965 =  ( n32 ) & ( n30642 )  ;
assign n30966 =  ( n32 ) & ( n30644 )  ;
assign n30967 =  ( n32 ) & ( n30646 )  ;
assign n30968 =  ( n33 ) & ( n30616 )  ;
assign n30969 =  ( n33 ) & ( n30618 )  ;
assign n30970 =  ( n33 ) & ( n30620 )  ;
assign n30971 =  ( n33 ) & ( n30622 )  ;
assign n30972 =  ( n33 ) & ( n30624 )  ;
assign n30973 =  ( n33 ) & ( n30626 )  ;
assign n30974 =  ( n33 ) & ( n30628 )  ;
assign n30975 =  ( n33 ) & ( n30630 )  ;
assign n30976 =  ( n33 ) & ( n30632 )  ;
assign n30977 =  ( n33 ) & ( n30634 )  ;
assign n30978 =  ( n33 ) & ( n30636 )  ;
assign n30979 =  ( n33 ) & ( n30638 )  ;
assign n30980 =  ( n33 ) & ( n30640 )  ;
assign n30981 =  ( n33 ) & ( n30642 )  ;
assign n30982 =  ( n33 ) & ( n30644 )  ;
assign n30983 =  ( n33 ) & ( n30646 )  ;
assign n30984 =  ( n34 ) & ( n30616 )  ;
assign n30985 =  ( n34 ) & ( n30618 )  ;
assign n30986 =  ( n34 ) & ( n30620 )  ;
assign n30987 =  ( n34 ) & ( n30622 )  ;
assign n30988 =  ( n34 ) & ( n30624 )  ;
assign n30989 =  ( n34 ) & ( n30626 )  ;
assign n30990 =  ( n34 ) & ( n30628 )  ;
assign n30991 =  ( n34 ) & ( n30630 )  ;
assign n30992 =  ( n34 ) & ( n30632 )  ;
assign n30993 =  ( n34 ) & ( n30634 )  ;
assign n30994 =  ( n34 ) & ( n30636 )  ;
assign n30995 =  ( n34 ) & ( n30638 )  ;
assign n30996 =  ( n34 ) & ( n30640 )  ;
assign n30997 =  ( n34 ) & ( n30642 )  ;
assign n30998 =  ( n34 ) & ( n30644 )  ;
assign n30999 =  ( n34 ) & ( n30646 )  ;
assign n31000 =  ( n35 ) & ( n30616 )  ;
assign n31001 =  ( n35 ) & ( n30618 )  ;
assign n31002 =  ( n35 ) & ( n30620 )  ;
assign n31003 =  ( n35 ) & ( n30622 )  ;
assign n31004 =  ( n35 ) & ( n30624 )  ;
assign n31005 =  ( n35 ) & ( n30626 )  ;
assign n31006 =  ( n35 ) & ( n30628 )  ;
assign n31007 =  ( n35 ) & ( n30630 )  ;
assign n31008 =  ( n35 ) & ( n30632 )  ;
assign n31009 =  ( n35 ) & ( n30634 )  ;
assign n31010 =  ( n35 ) & ( n30636 )  ;
assign n31011 =  ( n35 ) & ( n30638 )  ;
assign n31012 =  ( n35 ) & ( n30640 )  ;
assign n31013 =  ( n35 ) & ( n30642 )  ;
assign n31014 =  ( n35 ) & ( n30644 )  ;
assign n31015 =  ( n35 ) & ( n30646 )  ;
assign n31016 =  ( n36 ) & ( n30616 )  ;
assign n31017 =  ( n36 ) & ( n30618 )  ;
assign n31018 =  ( n36 ) & ( n30620 )  ;
assign n31019 =  ( n36 ) & ( n30622 )  ;
assign n31020 =  ( n36 ) & ( n30624 )  ;
assign n31021 =  ( n36 ) & ( n30626 )  ;
assign n31022 =  ( n36 ) & ( n30628 )  ;
assign n31023 =  ( n36 ) & ( n30630 )  ;
assign n31024 =  ( n36 ) & ( n30632 )  ;
assign n31025 =  ( n36 ) & ( n30634 )  ;
assign n31026 =  ( n36 ) & ( n30636 )  ;
assign n31027 =  ( n36 ) & ( n30638 )  ;
assign n31028 =  ( n36 ) & ( n30640 )  ;
assign n31029 =  ( n36 ) & ( n30642 )  ;
assign n31030 =  ( n36 ) & ( n30644 )  ;
assign n31031 =  ( n36 ) & ( n30646 )  ;
assign n31032 =  ( n37 ) & ( n30616 )  ;
assign n31033 =  ( n37 ) & ( n30618 )  ;
assign n31034 =  ( n37 ) & ( n30620 )  ;
assign n31035 =  ( n37 ) & ( n30622 )  ;
assign n31036 =  ( n37 ) & ( n30624 )  ;
assign n31037 =  ( n37 ) & ( n30626 )  ;
assign n31038 =  ( n37 ) & ( n30628 )  ;
assign n31039 =  ( n37 ) & ( n30630 )  ;
assign n31040 =  ( n37 ) & ( n30632 )  ;
assign n31041 =  ( n37 ) & ( n30634 )  ;
assign n31042 =  ( n37 ) & ( n30636 )  ;
assign n31043 =  ( n37 ) & ( n30638 )  ;
assign n31044 =  ( n37 ) & ( n30640 )  ;
assign n31045 =  ( n37 ) & ( n30642 )  ;
assign n31046 =  ( n37 ) & ( n30644 )  ;
assign n31047 =  ( n37 ) & ( n30646 )  ;
assign n31048 =  ( n38 ) & ( n30616 )  ;
assign n31049 =  ( n38 ) & ( n30618 )  ;
assign n31050 =  ( n38 ) & ( n30620 )  ;
assign n31051 =  ( n38 ) & ( n30622 )  ;
assign n31052 =  ( n38 ) & ( n30624 )  ;
assign n31053 =  ( n38 ) & ( n30626 )  ;
assign n31054 =  ( n38 ) & ( n30628 )  ;
assign n31055 =  ( n38 ) & ( n30630 )  ;
assign n31056 =  ( n38 ) & ( n30632 )  ;
assign n31057 =  ( n38 ) & ( n30634 )  ;
assign n31058 =  ( n38 ) & ( n30636 )  ;
assign n31059 =  ( n38 ) & ( n30638 )  ;
assign n31060 =  ( n38 ) & ( n30640 )  ;
assign n31061 =  ( n38 ) & ( n30642 )  ;
assign n31062 =  ( n38 ) & ( n30644 )  ;
assign n31063 =  ( n38 ) & ( n30646 )  ;
assign n31064 =  ( n39 ) & ( n30616 )  ;
assign n31065 =  ( n39 ) & ( n30618 )  ;
assign n31066 =  ( n39 ) & ( n30620 )  ;
assign n31067 =  ( n39 ) & ( n30622 )  ;
assign n31068 =  ( n39 ) & ( n30624 )  ;
assign n31069 =  ( n39 ) & ( n30626 )  ;
assign n31070 =  ( n39 ) & ( n30628 )  ;
assign n31071 =  ( n39 ) & ( n30630 )  ;
assign n31072 =  ( n39 ) & ( n30632 )  ;
assign n31073 =  ( n39 ) & ( n30634 )  ;
assign n31074 =  ( n39 ) & ( n30636 )  ;
assign n31075 =  ( n39 ) & ( n30638 )  ;
assign n31076 =  ( n39 ) & ( n30640 )  ;
assign n31077 =  ( n39 ) & ( n30642 )  ;
assign n31078 =  ( n39 ) & ( n30644 )  ;
assign n31079 =  ( n39 ) & ( n30646 )  ;
assign n31080 =  ( n40 ) & ( n30616 )  ;
assign n31081 =  ( n40 ) & ( n30618 )  ;
assign n31082 =  ( n40 ) & ( n30620 )  ;
assign n31083 =  ( n40 ) & ( n30622 )  ;
assign n31084 =  ( n40 ) & ( n30624 )  ;
assign n31085 =  ( n40 ) & ( n30626 )  ;
assign n31086 =  ( n40 ) & ( n30628 )  ;
assign n31087 =  ( n40 ) & ( n30630 )  ;
assign n31088 =  ( n40 ) & ( n30632 )  ;
assign n31089 =  ( n40 ) & ( n30634 )  ;
assign n31090 =  ( n40 ) & ( n30636 )  ;
assign n31091 =  ( n40 ) & ( n30638 )  ;
assign n31092 =  ( n40 ) & ( n30640 )  ;
assign n31093 =  ( n40 ) & ( n30642 )  ;
assign n31094 =  ( n40 ) & ( n30644 )  ;
assign n31095 =  ( n40 ) & ( n30646 )  ;
assign n31096 =  ( n41 ) & ( n30616 )  ;
assign n31097 =  ( n41 ) & ( n30618 )  ;
assign n31098 =  ( n41 ) & ( n30620 )  ;
assign n31099 =  ( n41 ) & ( n30622 )  ;
assign n31100 =  ( n41 ) & ( n30624 )  ;
assign n31101 =  ( n41 ) & ( n30626 )  ;
assign n31102 =  ( n41 ) & ( n30628 )  ;
assign n31103 =  ( n41 ) & ( n30630 )  ;
assign n31104 =  ( n41 ) & ( n30632 )  ;
assign n31105 =  ( n41 ) & ( n30634 )  ;
assign n31106 =  ( n41 ) & ( n30636 )  ;
assign n31107 =  ( n41 ) & ( n30638 )  ;
assign n31108 =  ( n41 ) & ( n30640 )  ;
assign n31109 =  ( n41 ) & ( n30642 )  ;
assign n31110 =  ( n41 ) & ( n30644 )  ;
assign n31111 =  ( n41 ) & ( n30646 )  ;
assign n31112 =  ( n42 ) & ( n30616 )  ;
assign n31113 =  ( n42 ) & ( n30618 )  ;
assign n31114 =  ( n42 ) & ( n30620 )  ;
assign n31115 =  ( n42 ) & ( n30622 )  ;
assign n31116 =  ( n42 ) & ( n30624 )  ;
assign n31117 =  ( n42 ) & ( n30626 )  ;
assign n31118 =  ( n42 ) & ( n30628 )  ;
assign n31119 =  ( n42 ) & ( n30630 )  ;
assign n31120 =  ( n42 ) & ( n30632 )  ;
assign n31121 =  ( n42 ) & ( n30634 )  ;
assign n31122 =  ( n42 ) & ( n30636 )  ;
assign n31123 =  ( n42 ) & ( n30638 )  ;
assign n31124 =  ( n42 ) & ( n30640 )  ;
assign n31125 =  ( n42 ) & ( n30642 )  ;
assign n31126 =  ( n42 ) & ( n30644 )  ;
assign n31127 =  ( n42 ) & ( n30646 )  ;
assign n31128 =  ( n43 ) & ( n30616 )  ;
assign n31129 =  ( n43 ) & ( n30618 )  ;
assign n31130 =  ( n43 ) & ( n30620 )  ;
assign n31131 =  ( n43 ) & ( n30622 )  ;
assign n31132 =  ( n43 ) & ( n30624 )  ;
assign n31133 =  ( n43 ) & ( n30626 )  ;
assign n31134 =  ( n43 ) & ( n30628 )  ;
assign n31135 =  ( n43 ) & ( n30630 )  ;
assign n31136 =  ( n43 ) & ( n30632 )  ;
assign n31137 =  ( n43 ) & ( n30634 )  ;
assign n31138 =  ( n43 ) & ( n30636 )  ;
assign n31139 =  ( n43 ) & ( n30638 )  ;
assign n31140 =  ( n43 ) & ( n30640 )  ;
assign n31141 =  ( n43 ) & ( n30642 )  ;
assign n31142 =  ( n43 ) & ( n30644 )  ;
assign n31143 =  ( n43 ) & ( n30646 )  ;
assign n31144 =  ( n31143 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n31145 =  ( n31142 ) ? ( VREG_0_1 ) : ( n31144 ) ;
assign n31146 =  ( n31141 ) ? ( VREG_0_2 ) : ( n31145 ) ;
assign n31147 =  ( n31140 ) ? ( VREG_0_3 ) : ( n31146 ) ;
assign n31148 =  ( n31139 ) ? ( VREG_0_4 ) : ( n31147 ) ;
assign n31149 =  ( n31138 ) ? ( VREG_0_5 ) : ( n31148 ) ;
assign n31150 =  ( n31137 ) ? ( VREG_0_6 ) : ( n31149 ) ;
assign n31151 =  ( n31136 ) ? ( VREG_0_7 ) : ( n31150 ) ;
assign n31152 =  ( n31135 ) ? ( VREG_0_8 ) : ( n31151 ) ;
assign n31153 =  ( n31134 ) ? ( VREG_0_9 ) : ( n31152 ) ;
assign n31154 =  ( n31133 ) ? ( VREG_0_10 ) : ( n31153 ) ;
assign n31155 =  ( n31132 ) ? ( VREG_0_11 ) : ( n31154 ) ;
assign n31156 =  ( n31131 ) ? ( VREG_0_12 ) : ( n31155 ) ;
assign n31157 =  ( n31130 ) ? ( VREG_0_13 ) : ( n31156 ) ;
assign n31158 =  ( n31129 ) ? ( VREG_0_14 ) : ( n31157 ) ;
assign n31159 =  ( n31128 ) ? ( VREG_0_15 ) : ( n31158 ) ;
assign n31160 =  ( n31127 ) ? ( VREG_1_0 ) : ( n31159 ) ;
assign n31161 =  ( n31126 ) ? ( VREG_1_1 ) : ( n31160 ) ;
assign n31162 =  ( n31125 ) ? ( VREG_1_2 ) : ( n31161 ) ;
assign n31163 =  ( n31124 ) ? ( VREG_1_3 ) : ( n31162 ) ;
assign n31164 =  ( n31123 ) ? ( VREG_1_4 ) : ( n31163 ) ;
assign n31165 =  ( n31122 ) ? ( VREG_1_5 ) : ( n31164 ) ;
assign n31166 =  ( n31121 ) ? ( VREG_1_6 ) : ( n31165 ) ;
assign n31167 =  ( n31120 ) ? ( VREG_1_7 ) : ( n31166 ) ;
assign n31168 =  ( n31119 ) ? ( VREG_1_8 ) : ( n31167 ) ;
assign n31169 =  ( n31118 ) ? ( VREG_1_9 ) : ( n31168 ) ;
assign n31170 =  ( n31117 ) ? ( VREG_1_10 ) : ( n31169 ) ;
assign n31171 =  ( n31116 ) ? ( VREG_1_11 ) : ( n31170 ) ;
assign n31172 =  ( n31115 ) ? ( VREG_1_12 ) : ( n31171 ) ;
assign n31173 =  ( n31114 ) ? ( VREG_1_13 ) : ( n31172 ) ;
assign n31174 =  ( n31113 ) ? ( VREG_1_14 ) : ( n31173 ) ;
assign n31175 =  ( n31112 ) ? ( VREG_1_15 ) : ( n31174 ) ;
assign n31176 =  ( n31111 ) ? ( VREG_2_0 ) : ( n31175 ) ;
assign n31177 =  ( n31110 ) ? ( VREG_2_1 ) : ( n31176 ) ;
assign n31178 =  ( n31109 ) ? ( VREG_2_2 ) : ( n31177 ) ;
assign n31179 =  ( n31108 ) ? ( VREG_2_3 ) : ( n31178 ) ;
assign n31180 =  ( n31107 ) ? ( VREG_2_4 ) : ( n31179 ) ;
assign n31181 =  ( n31106 ) ? ( VREG_2_5 ) : ( n31180 ) ;
assign n31182 =  ( n31105 ) ? ( VREG_2_6 ) : ( n31181 ) ;
assign n31183 =  ( n31104 ) ? ( VREG_2_7 ) : ( n31182 ) ;
assign n31184 =  ( n31103 ) ? ( VREG_2_8 ) : ( n31183 ) ;
assign n31185 =  ( n31102 ) ? ( VREG_2_9 ) : ( n31184 ) ;
assign n31186 =  ( n31101 ) ? ( VREG_2_10 ) : ( n31185 ) ;
assign n31187 =  ( n31100 ) ? ( VREG_2_11 ) : ( n31186 ) ;
assign n31188 =  ( n31099 ) ? ( VREG_2_12 ) : ( n31187 ) ;
assign n31189 =  ( n31098 ) ? ( VREG_2_13 ) : ( n31188 ) ;
assign n31190 =  ( n31097 ) ? ( VREG_2_14 ) : ( n31189 ) ;
assign n31191 =  ( n31096 ) ? ( VREG_2_15 ) : ( n31190 ) ;
assign n31192 =  ( n31095 ) ? ( VREG_3_0 ) : ( n31191 ) ;
assign n31193 =  ( n31094 ) ? ( VREG_3_1 ) : ( n31192 ) ;
assign n31194 =  ( n31093 ) ? ( VREG_3_2 ) : ( n31193 ) ;
assign n31195 =  ( n31092 ) ? ( VREG_3_3 ) : ( n31194 ) ;
assign n31196 =  ( n31091 ) ? ( VREG_3_4 ) : ( n31195 ) ;
assign n31197 =  ( n31090 ) ? ( VREG_3_5 ) : ( n31196 ) ;
assign n31198 =  ( n31089 ) ? ( VREG_3_6 ) : ( n31197 ) ;
assign n31199 =  ( n31088 ) ? ( VREG_3_7 ) : ( n31198 ) ;
assign n31200 =  ( n31087 ) ? ( VREG_3_8 ) : ( n31199 ) ;
assign n31201 =  ( n31086 ) ? ( VREG_3_9 ) : ( n31200 ) ;
assign n31202 =  ( n31085 ) ? ( VREG_3_10 ) : ( n31201 ) ;
assign n31203 =  ( n31084 ) ? ( VREG_3_11 ) : ( n31202 ) ;
assign n31204 =  ( n31083 ) ? ( VREG_3_12 ) : ( n31203 ) ;
assign n31205 =  ( n31082 ) ? ( VREG_3_13 ) : ( n31204 ) ;
assign n31206 =  ( n31081 ) ? ( VREG_3_14 ) : ( n31205 ) ;
assign n31207 =  ( n31080 ) ? ( VREG_3_15 ) : ( n31206 ) ;
assign n31208 =  ( n31079 ) ? ( VREG_4_0 ) : ( n31207 ) ;
assign n31209 =  ( n31078 ) ? ( VREG_4_1 ) : ( n31208 ) ;
assign n31210 =  ( n31077 ) ? ( VREG_4_2 ) : ( n31209 ) ;
assign n31211 =  ( n31076 ) ? ( VREG_4_3 ) : ( n31210 ) ;
assign n31212 =  ( n31075 ) ? ( VREG_4_4 ) : ( n31211 ) ;
assign n31213 =  ( n31074 ) ? ( VREG_4_5 ) : ( n31212 ) ;
assign n31214 =  ( n31073 ) ? ( VREG_4_6 ) : ( n31213 ) ;
assign n31215 =  ( n31072 ) ? ( VREG_4_7 ) : ( n31214 ) ;
assign n31216 =  ( n31071 ) ? ( VREG_4_8 ) : ( n31215 ) ;
assign n31217 =  ( n31070 ) ? ( VREG_4_9 ) : ( n31216 ) ;
assign n31218 =  ( n31069 ) ? ( VREG_4_10 ) : ( n31217 ) ;
assign n31219 =  ( n31068 ) ? ( VREG_4_11 ) : ( n31218 ) ;
assign n31220 =  ( n31067 ) ? ( VREG_4_12 ) : ( n31219 ) ;
assign n31221 =  ( n31066 ) ? ( VREG_4_13 ) : ( n31220 ) ;
assign n31222 =  ( n31065 ) ? ( VREG_4_14 ) : ( n31221 ) ;
assign n31223 =  ( n31064 ) ? ( VREG_4_15 ) : ( n31222 ) ;
assign n31224 =  ( n31063 ) ? ( VREG_5_0 ) : ( n31223 ) ;
assign n31225 =  ( n31062 ) ? ( VREG_5_1 ) : ( n31224 ) ;
assign n31226 =  ( n31061 ) ? ( VREG_5_2 ) : ( n31225 ) ;
assign n31227 =  ( n31060 ) ? ( VREG_5_3 ) : ( n31226 ) ;
assign n31228 =  ( n31059 ) ? ( VREG_5_4 ) : ( n31227 ) ;
assign n31229 =  ( n31058 ) ? ( VREG_5_5 ) : ( n31228 ) ;
assign n31230 =  ( n31057 ) ? ( VREG_5_6 ) : ( n31229 ) ;
assign n31231 =  ( n31056 ) ? ( VREG_5_7 ) : ( n31230 ) ;
assign n31232 =  ( n31055 ) ? ( VREG_5_8 ) : ( n31231 ) ;
assign n31233 =  ( n31054 ) ? ( VREG_5_9 ) : ( n31232 ) ;
assign n31234 =  ( n31053 ) ? ( VREG_5_10 ) : ( n31233 ) ;
assign n31235 =  ( n31052 ) ? ( VREG_5_11 ) : ( n31234 ) ;
assign n31236 =  ( n31051 ) ? ( VREG_5_12 ) : ( n31235 ) ;
assign n31237 =  ( n31050 ) ? ( VREG_5_13 ) : ( n31236 ) ;
assign n31238 =  ( n31049 ) ? ( VREG_5_14 ) : ( n31237 ) ;
assign n31239 =  ( n31048 ) ? ( VREG_5_15 ) : ( n31238 ) ;
assign n31240 =  ( n31047 ) ? ( VREG_6_0 ) : ( n31239 ) ;
assign n31241 =  ( n31046 ) ? ( VREG_6_1 ) : ( n31240 ) ;
assign n31242 =  ( n31045 ) ? ( VREG_6_2 ) : ( n31241 ) ;
assign n31243 =  ( n31044 ) ? ( VREG_6_3 ) : ( n31242 ) ;
assign n31244 =  ( n31043 ) ? ( VREG_6_4 ) : ( n31243 ) ;
assign n31245 =  ( n31042 ) ? ( VREG_6_5 ) : ( n31244 ) ;
assign n31246 =  ( n31041 ) ? ( VREG_6_6 ) : ( n31245 ) ;
assign n31247 =  ( n31040 ) ? ( VREG_6_7 ) : ( n31246 ) ;
assign n31248 =  ( n31039 ) ? ( VREG_6_8 ) : ( n31247 ) ;
assign n31249 =  ( n31038 ) ? ( VREG_6_9 ) : ( n31248 ) ;
assign n31250 =  ( n31037 ) ? ( VREG_6_10 ) : ( n31249 ) ;
assign n31251 =  ( n31036 ) ? ( VREG_6_11 ) : ( n31250 ) ;
assign n31252 =  ( n31035 ) ? ( VREG_6_12 ) : ( n31251 ) ;
assign n31253 =  ( n31034 ) ? ( VREG_6_13 ) : ( n31252 ) ;
assign n31254 =  ( n31033 ) ? ( VREG_6_14 ) : ( n31253 ) ;
assign n31255 =  ( n31032 ) ? ( VREG_6_15 ) : ( n31254 ) ;
assign n31256 =  ( n31031 ) ? ( VREG_7_0 ) : ( n31255 ) ;
assign n31257 =  ( n31030 ) ? ( VREG_7_1 ) : ( n31256 ) ;
assign n31258 =  ( n31029 ) ? ( VREG_7_2 ) : ( n31257 ) ;
assign n31259 =  ( n31028 ) ? ( VREG_7_3 ) : ( n31258 ) ;
assign n31260 =  ( n31027 ) ? ( VREG_7_4 ) : ( n31259 ) ;
assign n31261 =  ( n31026 ) ? ( VREG_7_5 ) : ( n31260 ) ;
assign n31262 =  ( n31025 ) ? ( VREG_7_6 ) : ( n31261 ) ;
assign n31263 =  ( n31024 ) ? ( VREG_7_7 ) : ( n31262 ) ;
assign n31264 =  ( n31023 ) ? ( VREG_7_8 ) : ( n31263 ) ;
assign n31265 =  ( n31022 ) ? ( VREG_7_9 ) : ( n31264 ) ;
assign n31266 =  ( n31021 ) ? ( VREG_7_10 ) : ( n31265 ) ;
assign n31267 =  ( n31020 ) ? ( VREG_7_11 ) : ( n31266 ) ;
assign n31268 =  ( n31019 ) ? ( VREG_7_12 ) : ( n31267 ) ;
assign n31269 =  ( n31018 ) ? ( VREG_7_13 ) : ( n31268 ) ;
assign n31270 =  ( n31017 ) ? ( VREG_7_14 ) : ( n31269 ) ;
assign n31271 =  ( n31016 ) ? ( VREG_7_15 ) : ( n31270 ) ;
assign n31272 =  ( n31015 ) ? ( VREG_8_0 ) : ( n31271 ) ;
assign n31273 =  ( n31014 ) ? ( VREG_8_1 ) : ( n31272 ) ;
assign n31274 =  ( n31013 ) ? ( VREG_8_2 ) : ( n31273 ) ;
assign n31275 =  ( n31012 ) ? ( VREG_8_3 ) : ( n31274 ) ;
assign n31276 =  ( n31011 ) ? ( VREG_8_4 ) : ( n31275 ) ;
assign n31277 =  ( n31010 ) ? ( VREG_8_5 ) : ( n31276 ) ;
assign n31278 =  ( n31009 ) ? ( VREG_8_6 ) : ( n31277 ) ;
assign n31279 =  ( n31008 ) ? ( VREG_8_7 ) : ( n31278 ) ;
assign n31280 =  ( n31007 ) ? ( VREG_8_8 ) : ( n31279 ) ;
assign n31281 =  ( n31006 ) ? ( VREG_8_9 ) : ( n31280 ) ;
assign n31282 =  ( n31005 ) ? ( VREG_8_10 ) : ( n31281 ) ;
assign n31283 =  ( n31004 ) ? ( VREG_8_11 ) : ( n31282 ) ;
assign n31284 =  ( n31003 ) ? ( VREG_8_12 ) : ( n31283 ) ;
assign n31285 =  ( n31002 ) ? ( VREG_8_13 ) : ( n31284 ) ;
assign n31286 =  ( n31001 ) ? ( VREG_8_14 ) : ( n31285 ) ;
assign n31287 =  ( n31000 ) ? ( VREG_8_15 ) : ( n31286 ) ;
assign n31288 =  ( n30999 ) ? ( VREG_9_0 ) : ( n31287 ) ;
assign n31289 =  ( n30998 ) ? ( VREG_9_1 ) : ( n31288 ) ;
assign n31290 =  ( n30997 ) ? ( VREG_9_2 ) : ( n31289 ) ;
assign n31291 =  ( n30996 ) ? ( VREG_9_3 ) : ( n31290 ) ;
assign n31292 =  ( n30995 ) ? ( VREG_9_4 ) : ( n31291 ) ;
assign n31293 =  ( n30994 ) ? ( VREG_9_5 ) : ( n31292 ) ;
assign n31294 =  ( n30993 ) ? ( VREG_9_6 ) : ( n31293 ) ;
assign n31295 =  ( n30992 ) ? ( VREG_9_7 ) : ( n31294 ) ;
assign n31296 =  ( n30991 ) ? ( VREG_9_8 ) : ( n31295 ) ;
assign n31297 =  ( n30990 ) ? ( VREG_9_9 ) : ( n31296 ) ;
assign n31298 =  ( n30989 ) ? ( VREG_9_10 ) : ( n31297 ) ;
assign n31299 =  ( n30988 ) ? ( VREG_9_11 ) : ( n31298 ) ;
assign n31300 =  ( n30987 ) ? ( VREG_9_12 ) : ( n31299 ) ;
assign n31301 =  ( n30986 ) ? ( VREG_9_13 ) : ( n31300 ) ;
assign n31302 =  ( n30985 ) ? ( VREG_9_14 ) : ( n31301 ) ;
assign n31303 =  ( n30984 ) ? ( VREG_9_15 ) : ( n31302 ) ;
assign n31304 =  ( n30983 ) ? ( VREG_10_0 ) : ( n31303 ) ;
assign n31305 =  ( n30982 ) ? ( VREG_10_1 ) : ( n31304 ) ;
assign n31306 =  ( n30981 ) ? ( VREG_10_2 ) : ( n31305 ) ;
assign n31307 =  ( n30980 ) ? ( VREG_10_3 ) : ( n31306 ) ;
assign n31308 =  ( n30979 ) ? ( VREG_10_4 ) : ( n31307 ) ;
assign n31309 =  ( n30978 ) ? ( VREG_10_5 ) : ( n31308 ) ;
assign n31310 =  ( n30977 ) ? ( VREG_10_6 ) : ( n31309 ) ;
assign n31311 =  ( n30976 ) ? ( VREG_10_7 ) : ( n31310 ) ;
assign n31312 =  ( n30975 ) ? ( VREG_10_8 ) : ( n31311 ) ;
assign n31313 =  ( n30974 ) ? ( VREG_10_9 ) : ( n31312 ) ;
assign n31314 =  ( n30973 ) ? ( VREG_10_10 ) : ( n31313 ) ;
assign n31315 =  ( n30972 ) ? ( VREG_10_11 ) : ( n31314 ) ;
assign n31316 =  ( n30971 ) ? ( VREG_10_12 ) : ( n31315 ) ;
assign n31317 =  ( n30970 ) ? ( VREG_10_13 ) : ( n31316 ) ;
assign n31318 =  ( n30969 ) ? ( VREG_10_14 ) : ( n31317 ) ;
assign n31319 =  ( n30968 ) ? ( VREG_10_15 ) : ( n31318 ) ;
assign n31320 =  ( n30967 ) ? ( VREG_11_0 ) : ( n31319 ) ;
assign n31321 =  ( n30966 ) ? ( VREG_11_1 ) : ( n31320 ) ;
assign n31322 =  ( n30965 ) ? ( VREG_11_2 ) : ( n31321 ) ;
assign n31323 =  ( n30964 ) ? ( VREG_11_3 ) : ( n31322 ) ;
assign n31324 =  ( n30963 ) ? ( VREG_11_4 ) : ( n31323 ) ;
assign n31325 =  ( n30962 ) ? ( VREG_11_5 ) : ( n31324 ) ;
assign n31326 =  ( n30961 ) ? ( VREG_11_6 ) : ( n31325 ) ;
assign n31327 =  ( n30960 ) ? ( VREG_11_7 ) : ( n31326 ) ;
assign n31328 =  ( n30959 ) ? ( VREG_11_8 ) : ( n31327 ) ;
assign n31329 =  ( n30958 ) ? ( VREG_11_9 ) : ( n31328 ) ;
assign n31330 =  ( n30957 ) ? ( VREG_11_10 ) : ( n31329 ) ;
assign n31331 =  ( n30956 ) ? ( VREG_11_11 ) : ( n31330 ) ;
assign n31332 =  ( n30955 ) ? ( VREG_11_12 ) : ( n31331 ) ;
assign n31333 =  ( n30954 ) ? ( VREG_11_13 ) : ( n31332 ) ;
assign n31334 =  ( n30953 ) ? ( VREG_11_14 ) : ( n31333 ) ;
assign n31335 =  ( n30952 ) ? ( VREG_11_15 ) : ( n31334 ) ;
assign n31336 =  ( n30951 ) ? ( VREG_12_0 ) : ( n31335 ) ;
assign n31337 =  ( n30950 ) ? ( VREG_12_1 ) : ( n31336 ) ;
assign n31338 =  ( n30949 ) ? ( VREG_12_2 ) : ( n31337 ) ;
assign n31339 =  ( n30948 ) ? ( VREG_12_3 ) : ( n31338 ) ;
assign n31340 =  ( n30947 ) ? ( VREG_12_4 ) : ( n31339 ) ;
assign n31341 =  ( n30946 ) ? ( VREG_12_5 ) : ( n31340 ) ;
assign n31342 =  ( n30945 ) ? ( VREG_12_6 ) : ( n31341 ) ;
assign n31343 =  ( n30944 ) ? ( VREG_12_7 ) : ( n31342 ) ;
assign n31344 =  ( n30943 ) ? ( VREG_12_8 ) : ( n31343 ) ;
assign n31345 =  ( n30942 ) ? ( VREG_12_9 ) : ( n31344 ) ;
assign n31346 =  ( n30941 ) ? ( VREG_12_10 ) : ( n31345 ) ;
assign n31347 =  ( n30940 ) ? ( VREG_12_11 ) : ( n31346 ) ;
assign n31348 =  ( n30939 ) ? ( VREG_12_12 ) : ( n31347 ) ;
assign n31349 =  ( n30938 ) ? ( VREG_12_13 ) : ( n31348 ) ;
assign n31350 =  ( n30937 ) ? ( VREG_12_14 ) : ( n31349 ) ;
assign n31351 =  ( n30936 ) ? ( VREG_12_15 ) : ( n31350 ) ;
assign n31352 =  ( n30935 ) ? ( VREG_13_0 ) : ( n31351 ) ;
assign n31353 =  ( n30934 ) ? ( VREG_13_1 ) : ( n31352 ) ;
assign n31354 =  ( n30933 ) ? ( VREG_13_2 ) : ( n31353 ) ;
assign n31355 =  ( n30932 ) ? ( VREG_13_3 ) : ( n31354 ) ;
assign n31356 =  ( n30931 ) ? ( VREG_13_4 ) : ( n31355 ) ;
assign n31357 =  ( n30930 ) ? ( VREG_13_5 ) : ( n31356 ) ;
assign n31358 =  ( n30929 ) ? ( VREG_13_6 ) : ( n31357 ) ;
assign n31359 =  ( n30928 ) ? ( VREG_13_7 ) : ( n31358 ) ;
assign n31360 =  ( n30927 ) ? ( VREG_13_8 ) : ( n31359 ) ;
assign n31361 =  ( n30926 ) ? ( VREG_13_9 ) : ( n31360 ) ;
assign n31362 =  ( n30925 ) ? ( VREG_13_10 ) : ( n31361 ) ;
assign n31363 =  ( n30924 ) ? ( VREG_13_11 ) : ( n31362 ) ;
assign n31364 =  ( n30923 ) ? ( VREG_13_12 ) : ( n31363 ) ;
assign n31365 =  ( n30922 ) ? ( VREG_13_13 ) : ( n31364 ) ;
assign n31366 =  ( n30921 ) ? ( VREG_13_14 ) : ( n31365 ) ;
assign n31367 =  ( n30920 ) ? ( VREG_13_15 ) : ( n31366 ) ;
assign n31368 =  ( n30919 ) ? ( VREG_14_0 ) : ( n31367 ) ;
assign n31369 =  ( n30918 ) ? ( VREG_14_1 ) : ( n31368 ) ;
assign n31370 =  ( n30917 ) ? ( VREG_14_2 ) : ( n31369 ) ;
assign n31371 =  ( n30916 ) ? ( VREG_14_3 ) : ( n31370 ) ;
assign n31372 =  ( n30915 ) ? ( VREG_14_4 ) : ( n31371 ) ;
assign n31373 =  ( n30914 ) ? ( VREG_14_5 ) : ( n31372 ) ;
assign n31374 =  ( n30913 ) ? ( VREG_14_6 ) : ( n31373 ) ;
assign n31375 =  ( n30912 ) ? ( VREG_14_7 ) : ( n31374 ) ;
assign n31376 =  ( n30911 ) ? ( VREG_14_8 ) : ( n31375 ) ;
assign n31377 =  ( n30910 ) ? ( VREG_14_9 ) : ( n31376 ) ;
assign n31378 =  ( n30909 ) ? ( VREG_14_10 ) : ( n31377 ) ;
assign n31379 =  ( n30908 ) ? ( VREG_14_11 ) : ( n31378 ) ;
assign n31380 =  ( n30907 ) ? ( VREG_14_12 ) : ( n31379 ) ;
assign n31381 =  ( n30906 ) ? ( VREG_14_13 ) : ( n31380 ) ;
assign n31382 =  ( n30905 ) ? ( VREG_14_14 ) : ( n31381 ) ;
assign n31383 =  ( n30904 ) ? ( VREG_14_15 ) : ( n31382 ) ;
assign n31384 =  ( n30903 ) ? ( VREG_15_0 ) : ( n31383 ) ;
assign n31385 =  ( n30902 ) ? ( VREG_15_1 ) : ( n31384 ) ;
assign n31386 =  ( n30901 ) ? ( VREG_15_2 ) : ( n31385 ) ;
assign n31387 =  ( n30900 ) ? ( VREG_15_3 ) : ( n31386 ) ;
assign n31388 =  ( n30899 ) ? ( VREG_15_4 ) : ( n31387 ) ;
assign n31389 =  ( n30898 ) ? ( VREG_15_5 ) : ( n31388 ) ;
assign n31390 =  ( n30897 ) ? ( VREG_15_6 ) : ( n31389 ) ;
assign n31391 =  ( n30896 ) ? ( VREG_15_7 ) : ( n31390 ) ;
assign n31392 =  ( n30895 ) ? ( VREG_15_8 ) : ( n31391 ) ;
assign n31393 =  ( n30894 ) ? ( VREG_15_9 ) : ( n31392 ) ;
assign n31394 =  ( n30893 ) ? ( VREG_15_10 ) : ( n31393 ) ;
assign n31395 =  ( n30892 ) ? ( VREG_15_11 ) : ( n31394 ) ;
assign n31396 =  ( n30891 ) ? ( VREG_15_12 ) : ( n31395 ) ;
assign n31397 =  ( n30890 ) ? ( VREG_15_13 ) : ( n31396 ) ;
assign n31398 =  ( n30889 ) ? ( VREG_15_14 ) : ( n31397 ) ;
assign n31399 =  ( n30888 ) ? ( VREG_15_15 ) : ( n31398 ) ;
assign n31400 =  ( n30887 ) ? ( VREG_16_0 ) : ( n31399 ) ;
assign n31401 =  ( n30886 ) ? ( VREG_16_1 ) : ( n31400 ) ;
assign n31402 =  ( n30885 ) ? ( VREG_16_2 ) : ( n31401 ) ;
assign n31403 =  ( n30884 ) ? ( VREG_16_3 ) : ( n31402 ) ;
assign n31404 =  ( n30883 ) ? ( VREG_16_4 ) : ( n31403 ) ;
assign n31405 =  ( n30882 ) ? ( VREG_16_5 ) : ( n31404 ) ;
assign n31406 =  ( n30881 ) ? ( VREG_16_6 ) : ( n31405 ) ;
assign n31407 =  ( n30880 ) ? ( VREG_16_7 ) : ( n31406 ) ;
assign n31408 =  ( n30879 ) ? ( VREG_16_8 ) : ( n31407 ) ;
assign n31409 =  ( n30878 ) ? ( VREG_16_9 ) : ( n31408 ) ;
assign n31410 =  ( n30877 ) ? ( VREG_16_10 ) : ( n31409 ) ;
assign n31411 =  ( n30876 ) ? ( VREG_16_11 ) : ( n31410 ) ;
assign n31412 =  ( n30875 ) ? ( VREG_16_12 ) : ( n31411 ) ;
assign n31413 =  ( n30874 ) ? ( VREG_16_13 ) : ( n31412 ) ;
assign n31414 =  ( n30873 ) ? ( VREG_16_14 ) : ( n31413 ) ;
assign n31415 =  ( n30872 ) ? ( VREG_16_15 ) : ( n31414 ) ;
assign n31416 =  ( n30871 ) ? ( VREG_17_0 ) : ( n31415 ) ;
assign n31417 =  ( n30870 ) ? ( VREG_17_1 ) : ( n31416 ) ;
assign n31418 =  ( n30869 ) ? ( VREG_17_2 ) : ( n31417 ) ;
assign n31419 =  ( n30868 ) ? ( VREG_17_3 ) : ( n31418 ) ;
assign n31420 =  ( n30867 ) ? ( VREG_17_4 ) : ( n31419 ) ;
assign n31421 =  ( n30866 ) ? ( VREG_17_5 ) : ( n31420 ) ;
assign n31422 =  ( n30865 ) ? ( VREG_17_6 ) : ( n31421 ) ;
assign n31423 =  ( n30864 ) ? ( VREG_17_7 ) : ( n31422 ) ;
assign n31424 =  ( n30863 ) ? ( VREG_17_8 ) : ( n31423 ) ;
assign n31425 =  ( n30862 ) ? ( VREG_17_9 ) : ( n31424 ) ;
assign n31426 =  ( n30861 ) ? ( VREG_17_10 ) : ( n31425 ) ;
assign n31427 =  ( n30860 ) ? ( VREG_17_11 ) : ( n31426 ) ;
assign n31428 =  ( n30859 ) ? ( VREG_17_12 ) : ( n31427 ) ;
assign n31429 =  ( n30858 ) ? ( VREG_17_13 ) : ( n31428 ) ;
assign n31430 =  ( n30857 ) ? ( VREG_17_14 ) : ( n31429 ) ;
assign n31431 =  ( n30856 ) ? ( VREG_17_15 ) : ( n31430 ) ;
assign n31432 =  ( n30855 ) ? ( VREG_18_0 ) : ( n31431 ) ;
assign n31433 =  ( n30854 ) ? ( VREG_18_1 ) : ( n31432 ) ;
assign n31434 =  ( n30853 ) ? ( VREG_18_2 ) : ( n31433 ) ;
assign n31435 =  ( n30852 ) ? ( VREG_18_3 ) : ( n31434 ) ;
assign n31436 =  ( n30851 ) ? ( VREG_18_4 ) : ( n31435 ) ;
assign n31437 =  ( n30850 ) ? ( VREG_18_5 ) : ( n31436 ) ;
assign n31438 =  ( n30849 ) ? ( VREG_18_6 ) : ( n31437 ) ;
assign n31439 =  ( n30848 ) ? ( VREG_18_7 ) : ( n31438 ) ;
assign n31440 =  ( n30847 ) ? ( VREG_18_8 ) : ( n31439 ) ;
assign n31441 =  ( n30846 ) ? ( VREG_18_9 ) : ( n31440 ) ;
assign n31442 =  ( n30845 ) ? ( VREG_18_10 ) : ( n31441 ) ;
assign n31443 =  ( n30844 ) ? ( VREG_18_11 ) : ( n31442 ) ;
assign n31444 =  ( n30843 ) ? ( VREG_18_12 ) : ( n31443 ) ;
assign n31445 =  ( n30842 ) ? ( VREG_18_13 ) : ( n31444 ) ;
assign n31446 =  ( n30841 ) ? ( VREG_18_14 ) : ( n31445 ) ;
assign n31447 =  ( n30840 ) ? ( VREG_18_15 ) : ( n31446 ) ;
assign n31448 =  ( n30839 ) ? ( VREG_19_0 ) : ( n31447 ) ;
assign n31449 =  ( n30838 ) ? ( VREG_19_1 ) : ( n31448 ) ;
assign n31450 =  ( n30837 ) ? ( VREG_19_2 ) : ( n31449 ) ;
assign n31451 =  ( n30836 ) ? ( VREG_19_3 ) : ( n31450 ) ;
assign n31452 =  ( n30835 ) ? ( VREG_19_4 ) : ( n31451 ) ;
assign n31453 =  ( n30834 ) ? ( VREG_19_5 ) : ( n31452 ) ;
assign n31454 =  ( n30833 ) ? ( VREG_19_6 ) : ( n31453 ) ;
assign n31455 =  ( n30832 ) ? ( VREG_19_7 ) : ( n31454 ) ;
assign n31456 =  ( n30831 ) ? ( VREG_19_8 ) : ( n31455 ) ;
assign n31457 =  ( n30830 ) ? ( VREG_19_9 ) : ( n31456 ) ;
assign n31458 =  ( n30829 ) ? ( VREG_19_10 ) : ( n31457 ) ;
assign n31459 =  ( n30828 ) ? ( VREG_19_11 ) : ( n31458 ) ;
assign n31460 =  ( n30827 ) ? ( VREG_19_12 ) : ( n31459 ) ;
assign n31461 =  ( n30826 ) ? ( VREG_19_13 ) : ( n31460 ) ;
assign n31462 =  ( n30825 ) ? ( VREG_19_14 ) : ( n31461 ) ;
assign n31463 =  ( n30824 ) ? ( VREG_19_15 ) : ( n31462 ) ;
assign n31464 =  ( n30823 ) ? ( VREG_20_0 ) : ( n31463 ) ;
assign n31465 =  ( n30822 ) ? ( VREG_20_1 ) : ( n31464 ) ;
assign n31466 =  ( n30821 ) ? ( VREG_20_2 ) : ( n31465 ) ;
assign n31467 =  ( n30820 ) ? ( VREG_20_3 ) : ( n31466 ) ;
assign n31468 =  ( n30819 ) ? ( VREG_20_4 ) : ( n31467 ) ;
assign n31469 =  ( n30818 ) ? ( VREG_20_5 ) : ( n31468 ) ;
assign n31470 =  ( n30817 ) ? ( VREG_20_6 ) : ( n31469 ) ;
assign n31471 =  ( n30816 ) ? ( VREG_20_7 ) : ( n31470 ) ;
assign n31472 =  ( n30815 ) ? ( VREG_20_8 ) : ( n31471 ) ;
assign n31473 =  ( n30814 ) ? ( VREG_20_9 ) : ( n31472 ) ;
assign n31474 =  ( n30813 ) ? ( VREG_20_10 ) : ( n31473 ) ;
assign n31475 =  ( n30812 ) ? ( VREG_20_11 ) : ( n31474 ) ;
assign n31476 =  ( n30811 ) ? ( VREG_20_12 ) : ( n31475 ) ;
assign n31477 =  ( n30810 ) ? ( VREG_20_13 ) : ( n31476 ) ;
assign n31478 =  ( n30809 ) ? ( VREG_20_14 ) : ( n31477 ) ;
assign n31479 =  ( n30808 ) ? ( VREG_20_15 ) : ( n31478 ) ;
assign n31480 =  ( n30807 ) ? ( VREG_21_0 ) : ( n31479 ) ;
assign n31481 =  ( n30806 ) ? ( VREG_21_1 ) : ( n31480 ) ;
assign n31482 =  ( n30805 ) ? ( VREG_21_2 ) : ( n31481 ) ;
assign n31483 =  ( n30804 ) ? ( VREG_21_3 ) : ( n31482 ) ;
assign n31484 =  ( n30803 ) ? ( VREG_21_4 ) : ( n31483 ) ;
assign n31485 =  ( n30802 ) ? ( VREG_21_5 ) : ( n31484 ) ;
assign n31486 =  ( n30801 ) ? ( VREG_21_6 ) : ( n31485 ) ;
assign n31487 =  ( n30800 ) ? ( VREG_21_7 ) : ( n31486 ) ;
assign n31488 =  ( n30799 ) ? ( VREG_21_8 ) : ( n31487 ) ;
assign n31489 =  ( n30798 ) ? ( VREG_21_9 ) : ( n31488 ) ;
assign n31490 =  ( n30797 ) ? ( VREG_21_10 ) : ( n31489 ) ;
assign n31491 =  ( n30796 ) ? ( VREG_21_11 ) : ( n31490 ) ;
assign n31492 =  ( n30795 ) ? ( VREG_21_12 ) : ( n31491 ) ;
assign n31493 =  ( n30794 ) ? ( VREG_21_13 ) : ( n31492 ) ;
assign n31494 =  ( n30793 ) ? ( VREG_21_14 ) : ( n31493 ) ;
assign n31495 =  ( n30792 ) ? ( VREG_21_15 ) : ( n31494 ) ;
assign n31496 =  ( n30791 ) ? ( VREG_22_0 ) : ( n31495 ) ;
assign n31497 =  ( n30790 ) ? ( VREG_22_1 ) : ( n31496 ) ;
assign n31498 =  ( n30789 ) ? ( VREG_22_2 ) : ( n31497 ) ;
assign n31499 =  ( n30788 ) ? ( VREG_22_3 ) : ( n31498 ) ;
assign n31500 =  ( n30787 ) ? ( VREG_22_4 ) : ( n31499 ) ;
assign n31501 =  ( n30786 ) ? ( VREG_22_5 ) : ( n31500 ) ;
assign n31502 =  ( n30785 ) ? ( VREG_22_6 ) : ( n31501 ) ;
assign n31503 =  ( n30784 ) ? ( VREG_22_7 ) : ( n31502 ) ;
assign n31504 =  ( n30783 ) ? ( VREG_22_8 ) : ( n31503 ) ;
assign n31505 =  ( n30782 ) ? ( VREG_22_9 ) : ( n31504 ) ;
assign n31506 =  ( n30781 ) ? ( VREG_22_10 ) : ( n31505 ) ;
assign n31507 =  ( n30780 ) ? ( VREG_22_11 ) : ( n31506 ) ;
assign n31508 =  ( n30779 ) ? ( VREG_22_12 ) : ( n31507 ) ;
assign n31509 =  ( n30778 ) ? ( VREG_22_13 ) : ( n31508 ) ;
assign n31510 =  ( n30777 ) ? ( VREG_22_14 ) : ( n31509 ) ;
assign n31511 =  ( n30776 ) ? ( VREG_22_15 ) : ( n31510 ) ;
assign n31512 =  ( n30775 ) ? ( VREG_23_0 ) : ( n31511 ) ;
assign n31513 =  ( n30774 ) ? ( VREG_23_1 ) : ( n31512 ) ;
assign n31514 =  ( n30773 ) ? ( VREG_23_2 ) : ( n31513 ) ;
assign n31515 =  ( n30772 ) ? ( VREG_23_3 ) : ( n31514 ) ;
assign n31516 =  ( n30771 ) ? ( VREG_23_4 ) : ( n31515 ) ;
assign n31517 =  ( n30770 ) ? ( VREG_23_5 ) : ( n31516 ) ;
assign n31518 =  ( n30769 ) ? ( VREG_23_6 ) : ( n31517 ) ;
assign n31519 =  ( n30768 ) ? ( VREG_23_7 ) : ( n31518 ) ;
assign n31520 =  ( n30767 ) ? ( VREG_23_8 ) : ( n31519 ) ;
assign n31521 =  ( n30766 ) ? ( VREG_23_9 ) : ( n31520 ) ;
assign n31522 =  ( n30765 ) ? ( VREG_23_10 ) : ( n31521 ) ;
assign n31523 =  ( n30764 ) ? ( VREG_23_11 ) : ( n31522 ) ;
assign n31524 =  ( n30763 ) ? ( VREG_23_12 ) : ( n31523 ) ;
assign n31525 =  ( n30762 ) ? ( VREG_23_13 ) : ( n31524 ) ;
assign n31526 =  ( n30761 ) ? ( VREG_23_14 ) : ( n31525 ) ;
assign n31527 =  ( n30760 ) ? ( VREG_23_15 ) : ( n31526 ) ;
assign n31528 =  ( n30759 ) ? ( VREG_24_0 ) : ( n31527 ) ;
assign n31529 =  ( n30758 ) ? ( VREG_24_1 ) : ( n31528 ) ;
assign n31530 =  ( n30757 ) ? ( VREG_24_2 ) : ( n31529 ) ;
assign n31531 =  ( n30756 ) ? ( VREG_24_3 ) : ( n31530 ) ;
assign n31532 =  ( n30755 ) ? ( VREG_24_4 ) : ( n31531 ) ;
assign n31533 =  ( n30754 ) ? ( VREG_24_5 ) : ( n31532 ) ;
assign n31534 =  ( n30753 ) ? ( VREG_24_6 ) : ( n31533 ) ;
assign n31535 =  ( n30752 ) ? ( VREG_24_7 ) : ( n31534 ) ;
assign n31536 =  ( n30751 ) ? ( VREG_24_8 ) : ( n31535 ) ;
assign n31537 =  ( n30750 ) ? ( VREG_24_9 ) : ( n31536 ) ;
assign n31538 =  ( n30749 ) ? ( VREG_24_10 ) : ( n31537 ) ;
assign n31539 =  ( n30748 ) ? ( VREG_24_11 ) : ( n31538 ) ;
assign n31540 =  ( n30747 ) ? ( VREG_24_12 ) : ( n31539 ) ;
assign n31541 =  ( n30746 ) ? ( VREG_24_13 ) : ( n31540 ) ;
assign n31542 =  ( n30745 ) ? ( VREG_24_14 ) : ( n31541 ) ;
assign n31543 =  ( n30744 ) ? ( VREG_24_15 ) : ( n31542 ) ;
assign n31544 =  ( n30743 ) ? ( VREG_25_0 ) : ( n31543 ) ;
assign n31545 =  ( n30742 ) ? ( VREG_25_1 ) : ( n31544 ) ;
assign n31546 =  ( n30741 ) ? ( VREG_25_2 ) : ( n31545 ) ;
assign n31547 =  ( n30740 ) ? ( VREG_25_3 ) : ( n31546 ) ;
assign n31548 =  ( n30739 ) ? ( VREG_25_4 ) : ( n31547 ) ;
assign n31549 =  ( n30738 ) ? ( VREG_25_5 ) : ( n31548 ) ;
assign n31550 =  ( n30737 ) ? ( VREG_25_6 ) : ( n31549 ) ;
assign n31551 =  ( n30736 ) ? ( VREG_25_7 ) : ( n31550 ) ;
assign n31552 =  ( n30735 ) ? ( VREG_25_8 ) : ( n31551 ) ;
assign n31553 =  ( n30734 ) ? ( VREG_25_9 ) : ( n31552 ) ;
assign n31554 =  ( n30733 ) ? ( VREG_25_10 ) : ( n31553 ) ;
assign n31555 =  ( n30732 ) ? ( VREG_25_11 ) : ( n31554 ) ;
assign n31556 =  ( n30731 ) ? ( VREG_25_12 ) : ( n31555 ) ;
assign n31557 =  ( n30730 ) ? ( VREG_25_13 ) : ( n31556 ) ;
assign n31558 =  ( n30729 ) ? ( VREG_25_14 ) : ( n31557 ) ;
assign n31559 =  ( n30728 ) ? ( VREG_25_15 ) : ( n31558 ) ;
assign n31560 =  ( n30727 ) ? ( VREG_26_0 ) : ( n31559 ) ;
assign n31561 =  ( n30726 ) ? ( VREG_26_1 ) : ( n31560 ) ;
assign n31562 =  ( n30725 ) ? ( VREG_26_2 ) : ( n31561 ) ;
assign n31563 =  ( n30724 ) ? ( VREG_26_3 ) : ( n31562 ) ;
assign n31564 =  ( n30723 ) ? ( VREG_26_4 ) : ( n31563 ) ;
assign n31565 =  ( n30722 ) ? ( VREG_26_5 ) : ( n31564 ) ;
assign n31566 =  ( n30721 ) ? ( VREG_26_6 ) : ( n31565 ) ;
assign n31567 =  ( n30720 ) ? ( VREG_26_7 ) : ( n31566 ) ;
assign n31568 =  ( n30719 ) ? ( VREG_26_8 ) : ( n31567 ) ;
assign n31569 =  ( n30718 ) ? ( VREG_26_9 ) : ( n31568 ) ;
assign n31570 =  ( n30717 ) ? ( VREG_26_10 ) : ( n31569 ) ;
assign n31571 =  ( n30716 ) ? ( VREG_26_11 ) : ( n31570 ) ;
assign n31572 =  ( n30715 ) ? ( VREG_26_12 ) : ( n31571 ) ;
assign n31573 =  ( n30714 ) ? ( VREG_26_13 ) : ( n31572 ) ;
assign n31574 =  ( n30713 ) ? ( VREG_26_14 ) : ( n31573 ) ;
assign n31575 =  ( n30712 ) ? ( VREG_26_15 ) : ( n31574 ) ;
assign n31576 =  ( n30711 ) ? ( VREG_27_0 ) : ( n31575 ) ;
assign n31577 =  ( n30710 ) ? ( VREG_27_1 ) : ( n31576 ) ;
assign n31578 =  ( n30709 ) ? ( VREG_27_2 ) : ( n31577 ) ;
assign n31579 =  ( n30708 ) ? ( VREG_27_3 ) : ( n31578 ) ;
assign n31580 =  ( n30707 ) ? ( VREG_27_4 ) : ( n31579 ) ;
assign n31581 =  ( n30706 ) ? ( VREG_27_5 ) : ( n31580 ) ;
assign n31582 =  ( n30705 ) ? ( VREG_27_6 ) : ( n31581 ) ;
assign n31583 =  ( n30704 ) ? ( VREG_27_7 ) : ( n31582 ) ;
assign n31584 =  ( n30703 ) ? ( VREG_27_8 ) : ( n31583 ) ;
assign n31585 =  ( n30702 ) ? ( VREG_27_9 ) : ( n31584 ) ;
assign n31586 =  ( n30701 ) ? ( VREG_27_10 ) : ( n31585 ) ;
assign n31587 =  ( n30700 ) ? ( VREG_27_11 ) : ( n31586 ) ;
assign n31588 =  ( n30699 ) ? ( VREG_27_12 ) : ( n31587 ) ;
assign n31589 =  ( n30698 ) ? ( VREG_27_13 ) : ( n31588 ) ;
assign n31590 =  ( n30697 ) ? ( VREG_27_14 ) : ( n31589 ) ;
assign n31591 =  ( n30696 ) ? ( VREG_27_15 ) : ( n31590 ) ;
assign n31592 =  ( n30695 ) ? ( VREG_28_0 ) : ( n31591 ) ;
assign n31593 =  ( n30694 ) ? ( VREG_28_1 ) : ( n31592 ) ;
assign n31594 =  ( n30693 ) ? ( VREG_28_2 ) : ( n31593 ) ;
assign n31595 =  ( n30692 ) ? ( VREG_28_3 ) : ( n31594 ) ;
assign n31596 =  ( n30691 ) ? ( VREG_28_4 ) : ( n31595 ) ;
assign n31597 =  ( n30690 ) ? ( VREG_28_5 ) : ( n31596 ) ;
assign n31598 =  ( n30689 ) ? ( VREG_28_6 ) : ( n31597 ) ;
assign n31599 =  ( n30688 ) ? ( VREG_28_7 ) : ( n31598 ) ;
assign n31600 =  ( n30687 ) ? ( VREG_28_8 ) : ( n31599 ) ;
assign n31601 =  ( n30686 ) ? ( VREG_28_9 ) : ( n31600 ) ;
assign n31602 =  ( n30685 ) ? ( VREG_28_10 ) : ( n31601 ) ;
assign n31603 =  ( n30684 ) ? ( VREG_28_11 ) : ( n31602 ) ;
assign n31604 =  ( n30683 ) ? ( VREG_28_12 ) : ( n31603 ) ;
assign n31605 =  ( n30682 ) ? ( VREG_28_13 ) : ( n31604 ) ;
assign n31606 =  ( n30681 ) ? ( VREG_28_14 ) : ( n31605 ) ;
assign n31607 =  ( n30680 ) ? ( VREG_28_15 ) : ( n31606 ) ;
assign n31608 =  ( n30679 ) ? ( VREG_29_0 ) : ( n31607 ) ;
assign n31609 =  ( n30678 ) ? ( VREG_29_1 ) : ( n31608 ) ;
assign n31610 =  ( n30677 ) ? ( VREG_29_2 ) : ( n31609 ) ;
assign n31611 =  ( n30676 ) ? ( VREG_29_3 ) : ( n31610 ) ;
assign n31612 =  ( n30675 ) ? ( VREG_29_4 ) : ( n31611 ) ;
assign n31613 =  ( n30674 ) ? ( VREG_29_5 ) : ( n31612 ) ;
assign n31614 =  ( n30673 ) ? ( VREG_29_6 ) : ( n31613 ) ;
assign n31615 =  ( n30672 ) ? ( VREG_29_7 ) : ( n31614 ) ;
assign n31616 =  ( n30671 ) ? ( VREG_29_8 ) : ( n31615 ) ;
assign n31617 =  ( n30670 ) ? ( VREG_29_9 ) : ( n31616 ) ;
assign n31618 =  ( n30669 ) ? ( VREG_29_10 ) : ( n31617 ) ;
assign n31619 =  ( n30668 ) ? ( VREG_29_11 ) : ( n31618 ) ;
assign n31620 =  ( n30667 ) ? ( VREG_29_12 ) : ( n31619 ) ;
assign n31621 =  ( n30666 ) ? ( VREG_29_13 ) : ( n31620 ) ;
assign n31622 =  ( n30665 ) ? ( VREG_29_14 ) : ( n31621 ) ;
assign n31623 =  ( n30664 ) ? ( VREG_29_15 ) : ( n31622 ) ;
assign n31624 =  ( n30663 ) ? ( VREG_30_0 ) : ( n31623 ) ;
assign n31625 =  ( n30662 ) ? ( VREG_30_1 ) : ( n31624 ) ;
assign n31626 =  ( n30661 ) ? ( VREG_30_2 ) : ( n31625 ) ;
assign n31627 =  ( n30660 ) ? ( VREG_30_3 ) : ( n31626 ) ;
assign n31628 =  ( n30659 ) ? ( VREG_30_4 ) : ( n31627 ) ;
assign n31629 =  ( n30658 ) ? ( VREG_30_5 ) : ( n31628 ) ;
assign n31630 =  ( n30657 ) ? ( VREG_30_6 ) : ( n31629 ) ;
assign n31631 =  ( n30656 ) ? ( VREG_30_7 ) : ( n31630 ) ;
assign n31632 =  ( n30655 ) ? ( VREG_30_8 ) : ( n31631 ) ;
assign n31633 =  ( n30654 ) ? ( VREG_30_9 ) : ( n31632 ) ;
assign n31634 =  ( n30653 ) ? ( VREG_30_10 ) : ( n31633 ) ;
assign n31635 =  ( n30652 ) ? ( VREG_30_11 ) : ( n31634 ) ;
assign n31636 =  ( n30651 ) ? ( VREG_30_12 ) : ( n31635 ) ;
assign n31637 =  ( n30650 ) ? ( VREG_30_13 ) : ( n31636 ) ;
assign n31638 =  ( n30649 ) ? ( VREG_30_14 ) : ( n31637 ) ;
assign n31639 =  ( n30648 ) ? ( VREG_30_15 ) : ( n31638 ) ;
assign n31640 =  ( n30647 ) ? ( VREG_31_0 ) : ( n31639 ) ;
assign n31641 =  ( n30645 ) ? ( VREG_31_1 ) : ( n31640 ) ;
assign n31642 =  ( n30643 ) ? ( VREG_31_2 ) : ( n31641 ) ;
assign n31643 =  ( n30641 ) ? ( VREG_31_3 ) : ( n31642 ) ;
assign n31644 =  ( n30639 ) ? ( VREG_31_4 ) : ( n31643 ) ;
assign n31645 =  ( n30637 ) ? ( VREG_31_5 ) : ( n31644 ) ;
assign n31646 =  ( n30635 ) ? ( VREG_31_6 ) : ( n31645 ) ;
assign n31647 =  ( n30633 ) ? ( VREG_31_7 ) : ( n31646 ) ;
assign n31648 =  ( n30631 ) ? ( VREG_31_8 ) : ( n31647 ) ;
assign n31649 =  ( n30629 ) ? ( VREG_31_9 ) : ( n31648 ) ;
assign n31650 =  ( n30627 ) ? ( VREG_31_10 ) : ( n31649 ) ;
assign n31651 =  ( n30625 ) ? ( VREG_31_11 ) : ( n31650 ) ;
assign n31652 =  ( n30623 ) ? ( VREG_31_12 ) : ( n31651 ) ;
assign n31653 =  ( n30621 ) ? ( VREG_31_13 ) : ( n31652 ) ;
assign n31654 =  ( n30619 ) ? ( VREG_31_14 ) : ( n31653 ) ;
assign n31655 =  ( n30617 ) ? ( VREG_31_15 ) : ( n31654 ) ;
assign n31656 =  ( n31655 ) + ( n140 )  ;
assign n31657 =  ( n31655 ) - ( n140 )  ;
assign n31658 =  ( n31655 ) & ( n140 )  ;
assign n31659 =  ( n31655 ) | ( n140 )  ;
assign n31660 =  ( ( n31655 ) * ( n140 ))  ;
assign n31661 =  ( n148 ) ? ( n31660 ) : ( VREG_0_8 ) ;
assign n31662 =  ( n146 ) ? ( n31659 ) : ( n31661 ) ;
assign n31663 =  ( n144 ) ? ( n31658 ) : ( n31662 ) ;
assign n31664 =  ( n142 ) ? ( n31657 ) : ( n31663 ) ;
assign n31665 =  ( n10 ) ? ( n31656 ) : ( n31664 ) ;
assign n31666 =  ( n77 ) & ( n30616 )  ;
assign n31667 =  ( n77 ) & ( n30618 )  ;
assign n31668 =  ( n77 ) & ( n30620 )  ;
assign n31669 =  ( n77 ) & ( n30622 )  ;
assign n31670 =  ( n77 ) & ( n30624 )  ;
assign n31671 =  ( n77 ) & ( n30626 )  ;
assign n31672 =  ( n77 ) & ( n30628 )  ;
assign n31673 =  ( n77 ) & ( n30630 )  ;
assign n31674 =  ( n77 ) & ( n30632 )  ;
assign n31675 =  ( n77 ) & ( n30634 )  ;
assign n31676 =  ( n77 ) & ( n30636 )  ;
assign n31677 =  ( n77 ) & ( n30638 )  ;
assign n31678 =  ( n77 ) & ( n30640 )  ;
assign n31679 =  ( n77 ) & ( n30642 )  ;
assign n31680 =  ( n77 ) & ( n30644 )  ;
assign n31681 =  ( n77 ) & ( n30646 )  ;
assign n31682 =  ( n78 ) & ( n30616 )  ;
assign n31683 =  ( n78 ) & ( n30618 )  ;
assign n31684 =  ( n78 ) & ( n30620 )  ;
assign n31685 =  ( n78 ) & ( n30622 )  ;
assign n31686 =  ( n78 ) & ( n30624 )  ;
assign n31687 =  ( n78 ) & ( n30626 )  ;
assign n31688 =  ( n78 ) & ( n30628 )  ;
assign n31689 =  ( n78 ) & ( n30630 )  ;
assign n31690 =  ( n78 ) & ( n30632 )  ;
assign n31691 =  ( n78 ) & ( n30634 )  ;
assign n31692 =  ( n78 ) & ( n30636 )  ;
assign n31693 =  ( n78 ) & ( n30638 )  ;
assign n31694 =  ( n78 ) & ( n30640 )  ;
assign n31695 =  ( n78 ) & ( n30642 )  ;
assign n31696 =  ( n78 ) & ( n30644 )  ;
assign n31697 =  ( n78 ) & ( n30646 )  ;
assign n31698 =  ( n79 ) & ( n30616 )  ;
assign n31699 =  ( n79 ) & ( n30618 )  ;
assign n31700 =  ( n79 ) & ( n30620 )  ;
assign n31701 =  ( n79 ) & ( n30622 )  ;
assign n31702 =  ( n79 ) & ( n30624 )  ;
assign n31703 =  ( n79 ) & ( n30626 )  ;
assign n31704 =  ( n79 ) & ( n30628 )  ;
assign n31705 =  ( n79 ) & ( n30630 )  ;
assign n31706 =  ( n79 ) & ( n30632 )  ;
assign n31707 =  ( n79 ) & ( n30634 )  ;
assign n31708 =  ( n79 ) & ( n30636 )  ;
assign n31709 =  ( n79 ) & ( n30638 )  ;
assign n31710 =  ( n79 ) & ( n30640 )  ;
assign n31711 =  ( n79 ) & ( n30642 )  ;
assign n31712 =  ( n79 ) & ( n30644 )  ;
assign n31713 =  ( n79 ) & ( n30646 )  ;
assign n31714 =  ( n80 ) & ( n30616 )  ;
assign n31715 =  ( n80 ) & ( n30618 )  ;
assign n31716 =  ( n80 ) & ( n30620 )  ;
assign n31717 =  ( n80 ) & ( n30622 )  ;
assign n31718 =  ( n80 ) & ( n30624 )  ;
assign n31719 =  ( n80 ) & ( n30626 )  ;
assign n31720 =  ( n80 ) & ( n30628 )  ;
assign n31721 =  ( n80 ) & ( n30630 )  ;
assign n31722 =  ( n80 ) & ( n30632 )  ;
assign n31723 =  ( n80 ) & ( n30634 )  ;
assign n31724 =  ( n80 ) & ( n30636 )  ;
assign n31725 =  ( n80 ) & ( n30638 )  ;
assign n31726 =  ( n80 ) & ( n30640 )  ;
assign n31727 =  ( n80 ) & ( n30642 )  ;
assign n31728 =  ( n80 ) & ( n30644 )  ;
assign n31729 =  ( n80 ) & ( n30646 )  ;
assign n31730 =  ( n81 ) & ( n30616 )  ;
assign n31731 =  ( n81 ) & ( n30618 )  ;
assign n31732 =  ( n81 ) & ( n30620 )  ;
assign n31733 =  ( n81 ) & ( n30622 )  ;
assign n31734 =  ( n81 ) & ( n30624 )  ;
assign n31735 =  ( n81 ) & ( n30626 )  ;
assign n31736 =  ( n81 ) & ( n30628 )  ;
assign n31737 =  ( n81 ) & ( n30630 )  ;
assign n31738 =  ( n81 ) & ( n30632 )  ;
assign n31739 =  ( n81 ) & ( n30634 )  ;
assign n31740 =  ( n81 ) & ( n30636 )  ;
assign n31741 =  ( n81 ) & ( n30638 )  ;
assign n31742 =  ( n81 ) & ( n30640 )  ;
assign n31743 =  ( n81 ) & ( n30642 )  ;
assign n31744 =  ( n81 ) & ( n30644 )  ;
assign n31745 =  ( n81 ) & ( n30646 )  ;
assign n31746 =  ( n82 ) & ( n30616 )  ;
assign n31747 =  ( n82 ) & ( n30618 )  ;
assign n31748 =  ( n82 ) & ( n30620 )  ;
assign n31749 =  ( n82 ) & ( n30622 )  ;
assign n31750 =  ( n82 ) & ( n30624 )  ;
assign n31751 =  ( n82 ) & ( n30626 )  ;
assign n31752 =  ( n82 ) & ( n30628 )  ;
assign n31753 =  ( n82 ) & ( n30630 )  ;
assign n31754 =  ( n82 ) & ( n30632 )  ;
assign n31755 =  ( n82 ) & ( n30634 )  ;
assign n31756 =  ( n82 ) & ( n30636 )  ;
assign n31757 =  ( n82 ) & ( n30638 )  ;
assign n31758 =  ( n82 ) & ( n30640 )  ;
assign n31759 =  ( n82 ) & ( n30642 )  ;
assign n31760 =  ( n82 ) & ( n30644 )  ;
assign n31761 =  ( n82 ) & ( n30646 )  ;
assign n31762 =  ( n83 ) & ( n30616 )  ;
assign n31763 =  ( n83 ) & ( n30618 )  ;
assign n31764 =  ( n83 ) & ( n30620 )  ;
assign n31765 =  ( n83 ) & ( n30622 )  ;
assign n31766 =  ( n83 ) & ( n30624 )  ;
assign n31767 =  ( n83 ) & ( n30626 )  ;
assign n31768 =  ( n83 ) & ( n30628 )  ;
assign n31769 =  ( n83 ) & ( n30630 )  ;
assign n31770 =  ( n83 ) & ( n30632 )  ;
assign n31771 =  ( n83 ) & ( n30634 )  ;
assign n31772 =  ( n83 ) & ( n30636 )  ;
assign n31773 =  ( n83 ) & ( n30638 )  ;
assign n31774 =  ( n83 ) & ( n30640 )  ;
assign n31775 =  ( n83 ) & ( n30642 )  ;
assign n31776 =  ( n83 ) & ( n30644 )  ;
assign n31777 =  ( n83 ) & ( n30646 )  ;
assign n31778 =  ( n84 ) & ( n30616 )  ;
assign n31779 =  ( n84 ) & ( n30618 )  ;
assign n31780 =  ( n84 ) & ( n30620 )  ;
assign n31781 =  ( n84 ) & ( n30622 )  ;
assign n31782 =  ( n84 ) & ( n30624 )  ;
assign n31783 =  ( n84 ) & ( n30626 )  ;
assign n31784 =  ( n84 ) & ( n30628 )  ;
assign n31785 =  ( n84 ) & ( n30630 )  ;
assign n31786 =  ( n84 ) & ( n30632 )  ;
assign n31787 =  ( n84 ) & ( n30634 )  ;
assign n31788 =  ( n84 ) & ( n30636 )  ;
assign n31789 =  ( n84 ) & ( n30638 )  ;
assign n31790 =  ( n84 ) & ( n30640 )  ;
assign n31791 =  ( n84 ) & ( n30642 )  ;
assign n31792 =  ( n84 ) & ( n30644 )  ;
assign n31793 =  ( n84 ) & ( n30646 )  ;
assign n31794 =  ( n85 ) & ( n30616 )  ;
assign n31795 =  ( n85 ) & ( n30618 )  ;
assign n31796 =  ( n85 ) & ( n30620 )  ;
assign n31797 =  ( n85 ) & ( n30622 )  ;
assign n31798 =  ( n85 ) & ( n30624 )  ;
assign n31799 =  ( n85 ) & ( n30626 )  ;
assign n31800 =  ( n85 ) & ( n30628 )  ;
assign n31801 =  ( n85 ) & ( n30630 )  ;
assign n31802 =  ( n85 ) & ( n30632 )  ;
assign n31803 =  ( n85 ) & ( n30634 )  ;
assign n31804 =  ( n85 ) & ( n30636 )  ;
assign n31805 =  ( n85 ) & ( n30638 )  ;
assign n31806 =  ( n85 ) & ( n30640 )  ;
assign n31807 =  ( n85 ) & ( n30642 )  ;
assign n31808 =  ( n85 ) & ( n30644 )  ;
assign n31809 =  ( n85 ) & ( n30646 )  ;
assign n31810 =  ( n86 ) & ( n30616 )  ;
assign n31811 =  ( n86 ) & ( n30618 )  ;
assign n31812 =  ( n86 ) & ( n30620 )  ;
assign n31813 =  ( n86 ) & ( n30622 )  ;
assign n31814 =  ( n86 ) & ( n30624 )  ;
assign n31815 =  ( n86 ) & ( n30626 )  ;
assign n31816 =  ( n86 ) & ( n30628 )  ;
assign n31817 =  ( n86 ) & ( n30630 )  ;
assign n31818 =  ( n86 ) & ( n30632 )  ;
assign n31819 =  ( n86 ) & ( n30634 )  ;
assign n31820 =  ( n86 ) & ( n30636 )  ;
assign n31821 =  ( n86 ) & ( n30638 )  ;
assign n31822 =  ( n86 ) & ( n30640 )  ;
assign n31823 =  ( n86 ) & ( n30642 )  ;
assign n31824 =  ( n86 ) & ( n30644 )  ;
assign n31825 =  ( n86 ) & ( n30646 )  ;
assign n31826 =  ( n87 ) & ( n30616 )  ;
assign n31827 =  ( n87 ) & ( n30618 )  ;
assign n31828 =  ( n87 ) & ( n30620 )  ;
assign n31829 =  ( n87 ) & ( n30622 )  ;
assign n31830 =  ( n87 ) & ( n30624 )  ;
assign n31831 =  ( n87 ) & ( n30626 )  ;
assign n31832 =  ( n87 ) & ( n30628 )  ;
assign n31833 =  ( n87 ) & ( n30630 )  ;
assign n31834 =  ( n87 ) & ( n30632 )  ;
assign n31835 =  ( n87 ) & ( n30634 )  ;
assign n31836 =  ( n87 ) & ( n30636 )  ;
assign n31837 =  ( n87 ) & ( n30638 )  ;
assign n31838 =  ( n87 ) & ( n30640 )  ;
assign n31839 =  ( n87 ) & ( n30642 )  ;
assign n31840 =  ( n87 ) & ( n30644 )  ;
assign n31841 =  ( n87 ) & ( n30646 )  ;
assign n31842 =  ( n88 ) & ( n30616 )  ;
assign n31843 =  ( n88 ) & ( n30618 )  ;
assign n31844 =  ( n88 ) & ( n30620 )  ;
assign n31845 =  ( n88 ) & ( n30622 )  ;
assign n31846 =  ( n88 ) & ( n30624 )  ;
assign n31847 =  ( n88 ) & ( n30626 )  ;
assign n31848 =  ( n88 ) & ( n30628 )  ;
assign n31849 =  ( n88 ) & ( n30630 )  ;
assign n31850 =  ( n88 ) & ( n30632 )  ;
assign n31851 =  ( n88 ) & ( n30634 )  ;
assign n31852 =  ( n88 ) & ( n30636 )  ;
assign n31853 =  ( n88 ) & ( n30638 )  ;
assign n31854 =  ( n88 ) & ( n30640 )  ;
assign n31855 =  ( n88 ) & ( n30642 )  ;
assign n31856 =  ( n88 ) & ( n30644 )  ;
assign n31857 =  ( n88 ) & ( n30646 )  ;
assign n31858 =  ( n89 ) & ( n30616 )  ;
assign n31859 =  ( n89 ) & ( n30618 )  ;
assign n31860 =  ( n89 ) & ( n30620 )  ;
assign n31861 =  ( n89 ) & ( n30622 )  ;
assign n31862 =  ( n89 ) & ( n30624 )  ;
assign n31863 =  ( n89 ) & ( n30626 )  ;
assign n31864 =  ( n89 ) & ( n30628 )  ;
assign n31865 =  ( n89 ) & ( n30630 )  ;
assign n31866 =  ( n89 ) & ( n30632 )  ;
assign n31867 =  ( n89 ) & ( n30634 )  ;
assign n31868 =  ( n89 ) & ( n30636 )  ;
assign n31869 =  ( n89 ) & ( n30638 )  ;
assign n31870 =  ( n89 ) & ( n30640 )  ;
assign n31871 =  ( n89 ) & ( n30642 )  ;
assign n31872 =  ( n89 ) & ( n30644 )  ;
assign n31873 =  ( n89 ) & ( n30646 )  ;
assign n31874 =  ( n90 ) & ( n30616 )  ;
assign n31875 =  ( n90 ) & ( n30618 )  ;
assign n31876 =  ( n90 ) & ( n30620 )  ;
assign n31877 =  ( n90 ) & ( n30622 )  ;
assign n31878 =  ( n90 ) & ( n30624 )  ;
assign n31879 =  ( n90 ) & ( n30626 )  ;
assign n31880 =  ( n90 ) & ( n30628 )  ;
assign n31881 =  ( n90 ) & ( n30630 )  ;
assign n31882 =  ( n90 ) & ( n30632 )  ;
assign n31883 =  ( n90 ) & ( n30634 )  ;
assign n31884 =  ( n90 ) & ( n30636 )  ;
assign n31885 =  ( n90 ) & ( n30638 )  ;
assign n31886 =  ( n90 ) & ( n30640 )  ;
assign n31887 =  ( n90 ) & ( n30642 )  ;
assign n31888 =  ( n90 ) & ( n30644 )  ;
assign n31889 =  ( n90 ) & ( n30646 )  ;
assign n31890 =  ( n91 ) & ( n30616 )  ;
assign n31891 =  ( n91 ) & ( n30618 )  ;
assign n31892 =  ( n91 ) & ( n30620 )  ;
assign n31893 =  ( n91 ) & ( n30622 )  ;
assign n31894 =  ( n91 ) & ( n30624 )  ;
assign n31895 =  ( n91 ) & ( n30626 )  ;
assign n31896 =  ( n91 ) & ( n30628 )  ;
assign n31897 =  ( n91 ) & ( n30630 )  ;
assign n31898 =  ( n91 ) & ( n30632 )  ;
assign n31899 =  ( n91 ) & ( n30634 )  ;
assign n31900 =  ( n91 ) & ( n30636 )  ;
assign n31901 =  ( n91 ) & ( n30638 )  ;
assign n31902 =  ( n91 ) & ( n30640 )  ;
assign n31903 =  ( n91 ) & ( n30642 )  ;
assign n31904 =  ( n91 ) & ( n30644 )  ;
assign n31905 =  ( n91 ) & ( n30646 )  ;
assign n31906 =  ( n92 ) & ( n30616 )  ;
assign n31907 =  ( n92 ) & ( n30618 )  ;
assign n31908 =  ( n92 ) & ( n30620 )  ;
assign n31909 =  ( n92 ) & ( n30622 )  ;
assign n31910 =  ( n92 ) & ( n30624 )  ;
assign n31911 =  ( n92 ) & ( n30626 )  ;
assign n31912 =  ( n92 ) & ( n30628 )  ;
assign n31913 =  ( n92 ) & ( n30630 )  ;
assign n31914 =  ( n92 ) & ( n30632 )  ;
assign n31915 =  ( n92 ) & ( n30634 )  ;
assign n31916 =  ( n92 ) & ( n30636 )  ;
assign n31917 =  ( n92 ) & ( n30638 )  ;
assign n31918 =  ( n92 ) & ( n30640 )  ;
assign n31919 =  ( n92 ) & ( n30642 )  ;
assign n31920 =  ( n92 ) & ( n30644 )  ;
assign n31921 =  ( n92 ) & ( n30646 )  ;
assign n31922 =  ( n93 ) & ( n30616 )  ;
assign n31923 =  ( n93 ) & ( n30618 )  ;
assign n31924 =  ( n93 ) & ( n30620 )  ;
assign n31925 =  ( n93 ) & ( n30622 )  ;
assign n31926 =  ( n93 ) & ( n30624 )  ;
assign n31927 =  ( n93 ) & ( n30626 )  ;
assign n31928 =  ( n93 ) & ( n30628 )  ;
assign n31929 =  ( n93 ) & ( n30630 )  ;
assign n31930 =  ( n93 ) & ( n30632 )  ;
assign n31931 =  ( n93 ) & ( n30634 )  ;
assign n31932 =  ( n93 ) & ( n30636 )  ;
assign n31933 =  ( n93 ) & ( n30638 )  ;
assign n31934 =  ( n93 ) & ( n30640 )  ;
assign n31935 =  ( n93 ) & ( n30642 )  ;
assign n31936 =  ( n93 ) & ( n30644 )  ;
assign n31937 =  ( n93 ) & ( n30646 )  ;
assign n31938 =  ( n94 ) & ( n30616 )  ;
assign n31939 =  ( n94 ) & ( n30618 )  ;
assign n31940 =  ( n94 ) & ( n30620 )  ;
assign n31941 =  ( n94 ) & ( n30622 )  ;
assign n31942 =  ( n94 ) & ( n30624 )  ;
assign n31943 =  ( n94 ) & ( n30626 )  ;
assign n31944 =  ( n94 ) & ( n30628 )  ;
assign n31945 =  ( n94 ) & ( n30630 )  ;
assign n31946 =  ( n94 ) & ( n30632 )  ;
assign n31947 =  ( n94 ) & ( n30634 )  ;
assign n31948 =  ( n94 ) & ( n30636 )  ;
assign n31949 =  ( n94 ) & ( n30638 )  ;
assign n31950 =  ( n94 ) & ( n30640 )  ;
assign n31951 =  ( n94 ) & ( n30642 )  ;
assign n31952 =  ( n94 ) & ( n30644 )  ;
assign n31953 =  ( n94 ) & ( n30646 )  ;
assign n31954 =  ( n95 ) & ( n30616 )  ;
assign n31955 =  ( n95 ) & ( n30618 )  ;
assign n31956 =  ( n95 ) & ( n30620 )  ;
assign n31957 =  ( n95 ) & ( n30622 )  ;
assign n31958 =  ( n95 ) & ( n30624 )  ;
assign n31959 =  ( n95 ) & ( n30626 )  ;
assign n31960 =  ( n95 ) & ( n30628 )  ;
assign n31961 =  ( n95 ) & ( n30630 )  ;
assign n31962 =  ( n95 ) & ( n30632 )  ;
assign n31963 =  ( n95 ) & ( n30634 )  ;
assign n31964 =  ( n95 ) & ( n30636 )  ;
assign n31965 =  ( n95 ) & ( n30638 )  ;
assign n31966 =  ( n95 ) & ( n30640 )  ;
assign n31967 =  ( n95 ) & ( n30642 )  ;
assign n31968 =  ( n95 ) & ( n30644 )  ;
assign n31969 =  ( n95 ) & ( n30646 )  ;
assign n31970 =  ( n96 ) & ( n30616 )  ;
assign n31971 =  ( n96 ) & ( n30618 )  ;
assign n31972 =  ( n96 ) & ( n30620 )  ;
assign n31973 =  ( n96 ) & ( n30622 )  ;
assign n31974 =  ( n96 ) & ( n30624 )  ;
assign n31975 =  ( n96 ) & ( n30626 )  ;
assign n31976 =  ( n96 ) & ( n30628 )  ;
assign n31977 =  ( n96 ) & ( n30630 )  ;
assign n31978 =  ( n96 ) & ( n30632 )  ;
assign n31979 =  ( n96 ) & ( n30634 )  ;
assign n31980 =  ( n96 ) & ( n30636 )  ;
assign n31981 =  ( n96 ) & ( n30638 )  ;
assign n31982 =  ( n96 ) & ( n30640 )  ;
assign n31983 =  ( n96 ) & ( n30642 )  ;
assign n31984 =  ( n96 ) & ( n30644 )  ;
assign n31985 =  ( n96 ) & ( n30646 )  ;
assign n31986 =  ( n97 ) & ( n30616 )  ;
assign n31987 =  ( n97 ) & ( n30618 )  ;
assign n31988 =  ( n97 ) & ( n30620 )  ;
assign n31989 =  ( n97 ) & ( n30622 )  ;
assign n31990 =  ( n97 ) & ( n30624 )  ;
assign n31991 =  ( n97 ) & ( n30626 )  ;
assign n31992 =  ( n97 ) & ( n30628 )  ;
assign n31993 =  ( n97 ) & ( n30630 )  ;
assign n31994 =  ( n97 ) & ( n30632 )  ;
assign n31995 =  ( n97 ) & ( n30634 )  ;
assign n31996 =  ( n97 ) & ( n30636 )  ;
assign n31997 =  ( n97 ) & ( n30638 )  ;
assign n31998 =  ( n97 ) & ( n30640 )  ;
assign n31999 =  ( n97 ) & ( n30642 )  ;
assign n32000 =  ( n97 ) & ( n30644 )  ;
assign n32001 =  ( n97 ) & ( n30646 )  ;
assign n32002 =  ( n98 ) & ( n30616 )  ;
assign n32003 =  ( n98 ) & ( n30618 )  ;
assign n32004 =  ( n98 ) & ( n30620 )  ;
assign n32005 =  ( n98 ) & ( n30622 )  ;
assign n32006 =  ( n98 ) & ( n30624 )  ;
assign n32007 =  ( n98 ) & ( n30626 )  ;
assign n32008 =  ( n98 ) & ( n30628 )  ;
assign n32009 =  ( n98 ) & ( n30630 )  ;
assign n32010 =  ( n98 ) & ( n30632 )  ;
assign n32011 =  ( n98 ) & ( n30634 )  ;
assign n32012 =  ( n98 ) & ( n30636 )  ;
assign n32013 =  ( n98 ) & ( n30638 )  ;
assign n32014 =  ( n98 ) & ( n30640 )  ;
assign n32015 =  ( n98 ) & ( n30642 )  ;
assign n32016 =  ( n98 ) & ( n30644 )  ;
assign n32017 =  ( n98 ) & ( n30646 )  ;
assign n32018 =  ( n99 ) & ( n30616 )  ;
assign n32019 =  ( n99 ) & ( n30618 )  ;
assign n32020 =  ( n99 ) & ( n30620 )  ;
assign n32021 =  ( n99 ) & ( n30622 )  ;
assign n32022 =  ( n99 ) & ( n30624 )  ;
assign n32023 =  ( n99 ) & ( n30626 )  ;
assign n32024 =  ( n99 ) & ( n30628 )  ;
assign n32025 =  ( n99 ) & ( n30630 )  ;
assign n32026 =  ( n99 ) & ( n30632 )  ;
assign n32027 =  ( n99 ) & ( n30634 )  ;
assign n32028 =  ( n99 ) & ( n30636 )  ;
assign n32029 =  ( n99 ) & ( n30638 )  ;
assign n32030 =  ( n99 ) & ( n30640 )  ;
assign n32031 =  ( n99 ) & ( n30642 )  ;
assign n32032 =  ( n99 ) & ( n30644 )  ;
assign n32033 =  ( n99 ) & ( n30646 )  ;
assign n32034 =  ( n100 ) & ( n30616 )  ;
assign n32035 =  ( n100 ) & ( n30618 )  ;
assign n32036 =  ( n100 ) & ( n30620 )  ;
assign n32037 =  ( n100 ) & ( n30622 )  ;
assign n32038 =  ( n100 ) & ( n30624 )  ;
assign n32039 =  ( n100 ) & ( n30626 )  ;
assign n32040 =  ( n100 ) & ( n30628 )  ;
assign n32041 =  ( n100 ) & ( n30630 )  ;
assign n32042 =  ( n100 ) & ( n30632 )  ;
assign n32043 =  ( n100 ) & ( n30634 )  ;
assign n32044 =  ( n100 ) & ( n30636 )  ;
assign n32045 =  ( n100 ) & ( n30638 )  ;
assign n32046 =  ( n100 ) & ( n30640 )  ;
assign n32047 =  ( n100 ) & ( n30642 )  ;
assign n32048 =  ( n100 ) & ( n30644 )  ;
assign n32049 =  ( n100 ) & ( n30646 )  ;
assign n32050 =  ( n101 ) & ( n30616 )  ;
assign n32051 =  ( n101 ) & ( n30618 )  ;
assign n32052 =  ( n101 ) & ( n30620 )  ;
assign n32053 =  ( n101 ) & ( n30622 )  ;
assign n32054 =  ( n101 ) & ( n30624 )  ;
assign n32055 =  ( n101 ) & ( n30626 )  ;
assign n32056 =  ( n101 ) & ( n30628 )  ;
assign n32057 =  ( n101 ) & ( n30630 )  ;
assign n32058 =  ( n101 ) & ( n30632 )  ;
assign n32059 =  ( n101 ) & ( n30634 )  ;
assign n32060 =  ( n101 ) & ( n30636 )  ;
assign n32061 =  ( n101 ) & ( n30638 )  ;
assign n32062 =  ( n101 ) & ( n30640 )  ;
assign n32063 =  ( n101 ) & ( n30642 )  ;
assign n32064 =  ( n101 ) & ( n30644 )  ;
assign n32065 =  ( n101 ) & ( n30646 )  ;
assign n32066 =  ( n102 ) & ( n30616 )  ;
assign n32067 =  ( n102 ) & ( n30618 )  ;
assign n32068 =  ( n102 ) & ( n30620 )  ;
assign n32069 =  ( n102 ) & ( n30622 )  ;
assign n32070 =  ( n102 ) & ( n30624 )  ;
assign n32071 =  ( n102 ) & ( n30626 )  ;
assign n32072 =  ( n102 ) & ( n30628 )  ;
assign n32073 =  ( n102 ) & ( n30630 )  ;
assign n32074 =  ( n102 ) & ( n30632 )  ;
assign n32075 =  ( n102 ) & ( n30634 )  ;
assign n32076 =  ( n102 ) & ( n30636 )  ;
assign n32077 =  ( n102 ) & ( n30638 )  ;
assign n32078 =  ( n102 ) & ( n30640 )  ;
assign n32079 =  ( n102 ) & ( n30642 )  ;
assign n32080 =  ( n102 ) & ( n30644 )  ;
assign n32081 =  ( n102 ) & ( n30646 )  ;
assign n32082 =  ( n103 ) & ( n30616 )  ;
assign n32083 =  ( n103 ) & ( n30618 )  ;
assign n32084 =  ( n103 ) & ( n30620 )  ;
assign n32085 =  ( n103 ) & ( n30622 )  ;
assign n32086 =  ( n103 ) & ( n30624 )  ;
assign n32087 =  ( n103 ) & ( n30626 )  ;
assign n32088 =  ( n103 ) & ( n30628 )  ;
assign n32089 =  ( n103 ) & ( n30630 )  ;
assign n32090 =  ( n103 ) & ( n30632 )  ;
assign n32091 =  ( n103 ) & ( n30634 )  ;
assign n32092 =  ( n103 ) & ( n30636 )  ;
assign n32093 =  ( n103 ) & ( n30638 )  ;
assign n32094 =  ( n103 ) & ( n30640 )  ;
assign n32095 =  ( n103 ) & ( n30642 )  ;
assign n32096 =  ( n103 ) & ( n30644 )  ;
assign n32097 =  ( n103 ) & ( n30646 )  ;
assign n32098 =  ( n104 ) & ( n30616 )  ;
assign n32099 =  ( n104 ) & ( n30618 )  ;
assign n32100 =  ( n104 ) & ( n30620 )  ;
assign n32101 =  ( n104 ) & ( n30622 )  ;
assign n32102 =  ( n104 ) & ( n30624 )  ;
assign n32103 =  ( n104 ) & ( n30626 )  ;
assign n32104 =  ( n104 ) & ( n30628 )  ;
assign n32105 =  ( n104 ) & ( n30630 )  ;
assign n32106 =  ( n104 ) & ( n30632 )  ;
assign n32107 =  ( n104 ) & ( n30634 )  ;
assign n32108 =  ( n104 ) & ( n30636 )  ;
assign n32109 =  ( n104 ) & ( n30638 )  ;
assign n32110 =  ( n104 ) & ( n30640 )  ;
assign n32111 =  ( n104 ) & ( n30642 )  ;
assign n32112 =  ( n104 ) & ( n30644 )  ;
assign n32113 =  ( n104 ) & ( n30646 )  ;
assign n32114 =  ( n105 ) & ( n30616 )  ;
assign n32115 =  ( n105 ) & ( n30618 )  ;
assign n32116 =  ( n105 ) & ( n30620 )  ;
assign n32117 =  ( n105 ) & ( n30622 )  ;
assign n32118 =  ( n105 ) & ( n30624 )  ;
assign n32119 =  ( n105 ) & ( n30626 )  ;
assign n32120 =  ( n105 ) & ( n30628 )  ;
assign n32121 =  ( n105 ) & ( n30630 )  ;
assign n32122 =  ( n105 ) & ( n30632 )  ;
assign n32123 =  ( n105 ) & ( n30634 )  ;
assign n32124 =  ( n105 ) & ( n30636 )  ;
assign n32125 =  ( n105 ) & ( n30638 )  ;
assign n32126 =  ( n105 ) & ( n30640 )  ;
assign n32127 =  ( n105 ) & ( n30642 )  ;
assign n32128 =  ( n105 ) & ( n30644 )  ;
assign n32129 =  ( n105 ) & ( n30646 )  ;
assign n32130 =  ( n106 ) & ( n30616 )  ;
assign n32131 =  ( n106 ) & ( n30618 )  ;
assign n32132 =  ( n106 ) & ( n30620 )  ;
assign n32133 =  ( n106 ) & ( n30622 )  ;
assign n32134 =  ( n106 ) & ( n30624 )  ;
assign n32135 =  ( n106 ) & ( n30626 )  ;
assign n32136 =  ( n106 ) & ( n30628 )  ;
assign n32137 =  ( n106 ) & ( n30630 )  ;
assign n32138 =  ( n106 ) & ( n30632 )  ;
assign n32139 =  ( n106 ) & ( n30634 )  ;
assign n32140 =  ( n106 ) & ( n30636 )  ;
assign n32141 =  ( n106 ) & ( n30638 )  ;
assign n32142 =  ( n106 ) & ( n30640 )  ;
assign n32143 =  ( n106 ) & ( n30642 )  ;
assign n32144 =  ( n106 ) & ( n30644 )  ;
assign n32145 =  ( n106 ) & ( n30646 )  ;
assign n32146 =  ( n107 ) & ( n30616 )  ;
assign n32147 =  ( n107 ) & ( n30618 )  ;
assign n32148 =  ( n107 ) & ( n30620 )  ;
assign n32149 =  ( n107 ) & ( n30622 )  ;
assign n32150 =  ( n107 ) & ( n30624 )  ;
assign n32151 =  ( n107 ) & ( n30626 )  ;
assign n32152 =  ( n107 ) & ( n30628 )  ;
assign n32153 =  ( n107 ) & ( n30630 )  ;
assign n32154 =  ( n107 ) & ( n30632 )  ;
assign n32155 =  ( n107 ) & ( n30634 )  ;
assign n32156 =  ( n107 ) & ( n30636 )  ;
assign n32157 =  ( n107 ) & ( n30638 )  ;
assign n32158 =  ( n107 ) & ( n30640 )  ;
assign n32159 =  ( n107 ) & ( n30642 )  ;
assign n32160 =  ( n107 ) & ( n30644 )  ;
assign n32161 =  ( n107 ) & ( n30646 )  ;
assign n32162 =  ( n108 ) & ( n30616 )  ;
assign n32163 =  ( n108 ) & ( n30618 )  ;
assign n32164 =  ( n108 ) & ( n30620 )  ;
assign n32165 =  ( n108 ) & ( n30622 )  ;
assign n32166 =  ( n108 ) & ( n30624 )  ;
assign n32167 =  ( n108 ) & ( n30626 )  ;
assign n32168 =  ( n108 ) & ( n30628 )  ;
assign n32169 =  ( n108 ) & ( n30630 )  ;
assign n32170 =  ( n108 ) & ( n30632 )  ;
assign n32171 =  ( n108 ) & ( n30634 )  ;
assign n32172 =  ( n108 ) & ( n30636 )  ;
assign n32173 =  ( n108 ) & ( n30638 )  ;
assign n32174 =  ( n108 ) & ( n30640 )  ;
assign n32175 =  ( n108 ) & ( n30642 )  ;
assign n32176 =  ( n108 ) & ( n30644 )  ;
assign n32177 =  ( n108 ) & ( n30646 )  ;
assign n32178 =  ( n32177 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n32179 =  ( n32176 ) ? ( VREG_0_1 ) : ( n32178 ) ;
assign n32180 =  ( n32175 ) ? ( VREG_0_2 ) : ( n32179 ) ;
assign n32181 =  ( n32174 ) ? ( VREG_0_3 ) : ( n32180 ) ;
assign n32182 =  ( n32173 ) ? ( VREG_0_4 ) : ( n32181 ) ;
assign n32183 =  ( n32172 ) ? ( VREG_0_5 ) : ( n32182 ) ;
assign n32184 =  ( n32171 ) ? ( VREG_0_6 ) : ( n32183 ) ;
assign n32185 =  ( n32170 ) ? ( VREG_0_7 ) : ( n32184 ) ;
assign n32186 =  ( n32169 ) ? ( VREG_0_8 ) : ( n32185 ) ;
assign n32187 =  ( n32168 ) ? ( VREG_0_9 ) : ( n32186 ) ;
assign n32188 =  ( n32167 ) ? ( VREG_0_10 ) : ( n32187 ) ;
assign n32189 =  ( n32166 ) ? ( VREG_0_11 ) : ( n32188 ) ;
assign n32190 =  ( n32165 ) ? ( VREG_0_12 ) : ( n32189 ) ;
assign n32191 =  ( n32164 ) ? ( VREG_0_13 ) : ( n32190 ) ;
assign n32192 =  ( n32163 ) ? ( VREG_0_14 ) : ( n32191 ) ;
assign n32193 =  ( n32162 ) ? ( VREG_0_15 ) : ( n32192 ) ;
assign n32194 =  ( n32161 ) ? ( VREG_1_0 ) : ( n32193 ) ;
assign n32195 =  ( n32160 ) ? ( VREG_1_1 ) : ( n32194 ) ;
assign n32196 =  ( n32159 ) ? ( VREG_1_2 ) : ( n32195 ) ;
assign n32197 =  ( n32158 ) ? ( VREG_1_3 ) : ( n32196 ) ;
assign n32198 =  ( n32157 ) ? ( VREG_1_4 ) : ( n32197 ) ;
assign n32199 =  ( n32156 ) ? ( VREG_1_5 ) : ( n32198 ) ;
assign n32200 =  ( n32155 ) ? ( VREG_1_6 ) : ( n32199 ) ;
assign n32201 =  ( n32154 ) ? ( VREG_1_7 ) : ( n32200 ) ;
assign n32202 =  ( n32153 ) ? ( VREG_1_8 ) : ( n32201 ) ;
assign n32203 =  ( n32152 ) ? ( VREG_1_9 ) : ( n32202 ) ;
assign n32204 =  ( n32151 ) ? ( VREG_1_10 ) : ( n32203 ) ;
assign n32205 =  ( n32150 ) ? ( VREG_1_11 ) : ( n32204 ) ;
assign n32206 =  ( n32149 ) ? ( VREG_1_12 ) : ( n32205 ) ;
assign n32207 =  ( n32148 ) ? ( VREG_1_13 ) : ( n32206 ) ;
assign n32208 =  ( n32147 ) ? ( VREG_1_14 ) : ( n32207 ) ;
assign n32209 =  ( n32146 ) ? ( VREG_1_15 ) : ( n32208 ) ;
assign n32210 =  ( n32145 ) ? ( VREG_2_0 ) : ( n32209 ) ;
assign n32211 =  ( n32144 ) ? ( VREG_2_1 ) : ( n32210 ) ;
assign n32212 =  ( n32143 ) ? ( VREG_2_2 ) : ( n32211 ) ;
assign n32213 =  ( n32142 ) ? ( VREG_2_3 ) : ( n32212 ) ;
assign n32214 =  ( n32141 ) ? ( VREG_2_4 ) : ( n32213 ) ;
assign n32215 =  ( n32140 ) ? ( VREG_2_5 ) : ( n32214 ) ;
assign n32216 =  ( n32139 ) ? ( VREG_2_6 ) : ( n32215 ) ;
assign n32217 =  ( n32138 ) ? ( VREG_2_7 ) : ( n32216 ) ;
assign n32218 =  ( n32137 ) ? ( VREG_2_8 ) : ( n32217 ) ;
assign n32219 =  ( n32136 ) ? ( VREG_2_9 ) : ( n32218 ) ;
assign n32220 =  ( n32135 ) ? ( VREG_2_10 ) : ( n32219 ) ;
assign n32221 =  ( n32134 ) ? ( VREG_2_11 ) : ( n32220 ) ;
assign n32222 =  ( n32133 ) ? ( VREG_2_12 ) : ( n32221 ) ;
assign n32223 =  ( n32132 ) ? ( VREG_2_13 ) : ( n32222 ) ;
assign n32224 =  ( n32131 ) ? ( VREG_2_14 ) : ( n32223 ) ;
assign n32225 =  ( n32130 ) ? ( VREG_2_15 ) : ( n32224 ) ;
assign n32226 =  ( n32129 ) ? ( VREG_3_0 ) : ( n32225 ) ;
assign n32227 =  ( n32128 ) ? ( VREG_3_1 ) : ( n32226 ) ;
assign n32228 =  ( n32127 ) ? ( VREG_3_2 ) : ( n32227 ) ;
assign n32229 =  ( n32126 ) ? ( VREG_3_3 ) : ( n32228 ) ;
assign n32230 =  ( n32125 ) ? ( VREG_3_4 ) : ( n32229 ) ;
assign n32231 =  ( n32124 ) ? ( VREG_3_5 ) : ( n32230 ) ;
assign n32232 =  ( n32123 ) ? ( VREG_3_6 ) : ( n32231 ) ;
assign n32233 =  ( n32122 ) ? ( VREG_3_7 ) : ( n32232 ) ;
assign n32234 =  ( n32121 ) ? ( VREG_3_8 ) : ( n32233 ) ;
assign n32235 =  ( n32120 ) ? ( VREG_3_9 ) : ( n32234 ) ;
assign n32236 =  ( n32119 ) ? ( VREG_3_10 ) : ( n32235 ) ;
assign n32237 =  ( n32118 ) ? ( VREG_3_11 ) : ( n32236 ) ;
assign n32238 =  ( n32117 ) ? ( VREG_3_12 ) : ( n32237 ) ;
assign n32239 =  ( n32116 ) ? ( VREG_3_13 ) : ( n32238 ) ;
assign n32240 =  ( n32115 ) ? ( VREG_3_14 ) : ( n32239 ) ;
assign n32241 =  ( n32114 ) ? ( VREG_3_15 ) : ( n32240 ) ;
assign n32242 =  ( n32113 ) ? ( VREG_4_0 ) : ( n32241 ) ;
assign n32243 =  ( n32112 ) ? ( VREG_4_1 ) : ( n32242 ) ;
assign n32244 =  ( n32111 ) ? ( VREG_4_2 ) : ( n32243 ) ;
assign n32245 =  ( n32110 ) ? ( VREG_4_3 ) : ( n32244 ) ;
assign n32246 =  ( n32109 ) ? ( VREG_4_4 ) : ( n32245 ) ;
assign n32247 =  ( n32108 ) ? ( VREG_4_5 ) : ( n32246 ) ;
assign n32248 =  ( n32107 ) ? ( VREG_4_6 ) : ( n32247 ) ;
assign n32249 =  ( n32106 ) ? ( VREG_4_7 ) : ( n32248 ) ;
assign n32250 =  ( n32105 ) ? ( VREG_4_8 ) : ( n32249 ) ;
assign n32251 =  ( n32104 ) ? ( VREG_4_9 ) : ( n32250 ) ;
assign n32252 =  ( n32103 ) ? ( VREG_4_10 ) : ( n32251 ) ;
assign n32253 =  ( n32102 ) ? ( VREG_4_11 ) : ( n32252 ) ;
assign n32254 =  ( n32101 ) ? ( VREG_4_12 ) : ( n32253 ) ;
assign n32255 =  ( n32100 ) ? ( VREG_4_13 ) : ( n32254 ) ;
assign n32256 =  ( n32099 ) ? ( VREG_4_14 ) : ( n32255 ) ;
assign n32257 =  ( n32098 ) ? ( VREG_4_15 ) : ( n32256 ) ;
assign n32258 =  ( n32097 ) ? ( VREG_5_0 ) : ( n32257 ) ;
assign n32259 =  ( n32096 ) ? ( VREG_5_1 ) : ( n32258 ) ;
assign n32260 =  ( n32095 ) ? ( VREG_5_2 ) : ( n32259 ) ;
assign n32261 =  ( n32094 ) ? ( VREG_5_3 ) : ( n32260 ) ;
assign n32262 =  ( n32093 ) ? ( VREG_5_4 ) : ( n32261 ) ;
assign n32263 =  ( n32092 ) ? ( VREG_5_5 ) : ( n32262 ) ;
assign n32264 =  ( n32091 ) ? ( VREG_5_6 ) : ( n32263 ) ;
assign n32265 =  ( n32090 ) ? ( VREG_5_7 ) : ( n32264 ) ;
assign n32266 =  ( n32089 ) ? ( VREG_5_8 ) : ( n32265 ) ;
assign n32267 =  ( n32088 ) ? ( VREG_5_9 ) : ( n32266 ) ;
assign n32268 =  ( n32087 ) ? ( VREG_5_10 ) : ( n32267 ) ;
assign n32269 =  ( n32086 ) ? ( VREG_5_11 ) : ( n32268 ) ;
assign n32270 =  ( n32085 ) ? ( VREG_5_12 ) : ( n32269 ) ;
assign n32271 =  ( n32084 ) ? ( VREG_5_13 ) : ( n32270 ) ;
assign n32272 =  ( n32083 ) ? ( VREG_5_14 ) : ( n32271 ) ;
assign n32273 =  ( n32082 ) ? ( VREG_5_15 ) : ( n32272 ) ;
assign n32274 =  ( n32081 ) ? ( VREG_6_0 ) : ( n32273 ) ;
assign n32275 =  ( n32080 ) ? ( VREG_6_1 ) : ( n32274 ) ;
assign n32276 =  ( n32079 ) ? ( VREG_6_2 ) : ( n32275 ) ;
assign n32277 =  ( n32078 ) ? ( VREG_6_3 ) : ( n32276 ) ;
assign n32278 =  ( n32077 ) ? ( VREG_6_4 ) : ( n32277 ) ;
assign n32279 =  ( n32076 ) ? ( VREG_6_5 ) : ( n32278 ) ;
assign n32280 =  ( n32075 ) ? ( VREG_6_6 ) : ( n32279 ) ;
assign n32281 =  ( n32074 ) ? ( VREG_6_7 ) : ( n32280 ) ;
assign n32282 =  ( n32073 ) ? ( VREG_6_8 ) : ( n32281 ) ;
assign n32283 =  ( n32072 ) ? ( VREG_6_9 ) : ( n32282 ) ;
assign n32284 =  ( n32071 ) ? ( VREG_6_10 ) : ( n32283 ) ;
assign n32285 =  ( n32070 ) ? ( VREG_6_11 ) : ( n32284 ) ;
assign n32286 =  ( n32069 ) ? ( VREG_6_12 ) : ( n32285 ) ;
assign n32287 =  ( n32068 ) ? ( VREG_6_13 ) : ( n32286 ) ;
assign n32288 =  ( n32067 ) ? ( VREG_6_14 ) : ( n32287 ) ;
assign n32289 =  ( n32066 ) ? ( VREG_6_15 ) : ( n32288 ) ;
assign n32290 =  ( n32065 ) ? ( VREG_7_0 ) : ( n32289 ) ;
assign n32291 =  ( n32064 ) ? ( VREG_7_1 ) : ( n32290 ) ;
assign n32292 =  ( n32063 ) ? ( VREG_7_2 ) : ( n32291 ) ;
assign n32293 =  ( n32062 ) ? ( VREG_7_3 ) : ( n32292 ) ;
assign n32294 =  ( n32061 ) ? ( VREG_7_4 ) : ( n32293 ) ;
assign n32295 =  ( n32060 ) ? ( VREG_7_5 ) : ( n32294 ) ;
assign n32296 =  ( n32059 ) ? ( VREG_7_6 ) : ( n32295 ) ;
assign n32297 =  ( n32058 ) ? ( VREG_7_7 ) : ( n32296 ) ;
assign n32298 =  ( n32057 ) ? ( VREG_7_8 ) : ( n32297 ) ;
assign n32299 =  ( n32056 ) ? ( VREG_7_9 ) : ( n32298 ) ;
assign n32300 =  ( n32055 ) ? ( VREG_7_10 ) : ( n32299 ) ;
assign n32301 =  ( n32054 ) ? ( VREG_7_11 ) : ( n32300 ) ;
assign n32302 =  ( n32053 ) ? ( VREG_7_12 ) : ( n32301 ) ;
assign n32303 =  ( n32052 ) ? ( VREG_7_13 ) : ( n32302 ) ;
assign n32304 =  ( n32051 ) ? ( VREG_7_14 ) : ( n32303 ) ;
assign n32305 =  ( n32050 ) ? ( VREG_7_15 ) : ( n32304 ) ;
assign n32306 =  ( n32049 ) ? ( VREG_8_0 ) : ( n32305 ) ;
assign n32307 =  ( n32048 ) ? ( VREG_8_1 ) : ( n32306 ) ;
assign n32308 =  ( n32047 ) ? ( VREG_8_2 ) : ( n32307 ) ;
assign n32309 =  ( n32046 ) ? ( VREG_8_3 ) : ( n32308 ) ;
assign n32310 =  ( n32045 ) ? ( VREG_8_4 ) : ( n32309 ) ;
assign n32311 =  ( n32044 ) ? ( VREG_8_5 ) : ( n32310 ) ;
assign n32312 =  ( n32043 ) ? ( VREG_8_6 ) : ( n32311 ) ;
assign n32313 =  ( n32042 ) ? ( VREG_8_7 ) : ( n32312 ) ;
assign n32314 =  ( n32041 ) ? ( VREG_8_8 ) : ( n32313 ) ;
assign n32315 =  ( n32040 ) ? ( VREG_8_9 ) : ( n32314 ) ;
assign n32316 =  ( n32039 ) ? ( VREG_8_10 ) : ( n32315 ) ;
assign n32317 =  ( n32038 ) ? ( VREG_8_11 ) : ( n32316 ) ;
assign n32318 =  ( n32037 ) ? ( VREG_8_12 ) : ( n32317 ) ;
assign n32319 =  ( n32036 ) ? ( VREG_8_13 ) : ( n32318 ) ;
assign n32320 =  ( n32035 ) ? ( VREG_8_14 ) : ( n32319 ) ;
assign n32321 =  ( n32034 ) ? ( VREG_8_15 ) : ( n32320 ) ;
assign n32322 =  ( n32033 ) ? ( VREG_9_0 ) : ( n32321 ) ;
assign n32323 =  ( n32032 ) ? ( VREG_9_1 ) : ( n32322 ) ;
assign n32324 =  ( n32031 ) ? ( VREG_9_2 ) : ( n32323 ) ;
assign n32325 =  ( n32030 ) ? ( VREG_9_3 ) : ( n32324 ) ;
assign n32326 =  ( n32029 ) ? ( VREG_9_4 ) : ( n32325 ) ;
assign n32327 =  ( n32028 ) ? ( VREG_9_5 ) : ( n32326 ) ;
assign n32328 =  ( n32027 ) ? ( VREG_9_6 ) : ( n32327 ) ;
assign n32329 =  ( n32026 ) ? ( VREG_9_7 ) : ( n32328 ) ;
assign n32330 =  ( n32025 ) ? ( VREG_9_8 ) : ( n32329 ) ;
assign n32331 =  ( n32024 ) ? ( VREG_9_9 ) : ( n32330 ) ;
assign n32332 =  ( n32023 ) ? ( VREG_9_10 ) : ( n32331 ) ;
assign n32333 =  ( n32022 ) ? ( VREG_9_11 ) : ( n32332 ) ;
assign n32334 =  ( n32021 ) ? ( VREG_9_12 ) : ( n32333 ) ;
assign n32335 =  ( n32020 ) ? ( VREG_9_13 ) : ( n32334 ) ;
assign n32336 =  ( n32019 ) ? ( VREG_9_14 ) : ( n32335 ) ;
assign n32337 =  ( n32018 ) ? ( VREG_9_15 ) : ( n32336 ) ;
assign n32338 =  ( n32017 ) ? ( VREG_10_0 ) : ( n32337 ) ;
assign n32339 =  ( n32016 ) ? ( VREG_10_1 ) : ( n32338 ) ;
assign n32340 =  ( n32015 ) ? ( VREG_10_2 ) : ( n32339 ) ;
assign n32341 =  ( n32014 ) ? ( VREG_10_3 ) : ( n32340 ) ;
assign n32342 =  ( n32013 ) ? ( VREG_10_4 ) : ( n32341 ) ;
assign n32343 =  ( n32012 ) ? ( VREG_10_5 ) : ( n32342 ) ;
assign n32344 =  ( n32011 ) ? ( VREG_10_6 ) : ( n32343 ) ;
assign n32345 =  ( n32010 ) ? ( VREG_10_7 ) : ( n32344 ) ;
assign n32346 =  ( n32009 ) ? ( VREG_10_8 ) : ( n32345 ) ;
assign n32347 =  ( n32008 ) ? ( VREG_10_9 ) : ( n32346 ) ;
assign n32348 =  ( n32007 ) ? ( VREG_10_10 ) : ( n32347 ) ;
assign n32349 =  ( n32006 ) ? ( VREG_10_11 ) : ( n32348 ) ;
assign n32350 =  ( n32005 ) ? ( VREG_10_12 ) : ( n32349 ) ;
assign n32351 =  ( n32004 ) ? ( VREG_10_13 ) : ( n32350 ) ;
assign n32352 =  ( n32003 ) ? ( VREG_10_14 ) : ( n32351 ) ;
assign n32353 =  ( n32002 ) ? ( VREG_10_15 ) : ( n32352 ) ;
assign n32354 =  ( n32001 ) ? ( VREG_11_0 ) : ( n32353 ) ;
assign n32355 =  ( n32000 ) ? ( VREG_11_1 ) : ( n32354 ) ;
assign n32356 =  ( n31999 ) ? ( VREG_11_2 ) : ( n32355 ) ;
assign n32357 =  ( n31998 ) ? ( VREG_11_3 ) : ( n32356 ) ;
assign n32358 =  ( n31997 ) ? ( VREG_11_4 ) : ( n32357 ) ;
assign n32359 =  ( n31996 ) ? ( VREG_11_5 ) : ( n32358 ) ;
assign n32360 =  ( n31995 ) ? ( VREG_11_6 ) : ( n32359 ) ;
assign n32361 =  ( n31994 ) ? ( VREG_11_7 ) : ( n32360 ) ;
assign n32362 =  ( n31993 ) ? ( VREG_11_8 ) : ( n32361 ) ;
assign n32363 =  ( n31992 ) ? ( VREG_11_9 ) : ( n32362 ) ;
assign n32364 =  ( n31991 ) ? ( VREG_11_10 ) : ( n32363 ) ;
assign n32365 =  ( n31990 ) ? ( VREG_11_11 ) : ( n32364 ) ;
assign n32366 =  ( n31989 ) ? ( VREG_11_12 ) : ( n32365 ) ;
assign n32367 =  ( n31988 ) ? ( VREG_11_13 ) : ( n32366 ) ;
assign n32368 =  ( n31987 ) ? ( VREG_11_14 ) : ( n32367 ) ;
assign n32369 =  ( n31986 ) ? ( VREG_11_15 ) : ( n32368 ) ;
assign n32370 =  ( n31985 ) ? ( VREG_12_0 ) : ( n32369 ) ;
assign n32371 =  ( n31984 ) ? ( VREG_12_1 ) : ( n32370 ) ;
assign n32372 =  ( n31983 ) ? ( VREG_12_2 ) : ( n32371 ) ;
assign n32373 =  ( n31982 ) ? ( VREG_12_3 ) : ( n32372 ) ;
assign n32374 =  ( n31981 ) ? ( VREG_12_4 ) : ( n32373 ) ;
assign n32375 =  ( n31980 ) ? ( VREG_12_5 ) : ( n32374 ) ;
assign n32376 =  ( n31979 ) ? ( VREG_12_6 ) : ( n32375 ) ;
assign n32377 =  ( n31978 ) ? ( VREG_12_7 ) : ( n32376 ) ;
assign n32378 =  ( n31977 ) ? ( VREG_12_8 ) : ( n32377 ) ;
assign n32379 =  ( n31976 ) ? ( VREG_12_9 ) : ( n32378 ) ;
assign n32380 =  ( n31975 ) ? ( VREG_12_10 ) : ( n32379 ) ;
assign n32381 =  ( n31974 ) ? ( VREG_12_11 ) : ( n32380 ) ;
assign n32382 =  ( n31973 ) ? ( VREG_12_12 ) : ( n32381 ) ;
assign n32383 =  ( n31972 ) ? ( VREG_12_13 ) : ( n32382 ) ;
assign n32384 =  ( n31971 ) ? ( VREG_12_14 ) : ( n32383 ) ;
assign n32385 =  ( n31970 ) ? ( VREG_12_15 ) : ( n32384 ) ;
assign n32386 =  ( n31969 ) ? ( VREG_13_0 ) : ( n32385 ) ;
assign n32387 =  ( n31968 ) ? ( VREG_13_1 ) : ( n32386 ) ;
assign n32388 =  ( n31967 ) ? ( VREG_13_2 ) : ( n32387 ) ;
assign n32389 =  ( n31966 ) ? ( VREG_13_3 ) : ( n32388 ) ;
assign n32390 =  ( n31965 ) ? ( VREG_13_4 ) : ( n32389 ) ;
assign n32391 =  ( n31964 ) ? ( VREG_13_5 ) : ( n32390 ) ;
assign n32392 =  ( n31963 ) ? ( VREG_13_6 ) : ( n32391 ) ;
assign n32393 =  ( n31962 ) ? ( VREG_13_7 ) : ( n32392 ) ;
assign n32394 =  ( n31961 ) ? ( VREG_13_8 ) : ( n32393 ) ;
assign n32395 =  ( n31960 ) ? ( VREG_13_9 ) : ( n32394 ) ;
assign n32396 =  ( n31959 ) ? ( VREG_13_10 ) : ( n32395 ) ;
assign n32397 =  ( n31958 ) ? ( VREG_13_11 ) : ( n32396 ) ;
assign n32398 =  ( n31957 ) ? ( VREG_13_12 ) : ( n32397 ) ;
assign n32399 =  ( n31956 ) ? ( VREG_13_13 ) : ( n32398 ) ;
assign n32400 =  ( n31955 ) ? ( VREG_13_14 ) : ( n32399 ) ;
assign n32401 =  ( n31954 ) ? ( VREG_13_15 ) : ( n32400 ) ;
assign n32402 =  ( n31953 ) ? ( VREG_14_0 ) : ( n32401 ) ;
assign n32403 =  ( n31952 ) ? ( VREG_14_1 ) : ( n32402 ) ;
assign n32404 =  ( n31951 ) ? ( VREG_14_2 ) : ( n32403 ) ;
assign n32405 =  ( n31950 ) ? ( VREG_14_3 ) : ( n32404 ) ;
assign n32406 =  ( n31949 ) ? ( VREG_14_4 ) : ( n32405 ) ;
assign n32407 =  ( n31948 ) ? ( VREG_14_5 ) : ( n32406 ) ;
assign n32408 =  ( n31947 ) ? ( VREG_14_6 ) : ( n32407 ) ;
assign n32409 =  ( n31946 ) ? ( VREG_14_7 ) : ( n32408 ) ;
assign n32410 =  ( n31945 ) ? ( VREG_14_8 ) : ( n32409 ) ;
assign n32411 =  ( n31944 ) ? ( VREG_14_9 ) : ( n32410 ) ;
assign n32412 =  ( n31943 ) ? ( VREG_14_10 ) : ( n32411 ) ;
assign n32413 =  ( n31942 ) ? ( VREG_14_11 ) : ( n32412 ) ;
assign n32414 =  ( n31941 ) ? ( VREG_14_12 ) : ( n32413 ) ;
assign n32415 =  ( n31940 ) ? ( VREG_14_13 ) : ( n32414 ) ;
assign n32416 =  ( n31939 ) ? ( VREG_14_14 ) : ( n32415 ) ;
assign n32417 =  ( n31938 ) ? ( VREG_14_15 ) : ( n32416 ) ;
assign n32418 =  ( n31937 ) ? ( VREG_15_0 ) : ( n32417 ) ;
assign n32419 =  ( n31936 ) ? ( VREG_15_1 ) : ( n32418 ) ;
assign n32420 =  ( n31935 ) ? ( VREG_15_2 ) : ( n32419 ) ;
assign n32421 =  ( n31934 ) ? ( VREG_15_3 ) : ( n32420 ) ;
assign n32422 =  ( n31933 ) ? ( VREG_15_4 ) : ( n32421 ) ;
assign n32423 =  ( n31932 ) ? ( VREG_15_5 ) : ( n32422 ) ;
assign n32424 =  ( n31931 ) ? ( VREG_15_6 ) : ( n32423 ) ;
assign n32425 =  ( n31930 ) ? ( VREG_15_7 ) : ( n32424 ) ;
assign n32426 =  ( n31929 ) ? ( VREG_15_8 ) : ( n32425 ) ;
assign n32427 =  ( n31928 ) ? ( VREG_15_9 ) : ( n32426 ) ;
assign n32428 =  ( n31927 ) ? ( VREG_15_10 ) : ( n32427 ) ;
assign n32429 =  ( n31926 ) ? ( VREG_15_11 ) : ( n32428 ) ;
assign n32430 =  ( n31925 ) ? ( VREG_15_12 ) : ( n32429 ) ;
assign n32431 =  ( n31924 ) ? ( VREG_15_13 ) : ( n32430 ) ;
assign n32432 =  ( n31923 ) ? ( VREG_15_14 ) : ( n32431 ) ;
assign n32433 =  ( n31922 ) ? ( VREG_15_15 ) : ( n32432 ) ;
assign n32434 =  ( n31921 ) ? ( VREG_16_0 ) : ( n32433 ) ;
assign n32435 =  ( n31920 ) ? ( VREG_16_1 ) : ( n32434 ) ;
assign n32436 =  ( n31919 ) ? ( VREG_16_2 ) : ( n32435 ) ;
assign n32437 =  ( n31918 ) ? ( VREG_16_3 ) : ( n32436 ) ;
assign n32438 =  ( n31917 ) ? ( VREG_16_4 ) : ( n32437 ) ;
assign n32439 =  ( n31916 ) ? ( VREG_16_5 ) : ( n32438 ) ;
assign n32440 =  ( n31915 ) ? ( VREG_16_6 ) : ( n32439 ) ;
assign n32441 =  ( n31914 ) ? ( VREG_16_7 ) : ( n32440 ) ;
assign n32442 =  ( n31913 ) ? ( VREG_16_8 ) : ( n32441 ) ;
assign n32443 =  ( n31912 ) ? ( VREG_16_9 ) : ( n32442 ) ;
assign n32444 =  ( n31911 ) ? ( VREG_16_10 ) : ( n32443 ) ;
assign n32445 =  ( n31910 ) ? ( VREG_16_11 ) : ( n32444 ) ;
assign n32446 =  ( n31909 ) ? ( VREG_16_12 ) : ( n32445 ) ;
assign n32447 =  ( n31908 ) ? ( VREG_16_13 ) : ( n32446 ) ;
assign n32448 =  ( n31907 ) ? ( VREG_16_14 ) : ( n32447 ) ;
assign n32449 =  ( n31906 ) ? ( VREG_16_15 ) : ( n32448 ) ;
assign n32450 =  ( n31905 ) ? ( VREG_17_0 ) : ( n32449 ) ;
assign n32451 =  ( n31904 ) ? ( VREG_17_1 ) : ( n32450 ) ;
assign n32452 =  ( n31903 ) ? ( VREG_17_2 ) : ( n32451 ) ;
assign n32453 =  ( n31902 ) ? ( VREG_17_3 ) : ( n32452 ) ;
assign n32454 =  ( n31901 ) ? ( VREG_17_4 ) : ( n32453 ) ;
assign n32455 =  ( n31900 ) ? ( VREG_17_5 ) : ( n32454 ) ;
assign n32456 =  ( n31899 ) ? ( VREG_17_6 ) : ( n32455 ) ;
assign n32457 =  ( n31898 ) ? ( VREG_17_7 ) : ( n32456 ) ;
assign n32458 =  ( n31897 ) ? ( VREG_17_8 ) : ( n32457 ) ;
assign n32459 =  ( n31896 ) ? ( VREG_17_9 ) : ( n32458 ) ;
assign n32460 =  ( n31895 ) ? ( VREG_17_10 ) : ( n32459 ) ;
assign n32461 =  ( n31894 ) ? ( VREG_17_11 ) : ( n32460 ) ;
assign n32462 =  ( n31893 ) ? ( VREG_17_12 ) : ( n32461 ) ;
assign n32463 =  ( n31892 ) ? ( VREG_17_13 ) : ( n32462 ) ;
assign n32464 =  ( n31891 ) ? ( VREG_17_14 ) : ( n32463 ) ;
assign n32465 =  ( n31890 ) ? ( VREG_17_15 ) : ( n32464 ) ;
assign n32466 =  ( n31889 ) ? ( VREG_18_0 ) : ( n32465 ) ;
assign n32467 =  ( n31888 ) ? ( VREG_18_1 ) : ( n32466 ) ;
assign n32468 =  ( n31887 ) ? ( VREG_18_2 ) : ( n32467 ) ;
assign n32469 =  ( n31886 ) ? ( VREG_18_3 ) : ( n32468 ) ;
assign n32470 =  ( n31885 ) ? ( VREG_18_4 ) : ( n32469 ) ;
assign n32471 =  ( n31884 ) ? ( VREG_18_5 ) : ( n32470 ) ;
assign n32472 =  ( n31883 ) ? ( VREG_18_6 ) : ( n32471 ) ;
assign n32473 =  ( n31882 ) ? ( VREG_18_7 ) : ( n32472 ) ;
assign n32474 =  ( n31881 ) ? ( VREG_18_8 ) : ( n32473 ) ;
assign n32475 =  ( n31880 ) ? ( VREG_18_9 ) : ( n32474 ) ;
assign n32476 =  ( n31879 ) ? ( VREG_18_10 ) : ( n32475 ) ;
assign n32477 =  ( n31878 ) ? ( VREG_18_11 ) : ( n32476 ) ;
assign n32478 =  ( n31877 ) ? ( VREG_18_12 ) : ( n32477 ) ;
assign n32479 =  ( n31876 ) ? ( VREG_18_13 ) : ( n32478 ) ;
assign n32480 =  ( n31875 ) ? ( VREG_18_14 ) : ( n32479 ) ;
assign n32481 =  ( n31874 ) ? ( VREG_18_15 ) : ( n32480 ) ;
assign n32482 =  ( n31873 ) ? ( VREG_19_0 ) : ( n32481 ) ;
assign n32483 =  ( n31872 ) ? ( VREG_19_1 ) : ( n32482 ) ;
assign n32484 =  ( n31871 ) ? ( VREG_19_2 ) : ( n32483 ) ;
assign n32485 =  ( n31870 ) ? ( VREG_19_3 ) : ( n32484 ) ;
assign n32486 =  ( n31869 ) ? ( VREG_19_4 ) : ( n32485 ) ;
assign n32487 =  ( n31868 ) ? ( VREG_19_5 ) : ( n32486 ) ;
assign n32488 =  ( n31867 ) ? ( VREG_19_6 ) : ( n32487 ) ;
assign n32489 =  ( n31866 ) ? ( VREG_19_7 ) : ( n32488 ) ;
assign n32490 =  ( n31865 ) ? ( VREG_19_8 ) : ( n32489 ) ;
assign n32491 =  ( n31864 ) ? ( VREG_19_9 ) : ( n32490 ) ;
assign n32492 =  ( n31863 ) ? ( VREG_19_10 ) : ( n32491 ) ;
assign n32493 =  ( n31862 ) ? ( VREG_19_11 ) : ( n32492 ) ;
assign n32494 =  ( n31861 ) ? ( VREG_19_12 ) : ( n32493 ) ;
assign n32495 =  ( n31860 ) ? ( VREG_19_13 ) : ( n32494 ) ;
assign n32496 =  ( n31859 ) ? ( VREG_19_14 ) : ( n32495 ) ;
assign n32497 =  ( n31858 ) ? ( VREG_19_15 ) : ( n32496 ) ;
assign n32498 =  ( n31857 ) ? ( VREG_20_0 ) : ( n32497 ) ;
assign n32499 =  ( n31856 ) ? ( VREG_20_1 ) : ( n32498 ) ;
assign n32500 =  ( n31855 ) ? ( VREG_20_2 ) : ( n32499 ) ;
assign n32501 =  ( n31854 ) ? ( VREG_20_3 ) : ( n32500 ) ;
assign n32502 =  ( n31853 ) ? ( VREG_20_4 ) : ( n32501 ) ;
assign n32503 =  ( n31852 ) ? ( VREG_20_5 ) : ( n32502 ) ;
assign n32504 =  ( n31851 ) ? ( VREG_20_6 ) : ( n32503 ) ;
assign n32505 =  ( n31850 ) ? ( VREG_20_7 ) : ( n32504 ) ;
assign n32506 =  ( n31849 ) ? ( VREG_20_8 ) : ( n32505 ) ;
assign n32507 =  ( n31848 ) ? ( VREG_20_9 ) : ( n32506 ) ;
assign n32508 =  ( n31847 ) ? ( VREG_20_10 ) : ( n32507 ) ;
assign n32509 =  ( n31846 ) ? ( VREG_20_11 ) : ( n32508 ) ;
assign n32510 =  ( n31845 ) ? ( VREG_20_12 ) : ( n32509 ) ;
assign n32511 =  ( n31844 ) ? ( VREG_20_13 ) : ( n32510 ) ;
assign n32512 =  ( n31843 ) ? ( VREG_20_14 ) : ( n32511 ) ;
assign n32513 =  ( n31842 ) ? ( VREG_20_15 ) : ( n32512 ) ;
assign n32514 =  ( n31841 ) ? ( VREG_21_0 ) : ( n32513 ) ;
assign n32515 =  ( n31840 ) ? ( VREG_21_1 ) : ( n32514 ) ;
assign n32516 =  ( n31839 ) ? ( VREG_21_2 ) : ( n32515 ) ;
assign n32517 =  ( n31838 ) ? ( VREG_21_3 ) : ( n32516 ) ;
assign n32518 =  ( n31837 ) ? ( VREG_21_4 ) : ( n32517 ) ;
assign n32519 =  ( n31836 ) ? ( VREG_21_5 ) : ( n32518 ) ;
assign n32520 =  ( n31835 ) ? ( VREG_21_6 ) : ( n32519 ) ;
assign n32521 =  ( n31834 ) ? ( VREG_21_7 ) : ( n32520 ) ;
assign n32522 =  ( n31833 ) ? ( VREG_21_8 ) : ( n32521 ) ;
assign n32523 =  ( n31832 ) ? ( VREG_21_9 ) : ( n32522 ) ;
assign n32524 =  ( n31831 ) ? ( VREG_21_10 ) : ( n32523 ) ;
assign n32525 =  ( n31830 ) ? ( VREG_21_11 ) : ( n32524 ) ;
assign n32526 =  ( n31829 ) ? ( VREG_21_12 ) : ( n32525 ) ;
assign n32527 =  ( n31828 ) ? ( VREG_21_13 ) : ( n32526 ) ;
assign n32528 =  ( n31827 ) ? ( VREG_21_14 ) : ( n32527 ) ;
assign n32529 =  ( n31826 ) ? ( VREG_21_15 ) : ( n32528 ) ;
assign n32530 =  ( n31825 ) ? ( VREG_22_0 ) : ( n32529 ) ;
assign n32531 =  ( n31824 ) ? ( VREG_22_1 ) : ( n32530 ) ;
assign n32532 =  ( n31823 ) ? ( VREG_22_2 ) : ( n32531 ) ;
assign n32533 =  ( n31822 ) ? ( VREG_22_3 ) : ( n32532 ) ;
assign n32534 =  ( n31821 ) ? ( VREG_22_4 ) : ( n32533 ) ;
assign n32535 =  ( n31820 ) ? ( VREG_22_5 ) : ( n32534 ) ;
assign n32536 =  ( n31819 ) ? ( VREG_22_6 ) : ( n32535 ) ;
assign n32537 =  ( n31818 ) ? ( VREG_22_7 ) : ( n32536 ) ;
assign n32538 =  ( n31817 ) ? ( VREG_22_8 ) : ( n32537 ) ;
assign n32539 =  ( n31816 ) ? ( VREG_22_9 ) : ( n32538 ) ;
assign n32540 =  ( n31815 ) ? ( VREG_22_10 ) : ( n32539 ) ;
assign n32541 =  ( n31814 ) ? ( VREG_22_11 ) : ( n32540 ) ;
assign n32542 =  ( n31813 ) ? ( VREG_22_12 ) : ( n32541 ) ;
assign n32543 =  ( n31812 ) ? ( VREG_22_13 ) : ( n32542 ) ;
assign n32544 =  ( n31811 ) ? ( VREG_22_14 ) : ( n32543 ) ;
assign n32545 =  ( n31810 ) ? ( VREG_22_15 ) : ( n32544 ) ;
assign n32546 =  ( n31809 ) ? ( VREG_23_0 ) : ( n32545 ) ;
assign n32547 =  ( n31808 ) ? ( VREG_23_1 ) : ( n32546 ) ;
assign n32548 =  ( n31807 ) ? ( VREG_23_2 ) : ( n32547 ) ;
assign n32549 =  ( n31806 ) ? ( VREG_23_3 ) : ( n32548 ) ;
assign n32550 =  ( n31805 ) ? ( VREG_23_4 ) : ( n32549 ) ;
assign n32551 =  ( n31804 ) ? ( VREG_23_5 ) : ( n32550 ) ;
assign n32552 =  ( n31803 ) ? ( VREG_23_6 ) : ( n32551 ) ;
assign n32553 =  ( n31802 ) ? ( VREG_23_7 ) : ( n32552 ) ;
assign n32554 =  ( n31801 ) ? ( VREG_23_8 ) : ( n32553 ) ;
assign n32555 =  ( n31800 ) ? ( VREG_23_9 ) : ( n32554 ) ;
assign n32556 =  ( n31799 ) ? ( VREG_23_10 ) : ( n32555 ) ;
assign n32557 =  ( n31798 ) ? ( VREG_23_11 ) : ( n32556 ) ;
assign n32558 =  ( n31797 ) ? ( VREG_23_12 ) : ( n32557 ) ;
assign n32559 =  ( n31796 ) ? ( VREG_23_13 ) : ( n32558 ) ;
assign n32560 =  ( n31795 ) ? ( VREG_23_14 ) : ( n32559 ) ;
assign n32561 =  ( n31794 ) ? ( VREG_23_15 ) : ( n32560 ) ;
assign n32562 =  ( n31793 ) ? ( VREG_24_0 ) : ( n32561 ) ;
assign n32563 =  ( n31792 ) ? ( VREG_24_1 ) : ( n32562 ) ;
assign n32564 =  ( n31791 ) ? ( VREG_24_2 ) : ( n32563 ) ;
assign n32565 =  ( n31790 ) ? ( VREG_24_3 ) : ( n32564 ) ;
assign n32566 =  ( n31789 ) ? ( VREG_24_4 ) : ( n32565 ) ;
assign n32567 =  ( n31788 ) ? ( VREG_24_5 ) : ( n32566 ) ;
assign n32568 =  ( n31787 ) ? ( VREG_24_6 ) : ( n32567 ) ;
assign n32569 =  ( n31786 ) ? ( VREG_24_7 ) : ( n32568 ) ;
assign n32570 =  ( n31785 ) ? ( VREG_24_8 ) : ( n32569 ) ;
assign n32571 =  ( n31784 ) ? ( VREG_24_9 ) : ( n32570 ) ;
assign n32572 =  ( n31783 ) ? ( VREG_24_10 ) : ( n32571 ) ;
assign n32573 =  ( n31782 ) ? ( VREG_24_11 ) : ( n32572 ) ;
assign n32574 =  ( n31781 ) ? ( VREG_24_12 ) : ( n32573 ) ;
assign n32575 =  ( n31780 ) ? ( VREG_24_13 ) : ( n32574 ) ;
assign n32576 =  ( n31779 ) ? ( VREG_24_14 ) : ( n32575 ) ;
assign n32577 =  ( n31778 ) ? ( VREG_24_15 ) : ( n32576 ) ;
assign n32578 =  ( n31777 ) ? ( VREG_25_0 ) : ( n32577 ) ;
assign n32579 =  ( n31776 ) ? ( VREG_25_1 ) : ( n32578 ) ;
assign n32580 =  ( n31775 ) ? ( VREG_25_2 ) : ( n32579 ) ;
assign n32581 =  ( n31774 ) ? ( VREG_25_3 ) : ( n32580 ) ;
assign n32582 =  ( n31773 ) ? ( VREG_25_4 ) : ( n32581 ) ;
assign n32583 =  ( n31772 ) ? ( VREG_25_5 ) : ( n32582 ) ;
assign n32584 =  ( n31771 ) ? ( VREG_25_6 ) : ( n32583 ) ;
assign n32585 =  ( n31770 ) ? ( VREG_25_7 ) : ( n32584 ) ;
assign n32586 =  ( n31769 ) ? ( VREG_25_8 ) : ( n32585 ) ;
assign n32587 =  ( n31768 ) ? ( VREG_25_9 ) : ( n32586 ) ;
assign n32588 =  ( n31767 ) ? ( VREG_25_10 ) : ( n32587 ) ;
assign n32589 =  ( n31766 ) ? ( VREG_25_11 ) : ( n32588 ) ;
assign n32590 =  ( n31765 ) ? ( VREG_25_12 ) : ( n32589 ) ;
assign n32591 =  ( n31764 ) ? ( VREG_25_13 ) : ( n32590 ) ;
assign n32592 =  ( n31763 ) ? ( VREG_25_14 ) : ( n32591 ) ;
assign n32593 =  ( n31762 ) ? ( VREG_25_15 ) : ( n32592 ) ;
assign n32594 =  ( n31761 ) ? ( VREG_26_0 ) : ( n32593 ) ;
assign n32595 =  ( n31760 ) ? ( VREG_26_1 ) : ( n32594 ) ;
assign n32596 =  ( n31759 ) ? ( VREG_26_2 ) : ( n32595 ) ;
assign n32597 =  ( n31758 ) ? ( VREG_26_3 ) : ( n32596 ) ;
assign n32598 =  ( n31757 ) ? ( VREG_26_4 ) : ( n32597 ) ;
assign n32599 =  ( n31756 ) ? ( VREG_26_5 ) : ( n32598 ) ;
assign n32600 =  ( n31755 ) ? ( VREG_26_6 ) : ( n32599 ) ;
assign n32601 =  ( n31754 ) ? ( VREG_26_7 ) : ( n32600 ) ;
assign n32602 =  ( n31753 ) ? ( VREG_26_8 ) : ( n32601 ) ;
assign n32603 =  ( n31752 ) ? ( VREG_26_9 ) : ( n32602 ) ;
assign n32604 =  ( n31751 ) ? ( VREG_26_10 ) : ( n32603 ) ;
assign n32605 =  ( n31750 ) ? ( VREG_26_11 ) : ( n32604 ) ;
assign n32606 =  ( n31749 ) ? ( VREG_26_12 ) : ( n32605 ) ;
assign n32607 =  ( n31748 ) ? ( VREG_26_13 ) : ( n32606 ) ;
assign n32608 =  ( n31747 ) ? ( VREG_26_14 ) : ( n32607 ) ;
assign n32609 =  ( n31746 ) ? ( VREG_26_15 ) : ( n32608 ) ;
assign n32610 =  ( n31745 ) ? ( VREG_27_0 ) : ( n32609 ) ;
assign n32611 =  ( n31744 ) ? ( VREG_27_1 ) : ( n32610 ) ;
assign n32612 =  ( n31743 ) ? ( VREG_27_2 ) : ( n32611 ) ;
assign n32613 =  ( n31742 ) ? ( VREG_27_3 ) : ( n32612 ) ;
assign n32614 =  ( n31741 ) ? ( VREG_27_4 ) : ( n32613 ) ;
assign n32615 =  ( n31740 ) ? ( VREG_27_5 ) : ( n32614 ) ;
assign n32616 =  ( n31739 ) ? ( VREG_27_6 ) : ( n32615 ) ;
assign n32617 =  ( n31738 ) ? ( VREG_27_7 ) : ( n32616 ) ;
assign n32618 =  ( n31737 ) ? ( VREG_27_8 ) : ( n32617 ) ;
assign n32619 =  ( n31736 ) ? ( VREG_27_9 ) : ( n32618 ) ;
assign n32620 =  ( n31735 ) ? ( VREG_27_10 ) : ( n32619 ) ;
assign n32621 =  ( n31734 ) ? ( VREG_27_11 ) : ( n32620 ) ;
assign n32622 =  ( n31733 ) ? ( VREG_27_12 ) : ( n32621 ) ;
assign n32623 =  ( n31732 ) ? ( VREG_27_13 ) : ( n32622 ) ;
assign n32624 =  ( n31731 ) ? ( VREG_27_14 ) : ( n32623 ) ;
assign n32625 =  ( n31730 ) ? ( VREG_27_15 ) : ( n32624 ) ;
assign n32626 =  ( n31729 ) ? ( VREG_28_0 ) : ( n32625 ) ;
assign n32627 =  ( n31728 ) ? ( VREG_28_1 ) : ( n32626 ) ;
assign n32628 =  ( n31727 ) ? ( VREG_28_2 ) : ( n32627 ) ;
assign n32629 =  ( n31726 ) ? ( VREG_28_3 ) : ( n32628 ) ;
assign n32630 =  ( n31725 ) ? ( VREG_28_4 ) : ( n32629 ) ;
assign n32631 =  ( n31724 ) ? ( VREG_28_5 ) : ( n32630 ) ;
assign n32632 =  ( n31723 ) ? ( VREG_28_6 ) : ( n32631 ) ;
assign n32633 =  ( n31722 ) ? ( VREG_28_7 ) : ( n32632 ) ;
assign n32634 =  ( n31721 ) ? ( VREG_28_8 ) : ( n32633 ) ;
assign n32635 =  ( n31720 ) ? ( VREG_28_9 ) : ( n32634 ) ;
assign n32636 =  ( n31719 ) ? ( VREG_28_10 ) : ( n32635 ) ;
assign n32637 =  ( n31718 ) ? ( VREG_28_11 ) : ( n32636 ) ;
assign n32638 =  ( n31717 ) ? ( VREG_28_12 ) : ( n32637 ) ;
assign n32639 =  ( n31716 ) ? ( VREG_28_13 ) : ( n32638 ) ;
assign n32640 =  ( n31715 ) ? ( VREG_28_14 ) : ( n32639 ) ;
assign n32641 =  ( n31714 ) ? ( VREG_28_15 ) : ( n32640 ) ;
assign n32642 =  ( n31713 ) ? ( VREG_29_0 ) : ( n32641 ) ;
assign n32643 =  ( n31712 ) ? ( VREG_29_1 ) : ( n32642 ) ;
assign n32644 =  ( n31711 ) ? ( VREG_29_2 ) : ( n32643 ) ;
assign n32645 =  ( n31710 ) ? ( VREG_29_3 ) : ( n32644 ) ;
assign n32646 =  ( n31709 ) ? ( VREG_29_4 ) : ( n32645 ) ;
assign n32647 =  ( n31708 ) ? ( VREG_29_5 ) : ( n32646 ) ;
assign n32648 =  ( n31707 ) ? ( VREG_29_6 ) : ( n32647 ) ;
assign n32649 =  ( n31706 ) ? ( VREG_29_7 ) : ( n32648 ) ;
assign n32650 =  ( n31705 ) ? ( VREG_29_8 ) : ( n32649 ) ;
assign n32651 =  ( n31704 ) ? ( VREG_29_9 ) : ( n32650 ) ;
assign n32652 =  ( n31703 ) ? ( VREG_29_10 ) : ( n32651 ) ;
assign n32653 =  ( n31702 ) ? ( VREG_29_11 ) : ( n32652 ) ;
assign n32654 =  ( n31701 ) ? ( VREG_29_12 ) : ( n32653 ) ;
assign n32655 =  ( n31700 ) ? ( VREG_29_13 ) : ( n32654 ) ;
assign n32656 =  ( n31699 ) ? ( VREG_29_14 ) : ( n32655 ) ;
assign n32657 =  ( n31698 ) ? ( VREG_29_15 ) : ( n32656 ) ;
assign n32658 =  ( n31697 ) ? ( VREG_30_0 ) : ( n32657 ) ;
assign n32659 =  ( n31696 ) ? ( VREG_30_1 ) : ( n32658 ) ;
assign n32660 =  ( n31695 ) ? ( VREG_30_2 ) : ( n32659 ) ;
assign n32661 =  ( n31694 ) ? ( VREG_30_3 ) : ( n32660 ) ;
assign n32662 =  ( n31693 ) ? ( VREG_30_4 ) : ( n32661 ) ;
assign n32663 =  ( n31692 ) ? ( VREG_30_5 ) : ( n32662 ) ;
assign n32664 =  ( n31691 ) ? ( VREG_30_6 ) : ( n32663 ) ;
assign n32665 =  ( n31690 ) ? ( VREG_30_7 ) : ( n32664 ) ;
assign n32666 =  ( n31689 ) ? ( VREG_30_8 ) : ( n32665 ) ;
assign n32667 =  ( n31688 ) ? ( VREG_30_9 ) : ( n32666 ) ;
assign n32668 =  ( n31687 ) ? ( VREG_30_10 ) : ( n32667 ) ;
assign n32669 =  ( n31686 ) ? ( VREG_30_11 ) : ( n32668 ) ;
assign n32670 =  ( n31685 ) ? ( VREG_30_12 ) : ( n32669 ) ;
assign n32671 =  ( n31684 ) ? ( VREG_30_13 ) : ( n32670 ) ;
assign n32672 =  ( n31683 ) ? ( VREG_30_14 ) : ( n32671 ) ;
assign n32673 =  ( n31682 ) ? ( VREG_30_15 ) : ( n32672 ) ;
assign n32674 =  ( n31681 ) ? ( VREG_31_0 ) : ( n32673 ) ;
assign n32675 =  ( n31680 ) ? ( VREG_31_1 ) : ( n32674 ) ;
assign n32676 =  ( n31679 ) ? ( VREG_31_2 ) : ( n32675 ) ;
assign n32677 =  ( n31678 ) ? ( VREG_31_3 ) : ( n32676 ) ;
assign n32678 =  ( n31677 ) ? ( VREG_31_4 ) : ( n32677 ) ;
assign n32679 =  ( n31676 ) ? ( VREG_31_5 ) : ( n32678 ) ;
assign n32680 =  ( n31675 ) ? ( VREG_31_6 ) : ( n32679 ) ;
assign n32681 =  ( n31674 ) ? ( VREG_31_7 ) : ( n32680 ) ;
assign n32682 =  ( n31673 ) ? ( VREG_31_8 ) : ( n32681 ) ;
assign n32683 =  ( n31672 ) ? ( VREG_31_9 ) : ( n32682 ) ;
assign n32684 =  ( n31671 ) ? ( VREG_31_10 ) : ( n32683 ) ;
assign n32685 =  ( n31670 ) ? ( VREG_31_11 ) : ( n32684 ) ;
assign n32686 =  ( n31669 ) ? ( VREG_31_12 ) : ( n32685 ) ;
assign n32687 =  ( n31668 ) ? ( VREG_31_13 ) : ( n32686 ) ;
assign n32688 =  ( n31667 ) ? ( VREG_31_14 ) : ( n32687 ) ;
assign n32689 =  ( n31666 ) ? ( VREG_31_15 ) : ( n32688 ) ;
assign n32690 =  ( n31655 ) + ( n32689 )  ;
assign n32691 =  ( n31655 ) - ( n32689 )  ;
assign n32692 =  ( n31655 ) & ( n32689 )  ;
assign n32693 =  ( n31655 ) | ( n32689 )  ;
assign n32694 =  ( ( n31655 ) * ( n32689 ))  ;
assign n32695 =  ( n148 ) ? ( n32694 ) : ( VREG_0_8 ) ;
assign n32696 =  ( n146 ) ? ( n32693 ) : ( n32695 ) ;
assign n32697 =  ( n144 ) ? ( n32692 ) : ( n32696 ) ;
assign n32698 =  ( n142 ) ? ( n32691 ) : ( n32697 ) ;
assign n32699 =  ( n10 ) ? ( n32690 ) : ( n32698 ) ;
assign n32700 = n3030[8:8] ;
assign n32701 =  ( n32700 ) == ( 1'd0 )  ;
assign n32702 =  ( n32701 ) ? ( VREG_0_8 ) : ( n31665 ) ;
assign n32703 =  ( n32701 ) ? ( VREG_0_8 ) : ( n32699 ) ;
assign n32704 =  ( n3034 ) ? ( n32703 ) : ( VREG_0_8 ) ;
assign n32705 =  ( n2965 ) ? ( n32702 ) : ( n32704 ) ;
assign n32706 =  ( n1930 ) ? ( n32699 ) : ( n32705 ) ;
assign n32707 =  ( n879 ) ? ( n31665 ) : ( n32706 ) ;
assign n32708 =  ( n31655 ) + ( n164 )  ;
assign n32709 =  ( n31655 ) - ( n164 )  ;
assign n32710 =  ( n31655 ) & ( n164 )  ;
assign n32711 =  ( n31655 ) | ( n164 )  ;
assign n32712 =  ( ( n31655 ) * ( n164 ))  ;
assign n32713 =  ( n172 ) ? ( n32712 ) : ( VREG_0_8 ) ;
assign n32714 =  ( n170 ) ? ( n32711 ) : ( n32713 ) ;
assign n32715 =  ( n168 ) ? ( n32710 ) : ( n32714 ) ;
assign n32716 =  ( n166 ) ? ( n32709 ) : ( n32715 ) ;
assign n32717 =  ( n162 ) ? ( n32708 ) : ( n32716 ) ;
assign n32718 =  ( n31655 ) + ( n180 )  ;
assign n32719 =  ( n31655 ) - ( n180 )  ;
assign n32720 =  ( n31655 ) & ( n180 )  ;
assign n32721 =  ( n31655 ) | ( n180 )  ;
assign n32722 =  ( ( n31655 ) * ( n180 ))  ;
assign n32723 =  ( n172 ) ? ( n32722 ) : ( VREG_0_8 ) ;
assign n32724 =  ( n170 ) ? ( n32721 ) : ( n32723 ) ;
assign n32725 =  ( n168 ) ? ( n32720 ) : ( n32724 ) ;
assign n32726 =  ( n166 ) ? ( n32719 ) : ( n32725 ) ;
assign n32727 =  ( n162 ) ? ( n32718 ) : ( n32726 ) ;
assign n32728 =  ( n32701 ) ? ( VREG_0_8 ) : ( n32727 ) ;
assign n32729 =  ( n3051 ) ? ( n32728 ) : ( VREG_0_8 ) ;
assign n32730 =  ( n3040 ) ? ( n32717 ) : ( n32729 ) ;
assign n32731 =  ( n192 ) ? ( VREG_0_8 ) : ( VREG_0_8 ) ;
assign n32732 =  ( n157 ) ? ( n32730 ) : ( n32731 ) ;
assign n32733 =  ( n6 ) ? ( n32707 ) : ( n32732 ) ;
assign n32734 =  ( n4 ) ? ( n32733 ) : ( VREG_0_8 ) ;
assign n32735 =  ( 32'd9 ) == ( 32'd15 )  ;
assign n32736 =  ( n12 ) & ( n32735 )  ;
assign n32737 =  ( 32'd9 ) == ( 32'd14 )  ;
assign n32738 =  ( n12 ) & ( n32737 )  ;
assign n32739 =  ( 32'd9 ) == ( 32'd13 )  ;
assign n32740 =  ( n12 ) & ( n32739 )  ;
assign n32741 =  ( 32'd9 ) == ( 32'd12 )  ;
assign n32742 =  ( n12 ) & ( n32741 )  ;
assign n32743 =  ( 32'd9 ) == ( 32'd11 )  ;
assign n32744 =  ( n12 ) & ( n32743 )  ;
assign n32745 =  ( 32'd9 ) == ( 32'd10 )  ;
assign n32746 =  ( n12 ) & ( n32745 )  ;
assign n32747 =  ( 32'd9 ) == ( 32'd9 )  ;
assign n32748 =  ( n12 ) & ( n32747 )  ;
assign n32749 =  ( 32'd9 ) == ( 32'd8 )  ;
assign n32750 =  ( n12 ) & ( n32749 )  ;
assign n32751 =  ( 32'd9 ) == ( 32'd7 )  ;
assign n32752 =  ( n12 ) & ( n32751 )  ;
assign n32753 =  ( 32'd9 ) == ( 32'd6 )  ;
assign n32754 =  ( n12 ) & ( n32753 )  ;
assign n32755 =  ( 32'd9 ) == ( 32'd5 )  ;
assign n32756 =  ( n12 ) & ( n32755 )  ;
assign n32757 =  ( 32'd9 ) == ( 32'd4 )  ;
assign n32758 =  ( n12 ) & ( n32757 )  ;
assign n32759 =  ( 32'd9 ) == ( 32'd3 )  ;
assign n32760 =  ( n12 ) & ( n32759 )  ;
assign n32761 =  ( 32'd9 ) == ( 32'd2 )  ;
assign n32762 =  ( n12 ) & ( n32761 )  ;
assign n32763 =  ( 32'd9 ) == ( 32'd1 )  ;
assign n32764 =  ( n12 ) & ( n32763 )  ;
assign n32765 =  ( 32'd9 ) == ( 32'd0 )  ;
assign n32766 =  ( n12 ) & ( n32765 )  ;
assign n32767 =  ( n13 ) & ( n32735 )  ;
assign n32768 =  ( n13 ) & ( n32737 )  ;
assign n32769 =  ( n13 ) & ( n32739 )  ;
assign n32770 =  ( n13 ) & ( n32741 )  ;
assign n32771 =  ( n13 ) & ( n32743 )  ;
assign n32772 =  ( n13 ) & ( n32745 )  ;
assign n32773 =  ( n13 ) & ( n32747 )  ;
assign n32774 =  ( n13 ) & ( n32749 )  ;
assign n32775 =  ( n13 ) & ( n32751 )  ;
assign n32776 =  ( n13 ) & ( n32753 )  ;
assign n32777 =  ( n13 ) & ( n32755 )  ;
assign n32778 =  ( n13 ) & ( n32757 )  ;
assign n32779 =  ( n13 ) & ( n32759 )  ;
assign n32780 =  ( n13 ) & ( n32761 )  ;
assign n32781 =  ( n13 ) & ( n32763 )  ;
assign n32782 =  ( n13 ) & ( n32765 )  ;
assign n32783 =  ( n14 ) & ( n32735 )  ;
assign n32784 =  ( n14 ) & ( n32737 )  ;
assign n32785 =  ( n14 ) & ( n32739 )  ;
assign n32786 =  ( n14 ) & ( n32741 )  ;
assign n32787 =  ( n14 ) & ( n32743 )  ;
assign n32788 =  ( n14 ) & ( n32745 )  ;
assign n32789 =  ( n14 ) & ( n32747 )  ;
assign n32790 =  ( n14 ) & ( n32749 )  ;
assign n32791 =  ( n14 ) & ( n32751 )  ;
assign n32792 =  ( n14 ) & ( n32753 )  ;
assign n32793 =  ( n14 ) & ( n32755 )  ;
assign n32794 =  ( n14 ) & ( n32757 )  ;
assign n32795 =  ( n14 ) & ( n32759 )  ;
assign n32796 =  ( n14 ) & ( n32761 )  ;
assign n32797 =  ( n14 ) & ( n32763 )  ;
assign n32798 =  ( n14 ) & ( n32765 )  ;
assign n32799 =  ( n15 ) & ( n32735 )  ;
assign n32800 =  ( n15 ) & ( n32737 )  ;
assign n32801 =  ( n15 ) & ( n32739 )  ;
assign n32802 =  ( n15 ) & ( n32741 )  ;
assign n32803 =  ( n15 ) & ( n32743 )  ;
assign n32804 =  ( n15 ) & ( n32745 )  ;
assign n32805 =  ( n15 ) & ( n32747 )  ;
assign n32806 =  ( n15 ) & ( n32749 )  ;
assign n32807 =  ( n15 ) & ( n32751 )  ;
assign n32808 =  ( n15 ) & ( n32753 )  ;
assign n32809 =  ( n15 ) & ( n32755 )  ;
assign n32810 =  ( n15 ) & ( n32757 )  ;
assign n32811 =  ( n15 ) & ( n32759 )  ;
assign n32812 =  ( n15 ) & ( n32761 )  ;
assign n32813 =  ( n15 ) & ( n32763 )  ;
assign n32814 =  ( n15 ) & ( n32765 )  ;
assign n32815 =  ( n16 ) & ( n32735 )  ;
assign n32816 =  ( n16 ) & ( n32737 )  ;
assign n32817 =  ( n16 ) & ( n32739 )  ;
assign n32818 =  ( n16 ) & ( n32741 )  ;
assign n32819 =  ( n16 ) & ( n32743 )  ;
assign n32820 =  ( n16 ) & ( n32745 )  ;
assign n32821 =  ( n16 ) & ( n32747 )  ;
assign n32822 =  ( n16 ) & ( n32749 )  ;
assign n32823 =  ( n16 ) & ( n32751 )  ;
assign n32824 =  ( n16 ) & ( n32753 )  ;
assign n32825 =  ( n16 ) & ( n32755 )  ;
assign n32826 =  ( n16 ) & ( n32757 )  ;
assign n32827 =  ( n16 ) & ( n32759 )  ;
assign n32828 =  ( n16 ) & ( n32761 )  ;
assign n32829 =  ( n16 ) & ( n32763 )  ;
assign n32830 =  ( n16 ) & ( n32765 )  ;
assign n32831 =  ( n17 ) & ( n32735 )  ;
assign n32832 =  ( n17 ) & ( n32737 )  ;
assign n32833 =  ( n17 ) & ( n32739 )  ;
assign n32834 =  ( n17 ) & ( n32741 )  ;
assign n32835 =  ( n17 ) & ( n32743 )  ;
assign n32836 =  ( n17 ) & ( n32745 )  ;
assign n32837 =  ( n17 ) & ( n32747 )  ;
assign n32838 =  ( n17 ) & ( n32749 )  ;
assign n32839 =  ( n17 ) & ( n32751 )  ;
assign n32840 =  ( n17 ) & ( n32753 )  ;
assign n32841 =  ( n17 ) & ( n32755 )  ;
assign n32842 =  ( n17 ) & ( n32757 )  ;
assign n32843 =  ( n17 ) & ( n32759 )  ;
assign n32844 =  ( n17 ) & ( n32761 )  ;
assign n32845 =  ( n17 ) & ( n32763 )  ;
assign n32846 =  ( n17 ) & ( n32765 )  ;
assign n32847 =  ( n18 ) & ( n32735 )  ;
assign n32848 =  ( n18 ) & ( n32737 )  ;
assign n32849 =  ( n18 ) & ( n32739 )  ;
assign n32850 =  ( n18 ) & ( n32741 )  ;
assign n32851 =  ( n18 ) & ( n32743 )  ;
assign n32852 =  ( n18 ) & ( n32745 )  ;
assign n32853 =  ( n18 ) & ( n32747 )  ;
assign n32854 =  ( n18 ) & ( n32749 )  ;
assign n32855 =  ( n18 ) & ( n32751 )  ;
assign n32856 =  ( n18 ) & ( n32753 )  ;
assign n32857 =  ( n18 ) & ( n32755 )  ;
assign n32858 =  ( n18 ) & ( n32757 )  ;
assign n32859 =  ( n18 ) & ( n32759 )  ;
assign n32860 =  ( n18 ) & ( n32761 )  ;
assign n32861 =  ( n18 ) & ( n32763 )  ;
assign n32862 =  ( n18 ) & ( n32765 )  ;
assign n32863 =  ( n19 ) & ( n32735 )  ;
assign n32864 =  ( n19 ) & ( n32737 )  ;
assign n32865 =  ( n19 ) & ( n32739 )  ;
assign n32866 =  ( n19 ) & ( n32741 )  ;
assign n32867 =  ( n19 ) & ( n32743 )  ;
assign n32868 =  ( n19 ) & ( n32745 )  ;
assign n32869 =  ( n19 ) & ( n32747 )  ;
assign n32870 =  ( n19 ) & ( n32749 )  ;
assign n32871 =  ( n19 ) & ( n32751 )  ;
assign n32872 =  ( n19 ) & ( n32753 )  ;
assign n32873 =  ( n19 ) & ( n32755 )  ;
assign n32874 =  ( n19 ) & ( n32757 )  ;
assign n32875 =  ( n19 ) & ( n32759 )  ;
assign n32876 =  ( n19 ) & ( n32761 )  ;
assign n32877 =  ( n19 ) & ( n32763 )  ;
assign n32878 =  ( n19 ) & ( n32765 )  ;
assign n32879 =  ( n20 ) & ( n32735 )  ;
assign n32880 =  ( n20 ) & ( n32737 )  ;
assign n32881 =  ( n20 ) & ( n32739 )  ;
assign n32882 =  ( n20 ) & ( n32741 )  ;
assign n32883 =  ( n20 ) & ( n32743 )  ;
assign n32884 =  ( n20 ) & ( n32745 )  ;
assign n32885 =  ( n20 ) & ( n32747 )  ;
assign n32886 =  ( n20 ) & ( n32749 )  ;
assign n32887 =  ( n20 ) & ( n32751 )  ;
assign n32888 =  ( n20 ) & ( n32753 )  ;
assign n32889 =  ( n20 ) & ( n32755 )  ;
assign n32890 =  ( n20 ) & ( n32757 )  ;
assign n32891 =  ( n20 ) & ( n32759 )  ;
assign n32892 =  ( n20 ) & ( n32761 )  ;
assign n32893 =  ( n20 ) & ( n32763 )  ;
assign n32894 =  ( n20 ) & ( n32765 )  ;
assign n32895 =  ( n21 ) & ( n32735 )  ;
assign n32896 =  ( n21 ) & ( n32737 )  ;
assign n32897 =  ( n21 ) & ( n32739 )  ;
assign n32898 =  ( n21 ) & ( n32741 )  ;
assign n32899 =  ( n21 ) & ( n32743 )  ;
assign n32900 =  ( n21 ) & ( n32745 )  ;
assign n32901 =  ( n21 ) & ( n32747 )  ;
assign n32902 =  ( n21 ) & ( n32749 )  ;
assign n32903 =  ( n21 ) & ( n32751 )  ;
assign n32904 =  ( n21 ) & ( n32753 )  ;
assign n32905 =  ( n21 ) & ( n32755 )  ;
assign n32906 =  ( n21 ) & ( n32757 )  ;
assign n32907 =  ( n21 ) & ( n32759 )  ;
assign n32908 =  ( n21 ) & ( n32761 )  ;
assign n32909 =  ( n21 ) & ( n32763 )  ;
assign n32910 =  ( n21 ) & ( n32765 )  ;
assign n32911 =  ( n22 ) & ( n32735 )  ;
assign n32912 =  ( n22 ) & ( n32737 )  ;
assign n32913 =  ( n22 ) & ( n32739 )  ;
assign n32914 =  ( n22 ) & ( n32741 )  ;
assign n32915 =  ( n22 ) & ( n32743 )  ;
assign n32916 =  ( n22 ) & ( n32745 )  ;
assign n32917 =  ( n22 ) & ( n32747 )  ;
assign n32918 =  ( n22 ) & ( n32749 )  ;
assign n32919 =  ( n22 ) & ( n32751 )  ;
assign n32920 =  ( n22 ) & ( n32753 )  ;
assign n32921 =  ( n22 ) & ( n32755 )  ;
assign n32922 =  ( n22 ) & ( n32757 )  ;
assign n32923 =  ( n22 ) & ( n32759 )  ;
assign n32924 =  ( n22 ) & ( n32761 )  ;
assign n32925 =  ( n22 ) & ( n32763 )  ;
assign n32926 =  ( n22 ) & ( n32765 )  ;
assign n32927 =  ( n23 ) & ( n32735 )  ;
assign n32928 =  ( n23 ) & ( n32737 )  ;
assign n32929 =  ( n23 ) & ( n32739 )  ;
assign n32930 =  ( n23 ) & ( n32741 )  ;
assign n32931 =  ( n23 ) & ( n32743 )  ;
assign n32932 =  ( n23 ) & ( n32745 )  ;
assign n32933 =  ( n23 ) & ( n32747 )  ;
assign n32934 =  ( n23 ) & ( n32749 )  ;
assign n32935 =  ( n23 ) & ( n32751 )  ;
assign n32936 =  ( n23 ) & ( n32753 )  ;
assign n32937 =  ( n23 ) & ( n32755 )  ;
assign n32938 =  ( n23 ) & ( n32757 )  ;
assign n32939 =  ( n23 ) & ( n32759 )  ;
assign n32940 =  ( n23 ) & ( n32761 )  ;
assign n32941 =  ( n23 ) & ( n32763 )  ;
assign n32942 =  ( n23 ) & ( n32765 )  ;
assign n32943 =  ( n24 ) & ( n32735 )  ;
assign n32944 =  ( n24 ) & ( n32737 )  ;
assign n32945 =  ( n24 ) & ( n32739 )  ;
assign n32946 =  ( n24 ) & ( n32741 )  ;
assign n32947 =  ( n24 ) & ( n32743 )  ;
assign n32948 =  ( n24 ) & ( n32745 )  ;
assign n32949 =  ( n24 ) & ( n32747 )  ;
assign n32950 =  ( n24 ) & ( n32749 )  ;
assign n32951 =  ( n24 ) & ( n32751 )  ;
assign n32952 =  ( n24 ) & ( n32753 )  ;
assign n32953 =  ( n24 ) & ( n32755 )  ;
assign n32954 =  ( n24 ) & ( n32757 )  ;
assign n32955 =  ( n24 ) & ( n32759 )  ;
assign n32956 =  ( n24 ) & ( n32761 )  ;
assign n32957 =  ( n24 ) & ( n32763 )  ;
assign n32958 =  ( n24 ) & ( n32765 )  ;
assign n32959 =  ( n25 ) & ( n32735 )  ;
assign n32960 =  ( n25 ) & ( n32737 )  ;
assign n32961 =  ( n25 ) & ( n32739 )  ;
assign n32962 =  ( n25 ) & ( n32741 )  ;
assign n32963 =  ( n25 ) & ( n32743 )  ;
assign n32964 =  ( n25 ) & ( n32745 )  ;
assign n32965 =  ( n25 ) & ( n32747 )  ;
assign n32966 =  ( n25 ) & ( n32749 )  ;
assign n32967 =  ( n25 ) & ( n32751 )  ;
assign n32968 =  ( n25 ) & ( n32753 )  ;
assign n32969 =  ( n25 ) & ( n32755 )  ;
assign n32970 =  ( n25 ) & ( n32757 )  ;
assign n32971 =  ( n25 ) & ( n32759 )  ;
assign n32972 =  ( n25 ) & ( n32761 )  ;
assign n32973 =  ( n25 ) & ( n32763 )  ;
assign n32974 =  ( n25 ) & ( n32765 )  ;
assign n32975 =  ( n26 ) & ( n32735 )  ;
assign n32976 =  ( n26 ) & ( n32737 )  ;
assign n32977 =  ( n26 ) & ( n32739 )  ;
assign n32978 =  ( n26 ) & ( n32741 )  ;
assign n32979 =  ( n26 ) & ( n32743 )  ;
assign n32980 =  ( n26 ) & ( n32745 )  ;
assign n32981 =  ( n26 ) & ( n32747 )  ;
assign n32982 =  ( n26 ) & ( n32749 )  ;
assign n32983 =  ( n26 ) & ( n32751 )  ;
assign n32984 =  ( n26 ) & ( n32753 )  ;
assign n32985 =  ( n26 ) & ( n32755 )  ;
assign n32986 =  ( n26 ) & ( n32757 )  ;
assign n32987 =  ( n26 ) & ( n32759 )  ;
assign n32988 =  ( n26 ) & ( n32761 )  ;
assign n32989 =  ( n26 ) & ( n32763 )  ;
assign n32990 =  ( n26 ) & ( n32765 )  ;
assign n32991 =  ( n27 ) & ( n32735 )  ;
assign n32992 =  ( n27 ) & ( n32737 )  ;
assign n32993 =  ( n27 ) & ( n32739 )  ;
assign n32994 =  ( n27 ) & ( n32741 )  ;
assign n32995 =  ( n27 ) & ( n32743 )  ;
assign n32996 =  ( n27 ) & ( n32745 )  ;
assign n32997 =  ( n27 ) & ( n32747 )  ;
assign n32998 =  ( n27 ) & ( n32749 )  ;
assign n32999 =  ( n27 ) & ( n32751 )  ;
assign n33000 =  ( n27 ) & ( n32753 )  ;
assign n33001 =  ( n27 ) & ( n32755 )  ;
assign n33002 =  ( n27 ) & ( n32757 )  ;
assign n33003 =  ( n27 ) & ( n32759 )  ;
assign n33004 =  ( n27 ) & ( n32761 )  ;
assign n33005 =  ( n27 ) & ( n32763 )  ;
assign n33006 =  ( n27 ) & ( n32765 )  ;
assign n33007 =  ( n28 ) & ( n32735 )  ;
assign n33008 =  ( n28 ) & ( n32737 )  ;
assign n33009 =  ( n28 ) & ( n32739 )  ;
assign n33010 =  ( n28 ) & ( n32741 )  ;
assign n33011 =  ( n28 ) & ( n32743 )  ;
assign n33012 =  ( n28 ) & ( n32745 )  ;
assign n33013 =  ( n28 ) & ( n32747 )  ;
assign n33014 =  ( n28 ) & ( n32749 )  ;
assign n33015 =  ( n28 ) & ( n32751 )  ;
assign n33016 =  ( n28 ) & ( n32753 )  ;
assign n33017 =  ( n28 ) & ( n32755 )  ;
assign n33018 =  ( n28 ) & ( n32757 )  ;
assign n33019 =  ( n28 ) & ( n32759 )  ;
assign n33020 =  ( n28 ) & ( n32761 )  ;
assign n33021 =  ( n28 ) & ( n32763 )  ;
assign n33022 =  ( n28 ) & ( n32765 )  ;
assign n33023 =  ( n29 ) & ( n32735 )  ;
assign n33024 =  ( n29 ) & ( n32737 )  ;
assign n33025 =  ( n29 ) & ( n32739 )  ;
assign n33026 =  ( n29 ) & ( n32741 )  ;
assign n33027 =  ( n29 ) & ( n32743 )  ;
assign n33028 =  ( n29 ) & ( n32745 )  ;
assign n33029 =  ( n29 ) & ( n32747 )  ;
assign n33030 =  ( n29 ) & ( n32749 )  ;
assign n33031 =  ( n29 ) & ( n32751 )  ;
assign n33032 =  ( n29 ) & ( n32753 )  ;
assign n33033 =  ( n29 ) & ( n32755 )  ;
assign n33034 =  ( n29 ) & ( n32757 )  ;
assign n33035 =  ( n29 ) & ( n32759 )  ;
assign n33036 =  ( n29 ) & ( n32761 )  ;
assign n33037 =  ( n29 ) & ( n32763 )  ;
assign n33038 =  ( n29 ) & ( n32765 )  ;
assign n33039 =  ( n30 ) & ( n32735 )  ;
assign n33040 =  ( n30 ) & ( n32737 )  ;
assign n33041 =  ( n30 ) & ( n32739 )  ;
assign n33042 =  ( n30 ) & ( n32741 )  ;
assign n33043 =  ( n30 ) & ( n32743 )  ;
assign n33044 =  ( n30 ) & ( n32745 )  ;
assign n33045 =  ( n30 ) & ( n32747 )  ;
assign n33046 =  ( n30 ) & ( n32749 )  ;
assign n33047 =  ( n30 ) & ( n32751 )  ;
assign n33048 =  ( n30 ) & ( n32753 )  ;
assign n33049 =  ( n30 ) & ( n32755 )  ;
assign n33050 =  ( n30 ) & ( n32757 )  ;
assign n33051 =  ( n30 ) & ( n32759 )  ;
assign n33052 =  ( n30 ) & ( n32761 )  ;
assign n33053 =  ( n30 ) & ( n32763 )  ;
assign n33054 =  ( n30 ) & ( n32765 )  ;
assign n33055 =  ( n31 ) & ( n32735 )  ;
assign n33056 =  ( n31 ) & ( n32737 )  ;
assign n33057 =  ( n31 ) & ( n32739 )  ;
assign n33058 =  ( n31 ) & ( n32741 )  ;
assign n33059 =  ( n31 ) & ( n32743 )  ;
assign n33060 =  ( n31 ) & ( n32745 )  ;
assign n33061 =  ( n31 ) & ( n32747 )  ;
assign n33062 =  ( n31 ) & ( n32749 )  ;
assign n33063 =  ( n31 ) & ( n32751 )  ;
assign n33064 =  ( n31 ) & ( n32753 )  ;
assign n33065 =  ( n31 ) & ( n32755 )  ;
assign n33066 =  ( n31 ) & ( n32757 )  ;
assign n33067 =  ( n31 ) & ( n32759 )  ;
assign n33068 =  ( n31 ) & ( n32761 )  ;
assign n33069 =  ( n31 ) & ( n32763 )  ;
assign n33070 =  ( n31 ) & ( n32765 )  ;
assign n33071 =  ( n32 ) & ( n32735 )  ;
assign n33072 =  ( n32 ) & ( n32737 )  ;
assign n33073 =  ( n32 ) & ( n32739 )  ;
assign n33074 =  ( n32 ) & ( n32741 )  ;
assign n33075 =  ( n32 ) & ( n32743 )  ;
assign n33076 =  ( n32 ) & ( n32745 )  ;
assign n33077 =  ( n32 ) & ( n32747 )  ;
assign n33078 =  ( n32 ) & ( n32749 )  ;
assign n33079 =  ( n32 ) & ( n32751 )  ;
assign n33080 =  ( n32 ) & ( n32753 )  ;
assign n33081 =  ( n32 ) & ( n32755 )  ;
assign n33082 =  ( n32 ) & ( n32757 )  ;
assign n33083 =  ( n32 ) & ( n32759 )  ;
assign n33084 =  ( n32 ) & ( n32761 )  ;
assign n33085 =  ( n32 ) & ( n32763 )  ;
assign n33086 =  ( n32 ) & ( n32765 )  ;
assign n33087 =  ( n33 ) & ( n32735 )  ;
assign n33088 =  ( n33 ) & ( n32737 )  ;
assign n33089 =  ( n33 ) & ( n32739 )  ;
assign n33090 =  ( n33 ) & ( n32741 )  ;
assign n33091 =  ( n33 ) & ( n32743 )  ;
assign n33092 =  ( n33 ) & ( n32745 )  ;
assign n33093 =  ( n33 ) & ( n32747 )  ;
assign n33094 =  ( n33 ) & ( n32749 )  ;
assign n33095 =  ( n33 ) & ( n32751 )  ;
assign n33096 =  ( n33 ) & ( n32753 )  ;
assign n33097 =  ( n33 ) & ( n32755 )  ;
assign n33098 =  ( n33 ) & ( n32757 )  ;
assign n33099 =  ( n33 ) & ( n32759 )  ;
assign n33100 =  ( n33 ) & ( n32761 )  ;
assign n33101 =  ( n33 ) & ( n32763 )  ;
assign n33102 =  ( n33 ) & ( n32765 )  ;
assign n33103 =  ( n34 ) & ( n32735 )  ;
assign n33104 =  ( n34 ) & ( n32737 )  ;
assign n33105 =  ( n34 ) & ( n32739 )  ;
assign n33106 =  ( n34 ) & ( n32741 )  ;
assign n33107 =  ( n34 ) & ( n32743 )  ;
assign n33108 =  ( n34 ) & ( n32745 )  ;
assign n33109 =  ( n34 ) & ( n32747 )  ;
assign n33110 =  ( n34 ) & ( n32749 )  ;
assign n33111 =  ( n34 ) & ( n32751 )  ;
assign n33112 =  ( n34 ) & ( n32753 )  ;
assign n33113 =  ( n34 ) & ( n32755 )  ;
assign n33114 =  ( n34 ) & ( n32757 )  ;
assign n33115 =  ( n34 ) & ( n32759 )  ;
assign n33116 =  ( n34 ) & ( n32761 )  ;
assign n33117 =  ( n34 ) & ( n32763 )  ;
assign n33118 =  ( n34 ) & ( n32765 )  ;
assign n33119 =  ( n35 ) & ( n32735 )  ;
assign n33120 =  ( n35 ) & ( n32737 )  ;
assign n33121 =  ( n35 ) & ( n32739 )  ;
assign n33122 =  ( n35 ) & ( n32741 )  ;
assign n33123 =  ( n35 ) & ( n32743 )  ;
assign n33124 =  ( n35 ) & ( n32745 )  ;
assign n33125 =  ( n35 ) & ( n32747 )  ;
assign n33126 =  ( n35 ) & ( n32749 )  ;
assign n33127 =  ( n35 ) & ( n32751 )  ;
assign n33128 =  ( n35 ) & ( n32753 )  ;
assign n33129 =  ( n35 ) & ( n32755 )  ;
assign n33130 =  ( n35 ) & ( n32757 )  ;
assign n33131 =  ( n35 ) & ( n32759 )  ;
assign n33132 =  ( n35 ) & ( n32761 )  ;
assign n33133 =  ( n35 ) & ( n32763 )  ;
assign n33134 =  ( n35 ) & ( n32765 )  ;
assign n33135 =  ( n36 ) & ( n32735 )  ;
assign n33136 =  ( n36 ) & ( n32737 )  ;
assign n33137 =  ( n36 ) & ( n32739 )  ;
assign n33138 =  ( n36 ) & ( n32741 )  ;
assign n33139 =  ( n36 ) & ( n32743 )  ;
assign n33140 =  ( n36 ) & ( n32745 )  ;
assign n33141 =  ( n36 ) & ( n32747 )  ;
assign n33142 =  ( n36 ) & ( n32749 )  ;
assign n33143 =  ( n36 ) & ( n32751 )  ;
assign n33144 =  ( n36 ) & ( n32753 )  ;
assign n33145 =  ( n36 ) & ( n32755 )  ;
assign n33146 =  ( n36 ) & ( n32757 )  ;
assign n33147 =  ( n36 ) & ( n32759 )  ;
assign n33148 =  ( n36 ) & ( n32761 )  ;
assign n33149 =  ( n36 ) & ( n32763 )  ;
assign n33150 =  ( n36 ) & ( n32765 )  ;
assign n33151 =  ( n37 ) & ( n32735 )  ;
assign n33152 =  ( n37 ) & ( n32737 )  ;
assign n33153 =  ( n37 ) & ( n32739 )  ;
assign n33154 =  ( n37 ) & ( n32741 )  ;
assign n33155 =  ( n37 ) & ( n32743 )  ;
assign n33156 =  ( n37 ) & ( n32745 )  ;
assign n33157 =  ( n37 ) & ( n32747 )  ;
assign n33158 =  ( n37 ) & ( n32749 )  ;
assign n33159 =  ( n37 ) & ( n32751 )  ;
assign n33160 =  ( n37 ) & ( n32753 )  ;
assign n33161 =  ( n37 ) & ( n32755 )  ;
assign n33162 =  ( n37 ) & ( n32757 )  ;
assign n33163 =  ( n37 ) & ( n32759 )  ;
assign n33164 =  ( n37 ) & ( n32761 )  ;
assign n33165 =  ( n37 ) & ( n32763 )  ;
assign n33166 =  ( n37 ) & ( n32765 )  ;
assign n33167 =  ( n38 ) & ( n32735 )  ;
assign n33168 =  ( n38 ) & ( n32737 )  ;
assign n33169 =  ( n38 ) & ( n32739 )  ;
assign n33170 =  ( n38 ) & ( n32741 )  ;
assign n33171 =  ( n38 ) & ( n32743 )  ;
assign n33172 =  ( n38 ) & ( n32745 )  ;
assign n33173 =  ( n38 ) & ( n32747 )  ;
assign n33174 =  ( n38 ) & ( n32749 )  ;
assign n33175 =  ( n38 ) & ( n32751 )  ;
assign n33176 =  ( n38 ) & ( n32753 )  ;
assign n33177 =  ( n38 ) & ( n32755 )  ;
assign n33178 =  ( n38 ) & ( n32757 )  ;
assign n33179 =  ( n38 ) & ( n32759 )  ;
assign n33180 =  ( n38 ) & ( n32761 )  ;
assign n33181 =  ( n38 ) & ( n32763 )  ;
assign n33182 =  ( n38 ) & ( n32765 )  ;
assign n33183 =  ( n39 ) & ( n32735 )  ;
assign n33184 =  ( n39 ) & ( n32737 )  ;
assign n33185 =  ( n39 ) & ( n32739 )  ;
assign n33186 =  ( n39 ) & ( n32741 )  ;
assign n33187 =  ( n39 ) & ( n32743 )  ;
assign n33188 =  ( n39 ) & ( n32745 )  ;
assign n33189 =  ( n39 ) & ( n32747 )  ;
assign n33190 =  ( n39 ) & ( n32749 )  ;
assign n33191 =  ( n39 ) & ( n32751 )  ;
assign n33192 =  ( n39 ) & ( n32753 )  ;
assign n33193 =  ( n39 ) & ( n32755 )  ;
assign n33194 =  ( n39 ) & ( n32757 )  ;
assign n33195 =  ( n39 ) & ( n32759 )  ;
assign n33196 =  ( n39 ) & ( n32761 )  ;
assign n33197 =  ( n39 ) & ( n32763 )  ;
assign n33198 =  ( n39 ) & ( n32765 )  ;
assign n33199 =  ( n40 ) & ( n32735 )  ;
assign n33200 =  ( n40 ) & ( n32737 )  ;
assign n33201 =  ( n40 ) & ( n32739 )  ;
assign n33202 =  ( n40 ) & ( n32741 )  ;
assign n33203 =  ( n40 ) & ( n32743 )  ;
assign n33204 =  ( n40 ) & ( n32745 )  ;
assign n33205 =  ( n40 ) & ( n32747 )  ;
assign n33206 =  ( n40 ) & ( n32749 )  ;
assign n33207 =  ( n40 ) & ( n32751 )  ;
assign n33208 =  ( n40 ) & ( n32753 )  ;
assign n33209 =  ( n40 ) & ( n32755 )  ;
assign n33210 =  ( n40 ) & ( n32757 )  ;
assign n33211 =  ( n40 ) & ( n32759 )  ;
assign n33212 =  ( n40 ) & ( n32761 )  ;
assign n33213 =  ( n40 ) & ( n32763 )  ;
assign n33214 =  ( n40 ) & ( n32765 )  ;
assign n33215 =  ( n41 ) & ( n32735 )  ;
assign n33216 =  ( n41 ) & ( n32737 )  ;
assign n33217 =  ( n41 ) & ( n32739 )  ;
assign n33218 =  ( n41 ) & ( n32741 )  ;
assign n33219 =  ( n41 ) & ( n32743 )  ;
assign n33220 =  ( n41 ) & ( n32745 )  ;
assign n33221 =  ( n41 ) & ( n32747 )  ;
assign n33222 =  ( n41 ) & ( n32749 )  ;
assign n33223 =  ( n41 ) & ( n32751 )  ;
assign n33224 =  ( n41 ) & ( n32753 )  ;
assign n33225 =  ( n41 ) & ( n32755 )  ;
assign n33226 =  ( n41 ) & ( n32757 )  ;
assign n33227 =  ( n41 ) & ( n32759 )  ;
assign n33228 =  ( n41 ) & ( n32761 )  ;
assign n33229 =  ( n41 ) & ( n32763 )  ;
assign n33230 =  ( n41 ) & ( n32765 )  ;
assign n33231 =  ( n42 ) & ( n32735 )  ;
assign n33232 =  ( n42 ) & ( n32737 )  ;
assign n33233 =  ( n42 ) & ( n32739 )  ;
assign n33234 =  ( n42 ) & ( n32741 )  ;
assign n33235 =  ( n42 ) & ( n32743 )  ;
assign n33236 =  ( n42 ) & ( n32745 )  ;
assign n33237 =  ( n42 ) & ( n32747 )  ;
assign n33238 =  ( n42 ) & ( n32749 )  ;
assign n33239 =  ( n42 ) & ( n32751 )  ;
assign n33240 =  ( n42 ) & ( n32753 )  ;
assign n33241 =  ( n42 ) & ( n32755 )  ;
assign n33242 =  ( n42 ) & ( n32757 )  ;
assign n33243 =  ( n42 ) & ( n32759 )  ;
assign n33244 =  ( n42 ) & ( n32761 )  ;
assign n33245 =  ( n42 ) & ( n32763 )  ;
assign n33246 =  ( n42 ) & ( n32765 )  ;
assign n33247 =  ( n43 ) & ( n32735 )  ;
assign n33248 =  ( n43 ) & ( n32737 )  ;
assign n33249 =  ( n43 ) & ( n32739 )  ;
assign n33250 =  ( n43 ) & ( n32741 )  ;
assign n33251 =  ( n43 ) & ( n32743 )  ;
assign n33252 =  ( n43 ) & ( n32745 )  ;
assign n33253 =  ( n43 ) & ( n32747 )  ;
assign n33254 =  ( n43 ) & ( n32749 )  ;
assign n33255 =  ( n43 ) & ( n32751 )  ;
assign n33256 =  ( n43 ) & ( n32753 )  ;
assign n33257 =  ( n43 ) & ( n32755 )  ;
assign n33258 =  ( n43 ) & ( n32757 )  ;
assign n33259 =  ( n43 ) & ( n32759 )  ;
assign n33260 =  ( n43 ) & ( n32761 )  ;
assign n33261 =  ( n43 ) & ( n32763 )  ;
assign n33262 =  ( n43 ) & ( n32765 )  ;
assign n33263 =  ( n33262 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n33264 =  ( n33261 ) ? ( VREG_0_1 ) : ( n33263 ) ;
assign n33265 =  ( n33260 ) ? ( VREG_0_2 ) : ( n33264 ) ;
assign n33266 =  ( n33259 ) ? ( VREG_0_3 ) : ( n33265 ) ;
assign n33267 =  ( n33258 ) ? ( VREG_0_4 ) : ( n33266 ) ;
assign n33268 =  ( n33257 ) ? ( VREG_0_5 ) : ( n33267 ) ;
assign n33269 =  ( n33256 ) ? ( VREG_0_6 ) : ( n33268 ) ;
assign n33270 =  ( n33255 ) ? ( VREG_0_7 ) : ( n33269 ) ;
assign n33271 =  ( n33254 ) ? ( VREG_0_8 ) : ( n33270 ) ;
assign n33272 =  ( n33253 ) ? ( VREG_0_9 ) : ( n33271 ) ;
assign n33273 =  ( n33252 ) ? ( VREG_0_10 ) : ( n33272 ) ;
assign n33274 =  ( n33251 ) ? ( VREG_0_11 ) : ( n33273 ) ;
assign n33275 =  ( n33250 ) ? ( VREG_0_12 ) : ( n33274 ) ;
assign n33276 =  ( n33249 ) ? ( VREG_0_13 ) : ( n33275 ) ;
assign n33277 =  ( n33248 ) ? ( VREG_0_14 ) : ( n33276 ) ;
assign n33278 =  ( n33247 ) ? ( VREG_0_15 ) : ( n33277 ) ;
assign n33279 =  ( n33246 ) ? ( VREG_1_0 ) : ( n33278 ) ;
assign n33280 =  ( n33245 ) ? ( VREG_1_1 ) : ( n33279 ) ;
assign n33281 =  ( n33244 ) ? ( VREG_1_2 ) : ( n33280 ) ;
assign n33282 =  ( n33243 ) ? ( VREG_1_3 ) : ( n33281 ) ;
assign n33283 =  ( n33242 ) ? ( VREG_1_4 ) : ( n33282 ) ;
assign n33284 =  ( n33241 ) ? ( VREG_1_5 ) : ( n33283 ) ;
assign n33285 =  ( n33240 ) ? ( VREG_1_6 ) : ( n33284 ) ;
assign n33286 =  ( n33239 ) ? ( VREG_1_7 ) : ( n33285 ) ;
assign n33287 =  ( n33238 ) ? ( VREG_1_8 ) : ( n33286 ) ;
assign n33288 =  ( n33237 ) ? ( VREG_1_9 ) : ( n33287 ) ;
assign n33289 =  ( n33236 ) ? ( VREG_1_10 ) : ( n33288 ) ;
assign n33290 =  ( n33235 ) ? ( VREG_1_11 ) : ( n33289 ) ;
assign n33291 =  ( n33234 ) ? ( VREG_1_12 ) : ( n33290 ) ;
assign n33292 =  ( n33233 ) ? ( VREG_1_13 ) : ( n33291 ) ;
assign n33293 =  ( n33232 ) ? ( VREG_1_14 ) : ( n33292 ) ;
assign n33294 =  ( n33231 ) ? ( VREG_1_15 ) : ( n33293 ) ;
assign n33295 =  ( n33230 ) ? ( VREG_2_0 ) : ( n33294 ) ;
assign n33296 =  ( n33229 ) ? ( VREG_2_1 ) : ( n33295 ) ;
assign n33297 =  ( n33228 ) ? ( VREG_2_2 ) : ( n33296 ) ;
assign n33298 =  ( n33227 ) ? ( VREG_2_3 ) : ( n33297 ) ;
assign n33299 =  ( n33226 ) ? ( VREG_2_4 ) : ( n33298 ) ;
assign n33300 =  ( n33225 ) ? ( VREG_2_5 ) : ( n33299 ) ;
assign n33301 =  ( n33224 ) ? ( VREG_2_6 ) : ( n33300 ) ;
assign n33302 =  ( n33223 ) ? ( VREG_2_7 ) : ( n33301 ) ;
assign n33303 =  ( n33222 ) ? ( VREG_2_8 ) : ( n33302 ) ;
assign n33304 =  ( n33221 ) ? ( VREG_2_9 ) : ( n33303 ) ;
assign n33305 =  ( n33220 ) ? ( VREG_2_10 ) : ( n33304 ) ;
assign n33306 =  ( n33219 ) ? ( VREG_2_11 ) : ( n33305 ) ;
assign n33307 =  ( n33218 ) ? ( VREG_2_12 ) : ( n33306 ) ;
assign n33308 =  ( n33217 ) ? ( VREG_2_13 ) : ( n33307 ) ;
assign n33309 =  ( n33216 ) ? ( VREG_2_14 ) : ( n33308 ) ;
assign n33310 =  ( n33215 ) ? ( VREG_2_15 ) : ( n33309 ) ;
assign n33311 =  ( n33214 ) ? ( VREG_3_0 ) : ( n33310 ) ;
assign n33312 =  ( n33213 ) ? ( VREG_3_1 ) : ( n33311 ) ;
assign n33313 =  ( n33212 ) ? ( VREG_3_2 ) : ( n33312 ) ;
assign n33314 =  ( n33211 ) ? ( VREG_3_3 ) : ( n33313 ) ;
assign n33315 =  ( n33210 ) ? ( VREG_3_4 ) : ( n33314 ) ;
assign n33316 =  ( n33209 ) ? ( VREG_3_5 ) : ( n33315 ) ;
assign n33317 =  ( n33208 ) ? ( VREG_3_6 ) : ( n33316 ) ;
assign n33318 =  ( n33207 ) ? ( VREG_3_7 ) : ( n33317 ) ;
assign n33319 =  ( n33206 ) ? ( VREG_3_8 ) : ( n33318 ) ;
assign n33320 =  ( n33205 ) ? ( VREG_3_9 ) : ( n33319 ) ;
assign n33321 =  ( n33204 ) ? ( VREG_3_10 ) : ( n33320 ) ;
assign n33322 =  ( n33203 ) ? ( VREG_3_11 ) : ( n33321 ) ;
assign n33323 =  ( n33202 ) ? ( VREG_3_12 ) : ( n33322 ) ;
assign n33324 =  ( n33201 ) ? ( VREG_3_13 ) : ( n33323 ) ;
assign n33325 =  ( n33200 ) ? ( VREG_3_14 ) : ( n33324 ) ;
assign n33326 =  ( n33199 ) ? ( VREG_3_15 ) : ( n33325 ) ;
assign n33327 =  ( n33198 ) ? ( VREG_4_0 ) : ( n33326 ) ;
assign n33328 =  ( n33197 ) ? ( VREG_4_1 ) : ( n33327 ) ;
assign n33329 =  ( n33196 ) ? ( VREG_4_2 ) : ( n33328 ) ;
assign n33330 =  ( n33195 ) ? ( VREG_4_3 ) : ( n33329 ) ;
assign n33331 =  ( n33194 ) ? ( VREG_4_4 ) : ( n33330 ) ;
assign n33332 =  ( n33193 ) ? ( VREG_4_5 ) : ( n33331 ) ;
assign n33333 =  ( n33192 ) ? ( VREG_4_6 ) : ( n33332 ) ;
assign n33334 =  ( n33191 ) ? ( VREG_4_7 ) : ( n33333 ) ;
assign n33335 =  ( n33190 ) ? ( VREG_4_8 ) : ( n33334 ) ;
assign n33336 =  ( n33189 ) ? ( VREG_4_9 ) : ( n33335 ) ;
assign n33337 =  ( n33188 ) ? ( VREG_4_10 ) : ( n33336 ) ;
assign n33338 =  ( n33187 ) ? ( VREG_4_11 ) : ( n33337 ) ;
assign n33339 =  ( n33186 ) ? ( VREG_4_12 ) : ( n33338 ) ;
assign n33340 =  ( n33185 ) ? ( VREG_4_13 ) : ( n33339 ) ;
assign n33341 =  ( n33184 ) ? ( VREG_4_14 ) : ( n33340 ) ;
assign n33342 =  ( n33183 ) ? ( VREG_4_15 ) : ( n33341 ) ;
assign n33343 =  ( n33182 ) ? ( VREG_5_0 ) : ( n33342 ) ;
assign n33344 =  ( n33181 ) ? ( VREG_5_1 ) : ( n33343 ) ;
assign n33345 =  ( n33180 ) ? ( VREG_5_2 ) : ( n33344 ) ;
assign n33346 =  ( n33179 ) ? ( VREG_5_3 ) : ( n33345 ) ;
assign n33347 =  ( n33178 ) ? ( VREG_5_4 ) : ( n33346 ) ;
assign n33348 =  ( n33177 ) ? ( VREG_5_5 ) : ( n33347 ) ;
assign n33349 =  ( n33176 ) ? ( VREG_5_6 ) : ( n33348 ) ;
assign n33350 =  ( n33175 ) ? ( VREG_5_7 ) : ( n33349 ) ;
assign n33351 =  ( n33174 ) ? ( VREG_5_8 ) : ( n33350 ) ;
assign n33352 =  ( n33173 ) ? ( VREG_5_9 ) : ( n33351 ) ;
assign n33353 =  ( n33172 ) ? ( VREG_5_10 ) : ( n33352 ) ;
assign n33354 =  ( n33171 ) ? ( VREG_5_11 ) : ( n33353 ) ;
assign n33355 =  ( n33170 ) ? ( VREG_5_12 ) : ( n33354 ) ;
assign n33356 =  ( n33169 ) ? ( VREG_5_13 ) : ( n33355 ) ;
assign n33357 =  ( n33168 ) ? ( VREG_5_14 ) : ( n33356 ) ;
assign n33358 =  ( n33167 ) ? ( VREG_5_15 ) : ( n33357 ) ;
assign n33359 =  ( n33166 ) ? ( VREG_6_0 ) : ( n33358 ) ;
assign n33360 =  ( n33165 ) ? ( VREG_6_1 ) : ( n33359 ) ;
assign n33361 =  ( n33164 ) ? ( VREG_6_2 ) : ( n33360 ) ;
assign n33362 =  ( n33163 ) ? ( VREG_6_3 ) : ( n33361 ) ;
assign n33363 =  ( n33162 ) ? ( VREG_6_4 ) : ( n33362 ) ;
assign n33364 =  ( n33161 ) ? ( VREG_6_5 ) : ( n33363 ) ;
assign n33365 =  ( n33160 ) ? ( VREG_6_6 ) : ( n33364 ) ;
assign n33366 =  ( n33159 ) ? ( VREG_6_7 ) : ( n33365 ) ;
assign n33367 =  ( n33158 ) ? ( VREG_6_8 ) : ( n33366 ) ;
assign n33368 =  ( n33157 ) ? ( VREG_6_9 ) : ( n33367 ) ;
assign n33369 =  ( n33156 ) ? ( VREG_6_10 ) : ( n33368 ) ;
assign n33370 =  ( n33155 ) ? ( VREG_6_11 ) : ( n33369 ) ;
assign n33371 =  ( n33154 ) ? ( VREG_6_12 ) : ( n33370 ) ;
assign n33372 =  ( n33153 ) ? ( VREG_6_13 ) : ( n33371 ) ;
assign n33373 =  ( n33152 ) ? ( VREG_6_14 ) : ( n33372 ) ;
assign n33374 =  ( n33151 ) ? ( VREG_6_15 ) : ( n33373 ) ;
assign n33375 =  ( n33150 ) ? ( VREG_7_0 ) : ( n33374 ) ;
assign n33376 =  ( n33149 ) ? ( VREG_7_1 ) : ( n33375 ) ;
assign n33377 =  ( n33148 ) ? ( VREG_7_2 ) : ( n33376 ) ;
assign n33378 =  ( n33147 ) ? ( VREG_7_3 ) : ( n33377 ) ;
assign n33379 =  ( n33146 ) ? ( VREG_7_4 ) : ( n33378 ) ;
assign n33380 =  ( n33145 ) ? ( VREG_7_5 ) : ( n33379 ) ;
assign n33381 =  ( n33144 ) ? ( VREG_7_6 ) : ( n33380 ) ;
assign n33382 =  ( n33143 ) ? ( VREG_7_7 ) : ( n33381 ) ;
assign n33383 =  ( n33142 ) ? ( VREG_7_8 ) : ( n33382 ) ;
assign n33384 =  ( n33141 ) ? ( VREG_7_9 ) : ( n33383 ) ;
assign n33385 =  ( n33140 ) ? ( VREG_7_10 ) : ( n33384 ) ;
assign n33386 =  ( n33139 ) ? ( VREG_7_11 ) : ( n33385 ) ;
assign n33387 =  ( n33138 ) ? ( VREG_7_12 ) : ( n33386 ) ;
assign n33388 =  ( n33137 ) ? ( VREG_7_13 ) : ( n33387 ) ;
assign n33389 =  ( n33136 ) ? ( VREG_7_14 ) : ( n33388 ) ;
assign n33390 =  ( n33135 ) ? ( VREG_7_15 ) : ( n33389 ) ;
assign n33391 =  ( n33134 ) ? ( VREG_8_0 ) : ( n33390 ) ;
assign n33392 =  ( n33133 ) ? ( VREG_8_1 ) : ( n33391 ) ;
assign n33393 =  ( n33132 ) ? ( VREG_8_2 ) : ( n33392 ) ;
assign n33394 =  ( n33131 ) ? ( VREG_8_3 ) : ( n33393 ) ;
assign n33395 =  ( n33130 ) ? ( VREG_8_4 ) : ( n33394 ) ;
assign n33396 =  ( n33129 ) ? ( VREG_8_5 ) : ( n33395 ) ;
assign n33397 =  ( n33128 ) ? ( VREG_8_6 ) : ( n33396 ) ;
assign n33398 =  ( n33127 ) ? ( VREG_8_7 ) : ( n33397 ) ;
assign n33399 =  ( n33126 ) ? ( VREG_8_8 ) : ( n33398 ) ;
assign n33400 =  ( n33125 ) ? ( VREG_8_9 ) : ( n33399 ) ;
assign n33401 =  ( n33124 ) ? ( VREG_8_10 ) : ( n33400 ) ;
assign n33402 =  ( n33123 ) ? ( VREG_8_11 ) : ( n33401 ) ;
assign n33403 =  ( n33122 ) ? ( VREG_8_12 ) : ( n33402 ) ;
assign n33404 =  ( n33121 ) ? ( VREG_8_13 ) : ( n33403 ) ;
assign n33405 =  ( n33120 ) ? ( VREG_8_14 ) : ( n33404 ) ;
assign n33406 =  ( n33119 ) ? ( VREG_8_15 ) : ( n33405 ) ;
assign n33407 =  ( n33118 ) ? ( VREG_9_0 ) : ( n33406 ) ;
assign n33408 =  ( n33117 ) ? ( VREG_9_1 ) : ( n33407 ) ;
assign n33409 =  ( n33116 ) ? ( VREG_9_2 ) : ( n33408 ) ;
assign n33410 =  ( n33115 ) ? ( VREG_9_3 ) : ( n33409 ) ;
assign n33411 =  ( n33114 ) ? ( VREG_9_4 ) : ( n33410 ) ;
assign n33412 =  ( n33113 ) ? ( VREG_9_5 ) : ( n33411 ) ;
assign n33413 =  ( n33112 ) ? ( VREG_9_6 ) : ( n33412 ) ;
assign n33414 =  ( n33111 ) ? ( VREG_9_7 ) : ( n33413 ) ;
assign n33415 =  ( n33110 ) ? ( VREG_9_8 ) : ( n33414 ) ;
assign n33416 =  ( n33109 ) ? ( VREG_9_9 ) : ( n33415 ) ;
assign n33417 =  ( n33108 ) ? ( VREG_9_10 ) : ( n33416 ) ;
assign n33418 =  ( n33107 ) ? ( VREG_9_11 ) : ( n33417 ) ;
assign n33419 =  ( n33106 ) ? ( VREG_9_12 ) : ( n33418 ) ;
assign n33420 =  ( n33105 ) ? ( VREG_9_13 ) : ( n33419 ) ;
assign n33421 =  ( n33104 ) ? ( VREG_9_14 ) : ( n33420 ) ;
assign n33422 =  ( n33103 ) ? ( VREG_9_15 ) : ( n33421 ) ;
assign n33423 =  ( n33102 ) ? ( VREG_10_0 ) : ( n33422 ) ;
assign n33424 =  ( n33101 ) ? ( VREG_10_1 ) : ( n33423 ) ;
assign n33425 =  ( n33100 ) ? ( VREG_10_2 ) : ( n33424 ) ;
assign n33426 =  ( n33099 ) ? ( VREG_10_3 ) : ( n33425 ) ;
assign n33427 =  ( n33098 ) ? ( VREG_10_4 ) : ( n33426 ) ;
assign n33428 =  ( n33097 ) ? ( VREG_10_5 ) : ( n33427 ) ;
assign n33429 =  ( n33096 ) ? ( VREG_10_6 ) : ( n33428 ) ;
assign n33430 =  ( n33095 ) ? ( VREG_10_7 ) : ( n33429 ) ;
assign n33431 =  ( n33094 ) ? ( VREG_10_8 ) : ( n33430 ) ;
assign n33432 =  ( n33093 ) ? ( VREG_10_9 ) : ( n33431 ) ;
assign n33433 =  ( n33092 ) ? ( VREG_10_10 ) : ( n33432 ) ;
assign n33434 =  ( n33091 ) ? ( VREG_10_11 ) : ( n33433 ) ;
assign n33435 =  ( n33090 ) ? ( VREG_10_12 ) : ( n33434 ) ;
assign n33436 =  ( n33089 ) ? ( VREG_10_13 ) : ( n33435 ) ;
assign n33437 =  ( n33088 ) ? ( VREG_10_14 ) : ( n33436 ) ;
assign n33438 =  ( n33087 ) ? ( VREG_10_15 ) : ( n33437 ) ;
assign n33439 =  ( n33086 ) ? ( VREG_11_0 ) : ( n33438 ) ;
assign n33440 =  ( n33085 ) ? ( VREG_11_1 ) : ( n33439 ) ;
assign n33441 =  ( n33084 ) ? ( VREG_11_2 ) : ( n33440 ) ;
assign n33442 =  ( n33083 ) ? ( VREG_11_3 ) : ( n33441 ) ;
assign n33443 =  ( n33082 ) ? ( VREG_11_4 ) : ( n33442 ) ;
assign n33444 =  ( n33081 ) ? ( VREG_11_5 ) : ( n33443 ) ;
assign n33445 =  ( n33080 ) ? ( VREG_11_6 ) : ( n33444 ) ;
assign n33446 =  ( n33079 ) ? ( VREG_11_7 ) : ( n33445 ) ;
assign n33447 =  ( n33078 ) ? ( VREG_11_8 ) : ( n33446 ) ;
assign n33448 =  ( n33077 ) ? ( VREG_11_9 ) : ( n33447 ) ;
assign n33449 =  ( n33076 ) ? ( VREG_11_10 ) : ( n33448 ) ;
assign n33450 =  ( n33075 ) ? ( VREG_11_11 ) : ( n33449 ) ;
assign n33451 =  ( n33074 ) ? ( VREG_11_12 ) : ( n33450 ) ;
assign n33452 =  ( n33073 ) ? ( VREG_11_13 ) : ( n33451 ) ;
assign n33453 =  ( n33072 ) ? ( VREG_11_14 ) : ( n33452 ) ;
assign n33454 =  ( n33071 ) ? ( VREG_11_15 ) : ( n33453 ) ;
assign n33455 =  ( n33070 ) ? ( VREG_12_0 ) : ( n33454 ) ;
assign n33456 =  ( n33069 ) ? ( VREG_12_1 ) : ( n33455 ) ;
assign n33457 =  ( n33068 ) ? ( VREG_12_2 ) : ( n33456 ) ;
assign n33458 =  ( n33067 ) ? ( VREG_12_3 ) : ( n33457 ) ;
assign n33459 =  ( n33066 ) ? ( VREG_12_4 ) : ( n33458 ) ;
assign n33460 =  ( n33065 ) ? ( VREG_12_5 ) : ( n33459 ) ;
assign n33461 =  ( n33064 ) ? ( VREG_12_6 ) : ( n33460 ) ;
assign n33462 =  ( n33063 ) ? ( VREG_12_7 ) : ( n33461 ) ;
assign n33463 =  ( n33062 ) ? ( VREG_12_8 ) : ( n33462 ) ;
assign n33464 =  ( n33061 ) ? ( VREG_12_9 ) : ( n33463 ) ;
assign n33465 =  ( n33060 ) ? ( VREG_12_10 ) : ( n33464 ) ;
assign n33466 =  ( n33059 ) ? ( VREG_12_11 ) : ( n33465 ) ;
assign n33467 =  ( n33058 ) ? ( VREG_12_12 ) : ( n33466 ) ;
assign n33468 =  ( n33057 ) ? ( VREG_12_13 ) : ( n33467 ) ;
assign n33469 =  ( n33056 ) ? ( VREG_12_14 ) : ( n33468 ) ;
assign n33470 =  ( n33055 ) ? ( VREG_12_15 ) : ( n33469 ) ;
assign n33471 =  ( n33054 ) ? ( VREG_13_0 ) : ( n33470 ) ;
assign n33472 =  ( n33053 ) ? ( VREG_13_1 ) : ( n33471 ) ;
assign n33473 =  ( n33052 ) ? ( VREG_13_2 ) : ( n33472 ) ;
assign n33474 =  ( n33051 ) ? ( VREG_13_3 ) : ( n33473 ) ;
assign n33475 =  ( n33050 ) ? ( VREG_13_4 ) : ( n33474 ) ;
assign n33476 =  ( n33049 ) ? ( VREG_13_5 ) : ( n33475 ) ;
assign n33477 =  ( n33048 ) ? ( VREG_13_6 ) : ( n33476 ) ;
assign n33478 =  ( n33047 ) ? ( VREG_13_7 ) : ( n33477 ) ;
assign n33479 =  ( n33046 ) ? ( VREG_13_8 ) : ( n33478 ) ;
assign n33480 =  ( n33045 ) ? ( VREG_13_9 ) : ( n33479 ) ;
assign n33481 =  ( n33044 ) ? ( VREG_13_10 ) : ( n33480 ) ;
assign n33482 =  ( n33043 ) ? ( VREG_13_11 ) : ( n33481 ) ;
assign n33483 =  ( n33042 ) ? ( VREG_13_12 ) : ( n33482 ) ;
assign n33484 =  ( n33041 ) ? ( VREG_13_13 ) : ( n33483 ) ;
assign n33485 =  ( n33040 ) ? ( VREG_13_14 ) : ( n33484 ) ;
assign n33486 =  ( n33039 ) ? ( VREG_13_15 ) : ( n33485 ) ;
assign n33487 =  ( n33038 ) ? ( VREG_14_0 ) : ( n33486 ) ;
assign n33488 =  ( n33037 ) ? ( VREG_14_1 ) : ( n33487 ) ;
assign n33489 =  ( n33036 ) ? ( VREG_14_2 ) : ( n33488 ) ;
assign n33490 =  ( n33035 ) ? ( VREG_14_3 ) : ( n33489 ) ;
assign n33491 =  ( n33034 ) ? ( VREG_14_4 ) : ( n33490 ) ;
assign n33492 =  ( n33033 ) ? ( VREG_14_5 ) : ( n33491 ) ;
assign n33493 =  ( n33032 ) ? ( VREG_14_6 ) : ( n33492 ) ;
assign n33494 =  ( n33031 ) ? ( VREG_14_7 ) : ( n33493 ) ;
assign n33495 =  ( n33030 ) ? ( VREG_14_8 ) : ( n33494 ) ;
assign n33496 =  ( n33029 ) ? ( VREG_14_9 ) : ( n33495 ) ;
assign n33497 =  ( n33028 ) ? ( VREG_14_10 ) : ( n33496 ) ;
assign n33498 =  ( n33027 ) ? ( VREG_14_11 ) : ( n33497 ) ;
assign n33499 =  ( n33026 ) ? ( VREG_14_12 ) : ( n33498 ) ;
assign n33500 =  ( n33025 ) ? ( VREG_14_13 ) : ( n33499 ) ;
assign n33501 =  ( n33024 ) ? ( VREG_14_14 ) : ( n33500 ) ;
assign n33502 =  ( n33023 ) ? ( VREG_14_15 ) : ( n33501 ) ;
assign n33503 =  ( n33022 ) ? ( VREG_15_0 ) : ( n33502 ) ;
assign n33504 =  ( n33021 ) ? ( VREG_15_1 ) : ( n33503 ) ;
assign n33505 =  ( n33020 ) ? ( VREG_15_2 ) : ( n33504 ) ;
assign n33506 =  ( n33019 ) ? ( VREG_15_3 ) : ( n33505 ) ;
assign n33507 =  ( n33018 ) ? ( VREG_15_4 ) : ( n33506 ) ;
assign n33508 =  ( n33017 ) ? ( VREG_15_5 ) : ( n33507 ) ;
assign n33509 =  ( n33016 ) ? ( VREG_15_6 ) : ( n33508 ) ;
assign n33510 =  ( n33015 ) ? ( VREG_15_7 ) : ( n33509 ) ;
assign n33511 =  ( n33014 ) ? ( VREG_15_8 ) : ( n33510 ) ;
assign n33512 =  ( n33013 ) ? ( VREG_15_9 ) : ( n33511 ) ;
assign n33513 =  ( n33012 ) ? ( VREG_15_10 ) : ( n33512 ) ;
assign n33514 =  ( n33011 ) ? ( VREG_15_11 ) : ( n33513 ) ;
assign n33515 =  ( n33010 ) ? ( VREG_15_12 ) : ( n33514 ) ;
assign n33516 =  ( n33009 ) ? ( VREG_15_13 ) : ( n33515 ) ;
assign n33517 =  ( n33008 ) ? ( VREG_15_14 ) : ( n33516 ) ;
assign n33518 =  ( n33007 ) ? ( VREG_15_15 ) : ( n33517 ) ;
assign n33519 =  ( n33006 ) ? ( VREG_16_0 ) : ( n33518 ) ;
assign n33520 =  ( n33005 ) ? ( VREG_16_1 ) : ( n33519 ) ;
assign n33521 =  ( n33004 ) ? ( VREG_16_2 ) : ( n33520 ) ;
assign n33522 =  ( n33003 ) ? ( VREG_16_3 ) : ( n33521 ) ;
assign n33523 =  ( n33002 ) ? ( VREG_16_4 ) : ( n33522 ) ;
assign n33524 =  ( n33001 ) ? ( VREG_16_5 ) : ( n33523 ) ;
assign n33525 =  ( n33000 ) ? ( VREG_16_6 ) : ( n33524 ) ;
assign n33526 =  ( n32999 ) ? ( VREG_16_7 ) : ( n33525 ) ;
assign n33527 =  ( n32998 ) ? ( VREG_16_8 ) : ( n33526 ) ;
assign n33528 =  ( n32997 ) ? ( VREG_16_9 ) : ( n33527 ) ;
assign n33529 =  ( n32996 ) ? ( VREG_16_10 ) : ( n33528 ) ;
assign n33530 =  ( n32995 ) ? ( VREG_16_11 ) : ( n33529 ) ;
assign n33531 =  ( n32994 ) ? ( VREG_16_12 ) : ( n33530 ) ;
assign n33532 =  ( n32993 ) ? ( VREG_16_13 ) : ( n33531 ) ;
assign n33533 =  ( n32992 ) ? ( VREG_16_14 ) : ( n33532 ) ;
assign n33534 =  ( n32991 ) ? ( VREG_16_15 ) : ( n33533 ) ;
assign n33535 =  ( n32990 ) ? ( VREG_17_0 ) : ( n33534 ) ;
assign n33536 =  ( n32989 ) ? ( VREG_17_1 ) : ( n33535 ) ;
assign n33537 =  ( n32988 ) ? ( VREG_17_2 ) : ( n33536 ) ;
assign n33538 =  ( n32987 ) ? ( VREG_17_3 ) : ( n33537 ) ;
assign n33539 =  ( n32986 ) ? ( VREG_17_4 ) : ( n33538 ) ;
assign n33540 =  ( n32985 ) ? ( VREG_17_5 ) : ( n33539 ) ;
assign n33541 =  ( n32984 ) ? ( VREG_17_6 ) : ( n33540 ) ;
assign n33542 =  ( n32983 ) ? ( VREG_17_7 ) : ( n33541 ) ;
assign n33543 =  ( n32982 ) ? ( VREG_17_8 ) : ( n33542 ) ;
assign n33544 =  ( n32981 ) ? ( VREG_17_9 ) : ( n33543 ) ;
assign n33545 =  ( n32980 ) ? ( VREG_17_10 ) : ( n33544 ) ;
assign n33546 =  ( n32979 ) ? ( VREG_17_11 ) : ( n33545 ) ;
assign n33547 =  ( n32978 ) ? ( VREG_17_12 ) : ( n33546 ) ;
assign n33548 =  ( n32977 ) ? ( VREG_17_13 ) : ( n33547 ) ;
assign n33549 =  ( n32976 ) ? ( VREG_17_14 ) : ( n33548 ) ;
assign n33550 =  ( n32975 ) ? ( VREG_17_15 ) : ( n33549 ) ;
assign n33551 =  ( n32974 ) ? ( VREG_18_0 ) : ( n33550 ) ;
assign n33552 =  ( n32973 ) ? ( VREG_18_1 ) : ( n33551 ) ;
assign n33553 =  ( n32972 ) ? ( VREG_18_2 ) : ( n33552 ) ;
assign n33554 =  ( n32971 ) ? ( VREG_18_3 ) : ( n33553 ) ;
assign n33555 =  ( n32970 ) ? ( VREG_18_4 ) : ( n33554 ) ;
assign n33556 =  ( n32969 ) ? ( VREG_18_5 ) : ( n33555 ) ;
assign n33557 =  ( n32968 ) ? ( VREG_18_6 ) : ( n33556 ) ;
assign n33558 =  ( n32967 ) ? ( VREG_18_7 ) : ( n33557 ) ;
assign n33559 =  ( n32966 ) ? ( VREG_18_8 ) : ( n33558 ) ;
assign n33560 =  ( n32965 ) ? ( VREG_18_9 ) : ( n33559 ) ;
assign n33561 =  ( n32964 ) ? ( VREG_18_10 ) : ( n33560 ) ;
assign n33562 =  ( n32963 ) ? ( VREG_18_11 ) : ( n33561 ) ;
assign n33563 =  ( n32962 ) ? ( VREG_18_12 ) : ( n33562 ) ;
assign n33564 =  ( n32961 ) ? ( VREG_18_13 ) : ( n33563 ) ;
assign n33565 =  ( n32960 ) ? ( VREG_18_14 ) : ( n33564 ) ;
assign n33566 =  ( n32959 ) ? ( VREG_18_15 ) : ( n33565 ) ;
assign n33567 =  ( n32958 ) ? ( VREG_19_0 ) : ( n33566 ) ;
assign n33568 =  ( n32957 ) ? ( VREG_19_1 ) : ( n33567 ) ;
assign n33569 =  ( n32956 ) ? ( VREG_19_2 ) : ( n33568 ) ;
assign n33570 =  ( n32955 ) ? ( VREG_19_3 ) : ( n33569 ) ;
assign n33571 =  ( n32954 ) ? ( VREG_19_4 ) : ( n33570 ) ;
assign n33572 =  ( n32953 ) ? ( VREG_19_5 ) : ( n33571 ) ;
assign n33573 =  ( n32952 ) ? ( VREG_19_6 ) : ( n33572 ) ;
assign n33574 =  ( n32951 ) ? ( VREG_19_7 ) : ( n33573 ) ;
assign n33575 =  ( n32950 ) ? ( VREG_19_8 ) : ( n33574 ) ;
assign n33576 =  ( n32949 ) ? ( VREG_19_9 ) : ( n33575 ) ;
assign n33577 =  ( n32948 ) ? ( VREG_19_10 ) : ( n33576 ) ;
assign n33578 =  ( n32947 ) ? ( VREG_19_11 ) : ( n33577 ) ;
assign n33579 =  ( n32946 ) ? ( VREG_19_12 ) : ( n33578 ) ;
assign n33580 =  ( n32945 ) ? ( VREG_19_13 ) : ( n33579 ) ;
assign n33581 =  ( n32944 ) ? ( VREG_19_14 ) : ( n33580 ) ;
assign n33582 =  ( n32943 ) ? ( VREG_19_15 ) : ( n33581 ) ;
assign n33583 =  ( n32942 ) ? ( VREG_20_0 ) : ( n33582 ) ;
assign n33584 =  ( n32941 ) ? ( VREG_20_1 ) : ( n33583 ) ;
assign n33585 =  ( n32940 ) ? ( VREG_20_2 ) : ( n33584 ) ;
assign n33586 =  ( n32939 ) ? ( VREG_20_3 ) : ( n33585 ) ;
assign n33587 =  ( n32938 ) ? ( VREG_20_4 ) : ( n33586 ) ;
assign n33588 =  ( n32937 ) ? ( VREG_20_5 ) : ( n33587 ) ;
assign n33589 =  ( n32936 ) ? ( VREG_20_6 ) : ( n33588 ) ;
assign n33590 =  ( n32935 ) ? ( VREG_20_7 ) : ( n33589 ) ;
assign n33591 =  ( n32934 ) ? ( VREG_20_8 ) : ( n33590 ) ;
assign n33592 =  ( n32933 ) ? ( VREG_20_9 ) : ( n33591 ) ;
assign n33593 =  ( n32932 ) ? ( VREG_20_10 ) : ( n33592 ) ;
assign n33594 =  ( n32931 ) ? ( VREG_20_11 ) : ( n33593 ) ;
assign n33595 =  ( n32930 ) ? ( VREG_20_12 ) : ( n33594 ) ;
assign n33596 =  ( n32929 ) ? ( VREG_20_13 ) : ( n33595 ) ;
assign n33597 =  ( n32928 ) ? ( VREG_20_14 ) : ( n33596 ) ;
assign n33598 =  ( n32927 ) ? ( VREG_20_15 ) : ( n33597 ) ;
assign n33599 =  ( n32926 ) ? ( VREG_21_0 ) : ( n33598 ) ;
assign n33600 =  ( n32925 ) ? ( VREG_21_1 ) : ( n33599 ) ;
assign n33601 =  ( n32924 ) ? ( VREG_21_2 ) : ( n33600 ) ;
assign n33602 =  ( n32923 ) ? ( VREG_21_3 ) : ( n33601 ) ;
assign n33603 =  ( n32922 ) ? ( VREG_21_4 ) : ( n33602 ) ;
assign n33604 =  ( n32921 ) ? ( VREG_21_5 ) : ( n33603 ) ;
assign n33605 =  ( n32920 ) ? ( VREG_21_6 ) : ( n33604 ) ;
assign n33606 =  ( n32919 ) ? ( VREG_21_7 ) : ( n33605 ) ;
assign n33607 =  ( n32918 ) ? ( VREG_21_8 ) : ( n33606 ) ;
assign n33608 =  ( n32917 ) ? ( VREG_21_9 ) : ( n33607 ) ;
assign n33609 =  ( n32916 ) ? ( VREG_21_10 ) : ( n33608 ) ;
assign n33610 =  ( n32915 ) ? ( VREG_21_11 ) : ( n33609 ) ;
assign n33611 =  ( n32914 ) ? ( VREG_21_12 ) : ( n33610 ) ;
assign n33612 =  ( n32913 ) ? ( VREG_21_13 ) : ( n33611 ) ;
assign n33613 =  ( n32912 ) ? ( VREG_21_14 ) : ( n33612 ) ;
assign n33614 =  ( n32911 ) ? ( VREG_21_15 ) : ( n33613 ) ;
assign n33615 =  ( n32910 ) ? ( VREG_22_0 ) : ( n33614 ) ;
assign n33616 =  ( n32909 ) ? ( VREG_22_1 ) : ( n33615 ) ;
assign n33617 =  ( n32908 ) ? ( VREG_22_2 ) : ( n33616 ) ;
assign n33618 =  ( n32907 ) ? ( VREG_22_3 ) : ( n33617 ) ;
assign n33619 =  ( n32906 ) ? ( VREG_22_4 ) : ( n33618 ) ;
assign n33620 =  ( n32905 ) ? ( VREG_22_5 ) : ( n33619 ) ;
assign n33621 =  ( n32904 ) ? ( VREG_22_6 ) : ( n33620 ) ;
assign n33622 =  ( n32903 ) ? ( VREG_22_7 ) : ( n33621 ) ;
assign n33623 =  ( n32902 ) ? ( VREG_22_8 ) : ( n33622 ) ;
assign n33624 =  ( n32901 ) ? ( VREG_22_9 ) : ( n33623 ) ;
assign n33625 =  ( n32900 ) ? ( VREG_22_10 ) : ( n33624 ) ;
assign n33626 =  ( n32899 ) ? ( VREG_22_11 ) : ( n33625 ) ;
assign n33627 =  ( n32898 ) ? ( VREG_22_12 ) : ( n33626 ) ;
assign n33628 =  ( n32897 ) ? ( VREG_22_13 ) : ( n33627 ) ;
assign n33629 =  ( n32896 ) ? ( VREG_22_14 ) : ( n33628 ) ;
assign n33630 =  ( n32895 ) ? ( VREG_22_15 ) : ( n33629 ) ;
assign n33631 =  ( n32894 ) ? ( VREG_23_0 ) : ( n33630 ) ;
assign n33632 =  ( n32893 ) ? ( VREG_23_1 ) : ( n33631 ) ;
assign n33633 =  ( n32892 ) ? ( VREG_23_2 ) : ( n33632 ) ;
assign n33634 =  ( n32891 ) ? ( VREG_23_3 ) : ( n33633 ) ;
assign n33635 =  ( n32890 ) ? ( VREG_23_4 ) : ( n33634 ) ;
assign n33636 =  ( n32889 ) ? ( VREG_23_5 ) : ( n33635 ) ;
assign n33637 =  ( n32888 ) ? ( VREG_23_6 ) : ( n33636 ) ;
assign n33638 =  ( n32887 ) ? ( VREG_23_7 ) : ( n33637 ) ;
assign n33639 =  ( n32886 ) ? ( VREG_23_8 ) : ( n33638 ) ;
assign n33640 =  ( n32885 ) ? ( VREG_23_9 ) : ( n33639 ) ;
assign n33641 =  ( n32884 ) ? ( VREG_23_10 ) : ( n33640 ) ;
assign n33642 =  ( n32883 ) ? ( VREG_23_11 ) : ( n33641 ) ;
assign n33643 =  ( n32882 ) ? ( VREG_23_12 ) : ( n33642 ) ;
assign n33644 =  ( n32881 ) ? ( VREG_23_13 ) : ( n33643 ) ;
assign n33645 =  ( n32880 ) ? ( VREG_23_14 ) : ( n33644 ) ;
assign n33646 =  ( n32879 ) ? ( VREG_23_15 ) : ( n33645 ) ;
assign n33647 =  ( n32878 ) ? ( VREG_24_0 ) : ( n33646 ) ;
assign n33648 =  ( n32877 ) ? ( VREG_24_1 ) : ( n33647 ) ;
assign n33649 =  ( n32876 ) ? ( VREG_24_2 ) : ( n33648 ) ;
assign n33650 =  ( n32875 ) ? ( VREG_24_3 ) : ( n33649 ) ;
assign n33651 =  ( n32874 ) ? ( VREG_24_4 ) : ( n33650 ) ;
assign n33652 =  ( n32873 ) ? ( VREG_24_5 ) : ( n33651 ) ;
assign n33653 =  ( n32872 ) ? ( VREG_24_6 ) : ( n33652 ) ;
assign n33654 =  ( n32871 ) ? ( VREG_24_7 ) : ( n33653 ) ;
assign n33655 =  ( n32870 ) ? ( VREG_24_8 ) : ( n33654 ) ;
assign n33656 =  ( n32869 ) ? ( VREG_24_9 ) : ( n33655 ) ;
assign n33657 =  ( n32868 ) ? ( VREG_24_10 ) : ( n33656 ) ;
assign n33658 =  ( n32867 ) ? ( VREG_24_11 ) : ( n33657 ) ;
assign n33659 =  ( n32866 ) ? ( VREG_24_12 ) : ( n33658 ) ;
assign n33660 =  ( n32865 ) ? ( VREG_24_13 ) : ( n33659 ) ;
assign n33661 =  ( n32864 ) ? ( VREG_24_14 ) : ( n33660 ) ;
assign n33662 =  ( n32863 ) ? ( VREG_24_15 ) : ( n33661 ) ;
assign n33663 =  ( n32862 ) ? ( VREG_25_0 ) : ( n33662 ) ;
assign n33664 =  ( n32861 ) ? ( VREG_25_1 ) : ( n33663 ) ;
assign n33665 =  ( n32860 ) ? ( VREG_25_2 ) : ( n33664 ) ;
assign n33666 =  ( n32859 ) ? ( VREG_25_3 ) : ( n33665 ) ;
assign n33667 =  ( n32858 ) ? ( VREG_25_4 ) : ( n33666 ) ;
assign n33668 =  ( n32857 ) ? ( VREG_25_5 ) : ( n33667 ) ;
assign n33669 =  ( n32856 ) ? ( VREG_25_6 ) : ( n33668 ) ;
assign n33670 =  ( n32855 ) ? ( VREG_25_7 ) : ( n33669 ) ;
assign n33671 =  ( n32854 ) ? ( VREG_25_8 ) : ( n33670 ) ;
assign n33672 =  ( n32853 ) ? ( VREG_25_9 ) : ( n33671 ) ;
assign n33673 =  ( n32852 ) ? ( VREG_25_10 ) : ( n33672 ) ;
assign n33674 =  ( n32851 ) ? ( VREG_25_11 ) : ( n33673 ) ;
assign n33675 =  ( n32850 ) ? ( VREG_25_12 ) : ( n33674 ) ;
assign n33676 =  ( n32849 ) ? ( VREG_25_13 ) : ( n33675 ) ;
assign n33677 =  ( n32848 ) ? ( VREG_25_14 ) : ( n33676 ) ;
assign n33678 =  ( n32847 ) ? ( VREG_25_15 ) : ( n33677 ) ;
assign n33679 =  ( n32846 ) ? ( VREG_26_0 ) : ( n33678 ) ;
assign n33680 =  ( n32845 ) ? ( VREG_26_1 ) : ( n33679 ) ;
assign n33681 =  ( n32844 ) ? ( VREG_26_2 ) : ( n33680 ) ;
assign n33682 =  ( n32843 ) ? ( VREG_26_3 ) : ( n33681 ) ;
assign n33683 =  ( n32842 ) ? ( VREG_26_4 ) : ( n33682 ) ;
assign n33684 =  ( n32841 ) ? ( VREG_26_5 ) : ( n33683 ) ;
assign n33685 =  ( n32840 ) ? ( VREG_26_6 ) : ( n33684 ) ;
assign n33686 =  ( n32839 ) ? ( VREG_26_7 ) : ( n33685 ) ;
assign n33687 =  ( n32838 ) ? ( VREG_26_8 ) : ( n33686 ) ;
assign n33688 =  ( n32837 ) ? ( VREG_26_9 ) : ( n33687 ) ;
assign n33689 =  ( n32836 ) ? ( VREG_26_10 ) : ( n33688 ) ;
assign n33690 =  ( n32835 ) ? ( VREG_26_11 ) : ( n33689 ) ;
assign n33691 =  ( n32834 ) ? ( VREG_26_12 ) : ( n33690 ) ;
assign n33692 =  ( n32833 ) ? ( VREG_26_13 ) : ( n33691 ) ;
assign n33693 =  ( n32832 ) ? ( VREG_26_14 ) : ( n33692 ) ;
assign n33694 =  ( n32831 ) ? ( VREG_26_15 ) : ( n33693 ) ;
assign n33695 =  ( n32830 ) ? ( VREG_27_0 ) : ( n33694 ) ;
assign n33696 =  ( n32829 ) ? ( VREG_27_1 ) : ( n33695 ) ;
assign n33697 =  ( n32828 ) ? ( VREG_27_2 ) : ( n33696 ) ;
assign n33698 =  ( n32827 ) ? ( VREG_27_3 ) : ( n33697 ) ;
assign n33699 =  ( n32826 ) ? ( VREG_27_4 ) : ( n33698 ) ;
assign n33700 =  ( n32825 ) ? ( VREG_27_5 ) : ( n33699 ) ;
assign n33701 =  ( n32824 ) ? ( VREG_27_6 ) : ( n33700 ) ;
assign n33702 =  ( n32823 ) ? ( VREG_27_7 ) : ( n33701 ) ;
assign n33703 =  ( n32822 ) ? ( VREG_27_8 ) : ( n33702 ) ;
assign n33704 =  ( n32821 ) ? ( VREG_27_9 ) : ( n33703 ) ;
assign n33705 =  ( n32820 ) ? ( VREG_27_10 ) : ( n33704 ) ;
assign n33706 =  ( n32819 ) ? ( VREG_27_11 ) : ( n33705 ) ;
assign n33707 =  ( n32818 ) ? ( VREG_27_12 ) : ( n33706 ) ;
assign n33708 =  ( n32817 ) ? ( VREG_27_13 ) : ( n33707 ) ;
assign n33709 =  ( n32816 ) ? ( VREG_27_14 ) : ( n33708 ) ;
assign n33710 =  ( n32815 ) ? ( VREG_27_15 ) : ( n33709 ) ;
assign n33711 =  ( n32814 ) ? ( VREG_28_0 ) : ( n33710 ) ;
assign n33712 =  ( n32813 ) ? ( VREG_28_1 ) : ( n33711 ) ;
assign n33713 =  ( n32812 ) ? ( VREG_28_2 ) : ( n33712 ) ;
assign n33714 =  ( n32811 ) ? ( VREG_28_3 ) : ( n33713 ) ;
assign n33715 =  ( n32810 ) ? ( VREG_28_4 ) : ( n33714 ) ;
assign n33716 =  ( n32809 ) ? ( VREG_28_5 ) : ( n33715 ) ;
assign n33717 =  ( n32808 ) ? ( VREG_28_6 ) : ( n33716 ) ;
assign n33718 =  ( n32807 ) ? ( VREG_28_7 ) : ( n33717 ) ;
assign n33719 =  ( n32806 ) ? ( VREG_28_8 ) : ( n33718 ) ;
assign n33720 =  ( n32805 ) ? ( VREG_28_9 ) : ( n33719 ) ;
assign n33721 =  ( n32804 ) ? ( VREG_28_10 ) : ( n33720 ) ;
assign n33722 =  ( n32803 ) ? ( VREG_28_11 ) : ( n33721 ) ;
assign n33723 =  ( n32802 ) ? ( VREG_28_12 ) : ( n33722 ) ;
assign n33724 =  ( n32801 ) ? ( VREG_28_13 ) : ( n33723 ) ;
assign n33725 =  ( n32800 ) ? ( VREG_28_14 ) : ( n33724 ) ;
assign n33726 =  ( n32799 ) ? ( VREG_28_15 ) : ( n33725 ) ;
assign n33727 =  ( n32798 ) ? ( VREG_29_0 ) : ( n33726 ) ;
assign n33728 =  ( n32797 ) ? ( VREG_29_1 ) : ( n33727 ) ;
assign n33729 =  ( n32796 ) ? ( VREG_29_2 ) : ( n33728 ) ;
assign n33730 =  ( n32795 ) ? ( VREG_29_3 ) : ( n33729 ) ;
assign n33731 =  ( n32794 ) ? ( VREG_29_4 ) : ( n33730 ) ;
assign n33732 =  ( n32793 ) ? ( VREG_29_5 ) : ( n33731 ) ;
assign n33733 =  ( n32792 ) ? ( VREG_29_6 ) : ( n33732 ) ;
assign n33734 =  ( n32791 ) ? ( VREG_29_7 ) : ( n33733 ) ;
assign n33735 =  ( n32790 ) ? ( VREG_29_8 ) : ( n33734 ) ;
assign n33736 =  ( n32789 ) ? ( VREG_29_9 ) : ( n33735 ) ;
assign n33737 =  ( n32788 ) ? ( VREG_29_10 ) : ( n33736 ) ;
assign n33738 =  ( n32787 ) ? ( VREG_29_11 ) : ( n33737 ) ;
assign n33739 =  ( n32786 ) ? ( VREG_29_12 ) : ( n33738 ) ;
assign n33740 =  ( n32785 ) ? ( VREG_29_13 ) : ( n33739 ) ;
assign n33741 =  ( n32784 ) ? ( VREG_29_14 ) : ( n33740 ) ;
assign n33742 =  ( n32783 ) ? ( VREG_29_15 ) : ( n33741 ) ;
assign n33743 =  ( n32782 ) ? ( VREG_30_0 ) : ( n33742 ) ;
assign n33744 =  ( n32781 ) ? ( VREG_30_1 ) : ( n33743 ) ;
assign n33745 =  ( n32780 ) ? ( VREG_30_2 ) : ( n33744 ) ;
assign n33746 =  ( n32779 ) ? ( VREG_30_3 ) : ( n33745 ) ;
assign n33747 =  ( n32778 ) ? ( VREG_30_4 ) : ( n33746 ) ;
assign n33748 =  ( n32777 ) ? ( VREG_30_5 ) : ( n33747 ) ;
assign n33749 =  ( n32776 ) ? ( VREG_30_6 ) : ( n33748 ) ;
assign n33750 =  ( n32775 ) ? ( VREG_30_7 ) : ( n33749 ) ;
assign n33751 =  ( n32774 ) ? ( VREG_30_8 ) : ( n33750 ) ;
assign n33752 =  ( n32773 ) ? ( VREG_30_9 ) : ( n33751 ) ;
assign n33753 =  ( n32772 ) ? ( VREG_30_10 ) : ( n33752 ) ;
assign n33754 =  ( n32771 ) ? ( VREG_30_11 ) : ( n33753 ) ;
assign n33755 =  ( n32770 ) ? ( VREG_30_12 ) : ( n33754 ) ;
assign n33756 =  ( n32769 ) ? ( VREG_30_13 ) : ( n33755 ) ;
assign n33757 =  ( n32768 ) ? ( VREG_30_14 ) : ( n33756 ) ;
assign n33758 =  ( n32767 ) ? ( VREG_30_15 ) : ( n33757 ) ;
assign n33759 =  ( n32766 ) ? ( VREG_31_0 ) : ( n33758 ) ;
assign n33760 =  ( n32764 ) ? ( VREG_31_1 ) : ( n33759 ) ;
assign n33761 =  ( n32762 ) ? ( VREG_31_2 ) : ( n33760 ) ;
assign n33762 =  ( n32760 ) ? ( VREG_31_3 ) : ( n33761 ) ;
assign n33763 =  ( n32758 ) ? ( VREG_31_4 ) : ( n33762 ) ;
assign n33764 =  ( n32756 ) ? ( VREG_31_5 ) : ( n33763 ) ;
assign n33765 =  ( n32754 ) ? ( VREG_31_6 ) : ( n33764 ) ;
assign n33766 =  ( n32752 ) ? ( VREG_31_7 ) : ( n33765 ) ;
assign n33767 =  ( n32750 ) ? ( VREG_31_8 ) : ( n33766 ) ;
assign n33768 =  ( n32748 ) ? ( VREG_31_9 ) : ( n33767 ) ;
assign n33769 =  ( n32746 ) ? ( VREG_31_10 ) : ( n33768 ) ;
assign n33770 =  ( n32744 ) ? ( VREG_31_11 ) : ( n33769 ) ;
assign n33771 =  ( n32742 ) ? ( VREG_31_12 ) : ( n33770 ) ;
assign n33772 =  ( n32740 ) ? ( VREG_31_13 ) : ( n33771 ) ;
assign n33773 =  ( n32738 ) ? ( VREG_31_14 ) : ( n33772 ) ;
assign n33774 =  ( n32736 ) ? ( VREG_31_15 ) : ( n33773 ) ;
assign n33775 =  ( n33774 ) + ( n140 )  ;
assign n33776 =  ( n33774 ) - ( n140 )  ;
assign n33777 =  ( n33774 ) & ( n140 )  ;
assign n33778 =  ( n33774 ) | ( n140 )  ;
assign n33779 =  ( ( n33774 ) * ( n140 ))  ;
assign n33780 =  ( n148 ) ? ( n33779 ) : ( VREG_0_9 ) ;
assign n33781 =  ( n146 ) ? ( n33778 ) : ( n33780 ) ;
assign n33782 =  ( n144 ) ? ( n33777 ) : ( n33781 ) ;
assign n33783 =  ( n142 ) ? ( n33776 ) : ( n33782 ) ;
assign n33784 =  ( n10 ) ? ( n33775 ) : ( n33783 ) ;
assign n33785 =  ( n77 ) & ( n32735 )  ;
assign n33786 =  ( n77 ) & ( n32737 )  ;
assign n33787 =  ( n77 ) & ( n32739 )  ;
assign n33788 =  ( n77 ) & ( n32741 )  ;
assign n33789 =  ( n77 ) & ( n32743 )  ;
assign n33790 =  ( n77 ) & ( n32745 )  ;
assign n33791 =  ( n77 ) & ( n32747 )  ;
assign n33792 =  ( n77 ) & ( n32749 )  ;
assign n33793 =  ( n77 ) & ( n32751 )  ;
assign n33794 =  ( n77 ) & ( n32753 )  ;
assign n33795 =  ( n77 ) & ( n32755 )  ;
assign n33796 =  ( n77 ) & ( n32757 )  ;
assign n33797 =  ( n77 ) & ( n32759 )  ;
assign n33798 =  ( n77 ) & ( n32761 )  ;
assign n33799 =  ( n77 ) & ( n32763 )  ;
assign n33800 =  ( n77 ) & ( n32765 )  ;
assign n33801 =  ( n78 ) & ( n32735 )  ;
assign n33802 =  ( n78 ) & ( n32737 )  ;
assign n33803 =  ( n78 ) & ( n32739 )  ;
assign n33804 =  ( n78 ) & ( n32741 )  ;
assign n33805 =  ( n78 ) & ( n32743 )  ;
assign n33806 =  ( n78 ) & ( n32745 )  ;
assign n33807 =  ( n78 ) & ( n32747 )  ;
assign n33808 =  ( n78 ) & ( n32749 )  ;
assign n33809 =  ( n78 ) & ( n32751 )  ;
assign n33810 =  ( n78 ) & ( n32753 )  ;
assign n33811 =  ( n78 ) & ( n32755 )  ;
assign n33812 =  ( n78 ) & ( n32757 )  ;
assign n33813 =  ( n78 ) & ( n32759 )  ;
assign n33814 =  ( n78 ) & ( n32761 )  ;
assign n33815 =  ( n78 ) & ( n32763 )  ;
assign n33816 =  ( n78 ) & ( n32765 )  ;
assign n33817 =  ( n79 ) & ( n32735 )  ;
assign n33818 =  ( n79 ) & ( n32737 )  ;
assign n33819 =  ( n79 ) & ( n32739 )  ;
assign n33820 =  ( n79 ) & ( n32741 )  ;
assign n33821 =  ( n79 ) & ( n32743 )  ;
assign n33822 =  ( n79 ) & ( n32745 )  ;
assign n33823 =  ( n79 ) & ( n32747 )  ;
assign n33824 =  ( n79 ) & ( n32749 )  ;
assign n33825 =  ( n79 ) & ( n32751 )  ;
assign n33826 =  ( n79 ) & ( n32753 )  ;
assign n33827 =  ( n79 ) & ( n32755 )  ;
assign n33828 =  ( n79 ) & ( n32757 )  ;
assign n33829 =  ( n79 ) & ( n32759 )  ;
assign n33830 =  ( n79 ) & ( n32761 )  ;
assign n33831 =  ( n79 ) & ( n32763 )  ;
assign n33832 =  ( n79 ) & ( n32765 )  ;
assign n33833 =  ( n80 ) & ( n32735 )  ;
assign n33834 =  ( n80 ) & ( n32737 )  ;
assign n33835 =  ( n80 ) & ( n32739 )  ;
assign n33836 =  ( n80 ) & ( n32741 )  ;
assign n33837 =  ( n80 ) & ( n32743 )  ;
assign n33838 =  ( n80 ) & ( n32745 )  ;
assign n33839 =  ( n80 ) & ( n32747 )  ;
assign n33840 =  ( n80 ) & ( n32749 )  ;
assign n33841 =  ( n80 ) & ( n32751 )  ;
assign n33842 =  ( n80 ) & ( n32753 )  ;
assign n33843 =  ( n80 ) & ( n32755 )  ;
assign n33844 =  ( n80 ) & ( n32757 )  ;
assign n33845 =  ( n80 ) & ( n32759 )  ;
assign n33846 =  ( n80 ) & ( n32761 )  ;
assign n33847 =  ( n80 ) & ( n32763 )  ;
assign n33848 =  ( n80 ) & ( n32765 )  ;
assign n33849 =  ( n81 ) & ( n32735 )  ;
assign n33850 =  ( n81 ) & ( n32737 )  ;
assign n33851 =  ( n81 ) & ( n32739 )  ;
assign n33852 =  ( n81 ) & ( n32741 )  ;
assign n33853 =  ( n81 ) & ( n32743 )  ;
assign n33854 =  ( n81 ) & ( n32745 )  ;
assign n33855 =  ( n81 ) & ( n32747 )  ;
assign n33856 =  ( n81 ) & ( n32749 )  ;
assign n33857 =  ( n81 ) & ( n32751 )  ;
assign n33858 =  ( n81 ) & ( n32753 )  ;
assign n33859 =  ( n81 ) & ( n32755 )  ;
assign n33860 =  ( n81 ) & ( n32757 )  ;
assign n33861 =  ( n81 ) & ( n32759 )  ;
assign n33862 =  ( n81 ) & ( n32761 )  ;
assign n33863 =  ( n81 ) & ( n32763 )  ;
assign n33864 =  ( n81 ) & ( n32765 )  ;
assign n33865 =  ( n82 ) & ( n32735 )  ;
assign n33866 =  ( n82 ) & ( n32737 )  ;
assign n33867 =  ( n82 ) & ( n32739 )  ;
assign n33868 =  ( n82 ) & ( n32741 )  ;
assign n33869 =  ( n82 ) & ( n32743 )  ;
assign n33870 =  ( n82 ) & ( n32745 )  ;
assign n33871 =  ( n82 ) & ( n32747 )  ;
assign n33872 =  ( n82 ) & ( n32749 )  ;
assign n33873 =  ( n82 ) & ( n32751 )  ;
assign n33874 =  ( n82 ) & ( n32753 )  ;
assign n33875 =  ( n82 ) & ( n32755 )  ;
assign n33876 =  ( n82 ) & ( n32757 )  ;
assign n33877 =  ( n82 ) & ( n32759 )  ;
assign n33878 =  ( n82 ) & ( n32761 )  ;
assign n33879 =  ( n82 ) & ( n32763 )  ;
assign n33880 =  ( n82 ) & ( n32765 )  ;
assign n33881 =  ( n83 ) & ( n32735 )  ;
assign n33882 =  ( n83 ) & ( n32737 )  ;
assign n33883 =  ( n83 ) & ( n32739 )  ;
assign n33884 =  ( n83 ) & ( n32741 )  ;
assign n33885 =  ( n83 ) & ( n32743 )  ;
assign n33886 =  ( n83 ) & ( n32745 )  ;
assign n33887 =  ( n83 ) & ( n32747 )  ;
assign n33888 =  ( n83 ) & ( n32749 )  ;
assign n33889 =  ( n83 ) & ( n32751 )  ;
assign n33890 =  ( n83 ) & ( n32753 )  ;
assign n33891 =  ( n83 ) & ( n32755 )  ;
assign n33892 =  ( n83 ) & ( n32757 )  ;
assign n33893 =  ( n83 ) & ( n32759 )  ;
assign n33894 =  ( n83 ) & ( n32761 )  ;
assign n33895 =  ( n83 ) & ( n32763 )  ;
assign n33896 =  ( n83 ) & ( n32765 )  ;
assign n33897 =  ( n84 ) & ( n32735 )  ;
assign n33898 =  ( n84 ) & ( n32737 )  ;
assign n33899 =  ( n84 ) & ( n32739 )  ;
assign n33900 =  ( n84 ) & ( n32741 )  ;
assign n33901 =  ( n84 ) & ( n32743 )  ;
assign n33902 =  ( n84 ) & ( n32745 )  ;
assign n33903 =  ( n84 ) & ( n32747 )  ;
assign n33904 =  ( n84 ) & ( n32749 )  ;
assign n33905 =  ( n84 ) & ( n32751 )  ;
assign n33906 =  ( n84 ) & ( n32753 )  ;
assign n33907 =  ( n84 ) & ( n32755 )  ;
assign n33908 =  ( n84 ) & ( n32757 )  ;
assign n33909 =  ( n84 ) & ( n32759 )  ;
assign n33910 =  ( n84 ) & ( n32761 )  ;
assign n33911 =  ( n84 ) & ( n32763 )  ;
assign n33912 =  ( n84 ) & ( n32765 )  ;
assign n33913 =  ( n85 ) & ( n32735 )  ;
assign n33914 =  ( n85 ) & ( n32737 )  ;
assign n33915 =  ( n85 ) & ( n32739 )  ;
assign n33916 =  ( n85 ) & ( n32741 )  ;
assign n33917 =  ( n85 ) & ( n32743 )  ;
assign n33918 =  ( n85 ) & ( n32745 )  ;
assign n33919 =  ( n85 ) & ( n32747 )  ;
assign n33920 =  ( n85 ) & ( n32749 )  ;
assign n33921 =  ( n85 ) & ( n32751 )  ;
assign n33922 =  ( n85 ) & ( n32753 )  ;
assign n33923 =  ( n85 ) & ( n32755 )  ;
assign n33924 =  ( n85 ) & ( n32757 )  ;
assign n33925 =  ( n85 ) & ( n32759 )  ;
assign n33926 =  ( n85 ) & ( n32761 )  ;
assign n33927 =  ( n85 ) & ( n32763 )  ;
assign n33928 =  ( n85 ) & ( n32765 )  ;
assign n33929 =  ( n86 ) & ( n32735 )  ;
assign n33930 =  ( n86 ) & ( n32737 )  ;
assign n33931 =  ( n86 ) & ( n32739 )  ;
assign n33932 =  ( n86 ) & ( n32741 )  ;
assign n33933 =  ( n86 ) & ( n32743 )  ;
assign n33934 =  ( n86 ) & ( n32745 )  ;
assign n33935 =  ( n86 ) & ( n32747 )  ;
assign n33936 =  ( n86 ) & ( n32749 )  ;
assign n33937 =  ( n86 ) & ( n32751 )  ;
assign n33938 =  ( n86 ) & ( n32753 )  ;
assign n33939 =  ( n86 ) & ( n32755 )  ;
assign n33940 =  ( n86 ) & ( n32757 )  ;
assign n33941 =  ( n86 ) & ( n32759 )  ;
assign n33942 =  ( n86 ) & ( n32761 )  ;
assign n33943 =  ( n86 ) & ( n32763 )  ;
assign n33944 =  ( n86 ) & ( n32765 )  ;
assign n33945 =  ( n87 ) & ( n32735 )  ;
assign n33946 =  ( n87 ) & ( n32737 )  ;
assign n33947 =  ( n87 ) & ( n32739 )  ;
assign n33948 =  ( n87 ) & ( n32741 )  ;
assign n33949 =  ( n87 ) & ( n32743 )  ;
assign n33950 =  ( n87 ) & ( n32745 )  ;
assign n33951 =  ( n87 ) & ( n32747 )  ;
assign n33952 =  ( n87 ) & ( n32749 )  ;
assign n33953 =  ( n87 ) & ( n32751 )  ;
assign n33954 =  ( n87 ) & ( n32753 )  ;
assign n33955 =  ( n87 ) & ( n32755 )  ;
assign n33956 =  ( n87 ) & ( n32757 )  ;
assign n33957 =  ( n87 ) & ( n32759 )  ;
assign n33958 =  ( n87 ) & ( n32761 )  ;
assign n33959 =  ( n87 ) & ( n32763 )  ;
assign n33960 =  ( n87 ) & ( n32765 )  ;
assign n33961 =  ( n88 ) & ( n32735 )  ;
assign n33962 =  ( n88 ) & ( n32737 )  ;
assign n33963 =  ( n88 ) & ( n32739 )  ;
assign n33964 =  ( n88 ) & ( n32741 )  ;
assign n33965 =  ( n88 ) & ( n32743 )  ;
assign n33966 =  ( n88 ) & ( n32745 )  ;
assign n33967 =  ( n88 ) & ( n32747 )  ;
assign n33968 =  ( n88 ) & ( n32749 )  ;
assign n33969 =  ( n88 ) & ( n32751 )  ;
assign n33970 =  ( n88 ) & ( n32753 )  ;
assign n33971 =  ( n88 ) & ( n32755 )  ;
assign n33972 =  ( n88 ) & ( n32757 )  ;
assign n33973 =  ( n88 ) & ( n32759 )  ;
assign n33974 =  ( n88 ) & ( n32761 )  ;
assign n33975 =  ( n88 ) & ( n32763 )  ;
assign n33976 =  ( n88 ) & ( n32765 )  ;
assign n33977 =  ( n89 ) & ( n32735 )  ;
assign n33978 =  ( n89 ) & ( n32737 )  ;
assign n33979 =  ( n89 ) & ( n32739 )  ;
assign n33980 =  ( n89 ) & ( n32741 )  ;
assign n33981 =  ( n89 ) & ( n32743 )  ;
assign n33982 =  ( n89 ) & ( n32745 )  ;
assign n33983 =  ( n89 ) & ( n32747 )  ;
assign n33984 =  ( n89 ) & ( n32749 )  ;
assign n33985 =  ( n89 ) & ( n32751 )  ;
assign n33986 =  ( n89 ) & ( n32753 )  ;
assign n33987 =  ( n89 ) & ( n32755 )  ;
assign n33988 =  ( n89 ) & ( n32757 )  ;
assign n33989 =  ( n89 ) & ( n32759 )  ;
assign n33990 =  ( n89 ) & ( n32761 )  ;
assign n33991 =  ( n89 ) & ( n32763 )  ;
assign n33992 =  ( n89 ) & ( n32765 )  ;
assign n33993 =  ( n90 ) & ( n32735 )  ;
assign n33994 =  ( n90 ) & ( n32737 )  ;
assign n33995 =  ( n90 ) & ( n32739 )  ;
assign n33996 =  ( n90 ) & ( n32741 )  ;
assign n33997 =  ( n90 ) & ( n32743 )  ;
assign n33998 =  ( n90 ) & ( n32745 )  ;
assign n33999 =  ( n90 ) & ( n32747 )  ;
assign n34000 =  ( n90 ) & ( n32749 )  ;
assign n34001 =  ( n90 ) & ( n32751 )  ;
assign n34002 =  ( n90 ) & ( n32753 )  ;
assign n34003 =  ( n90 ) & ( n32755 )  ;
assign n34004 =  ( n90 ) & ( n32757 )  ;
assign n34005 =  ( n90 ) & ( n32759 )  ;
assign n34006 =  ( n90 ) & ( n32761 )  ;
assign n34007 =  ( n90 ) & ( n32763 )  ;
assign n34008 =  ( n90 ) & ( n32765 )  ;
assign n34009 =  ( n91 ) & ( n32735 )  ;
assign n34010 =  ( n91 ) & ( n32737 )  ;
assign n34011 =  ( n91 ) & ( n32739 )  ;
assign n34012 =  ( n91 ) & ( n32741 )  ;
assign n34013 =  ( n91 ) & ( n32743 )  ;
assign n34014 =  ( n91 ) & ( n32745 )  ;
assign n34015 =  ( n91 ) & ( n32747 )  ;
assign n34016 =  ( n91 ) & ( n32749 )  ;
assign n34017 =  ( n91 ) & ( n32751 )  ;
assign n34018 =  ( n91 ) & ( n32753 )  ;
assign n34019 =  ( n91 ) & ( n32755 )  ;
assign n34020 =  ( n91 ) & ( n32757 )  ;
assign n34021 =  ( n91 ) & ( n32759 )  ;
assign n34022 =  ( n91 ) & ( n32761 )  ;
assign n34023 =  ( n91 ) & ( n32763 )  ;
assign n34024 =  ( n91 ) & ( n32765 )  ;
assign n34025 =  ( n92 ) & ( n32735 )  ;
assign n34026 =  ( n92 ) & ( n32737 )  ;
assign n34027 =  ( n92 ) & ( n32739 )  ;
assign n34028 =  ( n92 ) & ( n32741 )  ;
assign n34029 =  ( n92 ) & ( n32743 )  ;
assign n34030 =  ( n92 ) & ( n32745 )  ;
assign n34031 =  ( n92 ) & ( n32747 )  ;
assign n34032 =  ( n92 ) & ( n32749 )  ;
assign n34033 =  ( n92 ) & ( n32751 )  ;
assign n34034 =  ( n92 ) & ( n32753 )  ;
assign n34035 =  ( n92 ) & ( n32755 )  ;
assign n34036 =  ( n92 ) & ( n32757 )  ;
assign n34037 =  ( n92 ) & ( n32759 )  ;
assign n34038 =  ( n92 ) & ( n32761 )  ;
assign n34039 =  ( n92 ) & ( n32763 )  ;
assign n34040 =  ( n92 ) & ( n32765 )  ;
assign n34041 =  ( n93 ) & ( n32735 )  ;
assign n34042 =  ( n93 ) & ( n32737 )  ;
assign n34043 =  ( n93 ) & ( n32739 )  ;
assign n34044 =  ( n93 ) & ( n32741 )  ;
assign n34045 =  ( n93 ) & ( n32743 )  ;
assign n34046 =  ( n93 ) & ( n32745 )  ;
assign n34047 =  ( n93 ) & ( n32747 )  ;
assign n34048 =  ( n93 ) & ( n32749 )  ;
assign n34049 =  ( n93 ) & ( n32751 )  ;
assign n34050 =  ( n93 ) & ( n32753 )  ;
assign n34051 =  ( n93 ) & ( n32755 )  ;
assign n34052 =  ( n93 ) & ( n32757 )  ;
assign n34053 =  ( n93 ) & ( n32759 )  ;
assign n34054 =  ( n93 ) & ( n32761 )  ;
assign n34055 =  ( n93 ) & ( n32763 )  ;
assign n34056 =  ( n93 ) & ( n32765 )  ;
assign n34057 =  ( n94 ) & ( n32735 )  ;
assign n34058 =  ( n94 ) & ( n32737 )  ;
assign n34059 =  ( n94 ) & ( n32739 )  ;
assign n34060 =  ( n94 ) & ( n32741 )  ;
assign n34061 =  ( n94 ) & ( n32743 )  ;
assign n34062 =  ( n94 ) & ( n32745 )  ;
assign n34063 =  ( n94 ) & ( n32747 )  ;
assign n34064 =  ( n94 ) & ( n32749 )  ;
assign n34065 =  ( n94 ) & ( n32751 )  ;
assign n34066 =  ( n94 ) & ( n32753 )  ;
assign n34067 =  ( n94 ) & ( n32755 )  ;
assign n34068 =  ( n94 ) & ( n32757 )  ;
assign n34069 =  ( n94 ) & ( n32759 )  ;
assign n34070 =  ( n94 ) & ( n32761 )  ;
assign n34071 =  ( n94 ) & ( n32763 )  ;
assign n34072 =  ( n94 ) & ( n32765 )  ;
assign n34073 =  ( n95 ) & ( n32735 )  ;
assign n34074 =  ( n95 ) & ( n32737 )  ;
assign n34075 =  ( n95 ) & ( n32739 )  ;
assign n34076 =  ( n95 ) & ( n32741 )  ;
assign n34077 =  ( n95 ) & ( n32743 )  ;
assign n34078 =  ( n95 ) & ( n32745 )  ;
assign n34079 =  ( n95 ) & ( n32747 )  ;
assign n34080 =  ( n95 ) & ( n32749 )  ;
assign n34081 =  ( n95 ) & ( n32751 )  ;
assign n34082 =  ( n95 ) & ( n32753 )  ;
assign n34083 =  ( n95 ) & ( n32755 )  ;
assign n34084 =  ( n95 ) & ( n32757 )  ;
assign n34085 =  ( n95 ) & ( n32759 )  ;
assign n34086 =  ( n95 ) & ( n32761 )  ;
assign n34087 =  ( n95 ) & ( n32763 )  ;
assign n34088 =  ( n95 ) & ( n32765 )  ;
assign n34089 =  ( n96 ) & ( n32735 )  ;
assign n34090 =  ( n96 ) & ( n32737 )  ;
assign n34091 =  ( n96 ) & ( n32739 )  ;
assign n34092 =  ( n96 ) & ( n32741 )  ;
assign n34093 =  ( n96 ) & ( n32743 )  ;
assign n34094 =  ( n96 ) & ( n32745 )  ;
assign n34095 =  ( n96 ) & ( n32747 )  ;
assign n34096 =  ( n96 ) & ( n32749 )  ;
assign n34097 =  ( n96 ) & ( n32751 )  ;
assign n34098 =  ( n96 ) & ( n32753 )  ;
assign n34099 =  ( n96 ) & ( n32755 )  ;
assign n34100 =  ( n96 ) & ( n32757 )  ;
assign n34101 =  ( n96 ) & ( n32759 )  ;
assign n34102 =  ( n96 ) & ( n32761 )  ;
assign n34103 =  ( n96 ) & ( n32763 )  ;
assign n34104 =  ( n96 ) & ( n32765 )  ;
assign n34105 =  ( n97 ) & ( n32735 )  ;
assign n34106 =  ( n97 ) & ( n32737 )  ;
assign n34107 =  ( n97 ) & ( n32739 )  ;
assign n34108 =  ( n97 ) & ( n32741 )  ;
assign n34109 =  ( n97 ) & ( n32743 )  ;
assign n34110 =  ( n97 ) & ( n32745 )  ;
assign n34111 =  ( n97 ) & ( n32747 )  ;
assign n34112 =  ( n97 ) & ( n32749 )  ;
assign n34113 =  ( n97 ) & ( n32751 )  ;
assign n34114 =  ( n97 ) & ( n32753 )  ;
assign n34115 =  ( n97 ) & ( n32755 )  ;
assign n34116 =  ( n97 ) & ( n32757 )  ;
assign n34117 =  ( n97 ) & ( n32759 )  ;
assign n34118 =  ( n97 ) & ( n32761 )  ;
assign n34119 =  ( n97 ) & ( n32763 )  ;
assign n34120 =  ( n97 ) & ( n32765 )  ;
assign n34121 =  ( n98 ) & ( n32735 )  ;
assign n34122 =  ( n98 ) & ( n32737 )  ;
assign n34123 =  ( n98 ) & ( n32739 )  ;
assign n34124 =  ( n98 ) & ( n32741 )  ;
assign n34125 =  ( n98 ) & ( n32743 )  ;
assign n34126 =  ( n98 ) & ( n32745 )  ;
assign n34127 =  ( n98 ) & ( n32747 )  ;
assign n34128 =  ( n98 ) & ( n32749 )  ;
assign n34129 =  ( n98 ) & ( n32751 )  ;
assign n34130 =  ( n98 ) & ( n32753 )  ;
assign n34131 =  ( n98 ) & ( n32755 )  ;
assign n34132 =  ( n98 ) & ( n32757 )  ;
assign n34133 =  ( n98 ) & ( n32759 )  ;
assign n34134 =  ( n98 ) & ( n32761 )  ;
assign n34135 =  ( n98 ) & ( n32763 )  ;
assign n34136 =  ( n98 ) & ( n32765 )  ;
assign n34137 =  ( n99 ) & ( n32735 )  ;
assign n34138 =  ( n99 ) & ( n32737 )  ;
assign n34139 =  ( n99 ) & ( n32739 )  ;
assign n34140 =  ( n99 ) & ( n32741 )  ;
assign n34141 =  ( n99 ) & ( n32743 )  ;
assign n34142 =  ( n99 ) & ( n32745 )  ;
assign n34143 =  ( n99 ) & ( n32747 )  ;
assign n34144 =  ( n99 ) & ( n32749 )  ;
assign n34145 =  ( n99 ) & ( n32751 )  ;
assign n34146 =  ( n99 ) & ( n32753 )  ;
assign n34147 =  ( n99 ) & ( n32755 )  ;
assign n34148 =  ( n99 ) & ( n32757 )  ;
assign n34149 =  ( n99 ) & ( n32759 )  ;
assign n34150 =  ( n99 ) & ( n32761 )  ;
assign n34151 =  ( n99 ) & ( n32763 )  ;
assign n34152 =  ( n99 ) & ( n32765 )  ;
assign n34153 =  ( n100 ) & ( n32735 )  ;
assign n34154 =  ( n100 ) & ( n32737 )  ;
assign n34155 =  ( n100 ) & ( n32739 )  ;
assign n34156 =  ( n100 ) & ( n32741 )  ;
assign n34157 =  ( n100 ) & ( n32743 )  ;
assign n34158 =  ( n100 ) & ( n32745 )  ;
assign n34159 =  ( n100 ) & ( n32747 )  ;
assign n34160 =  ( n100 ) & ( n32749 )  ;
assign n34161 =  ( n100 ) & ( n32751 )  ;
assign n34162 =  ( n100 ) & ( n32753 )  ;
assign n34163 =  ( n100 ) & ( n32755 )  ;
assign n34164 =  ( n100 ) & ( n32757 )  ;
assign n34165 =  ( n100 ) & ( n32759 )  ;
assign n34166 =  ( n100 ) & ( n32761 )  ;
assign n34167 =  ( n100 ) & ( n32763 )  ;
assign n34168 =  ( n100 ) & ( n32765 )  ;
assign n34169 =  ( n101 ) & ( n32735 )  ;
assign n34170 =  ( n101 ) & ( n32737 )  ;
assign n34171 =  ( n101 ) & ( n32739 )  ;
assign n34172 =  ( n101 ) & ( n32741 )  ;
assign n34173 =  ( n101 ) & ( n32743 )  ;
assign n34174 =  ( n101 ) & ( n32745 )  ;
assign n34175 =  ( n101 ) & ( n32747 )  ;
assign n34176 =  ( n101 ) & ( n32749 )  ;
assign n34177 =  ( n101 ) & ( n32751 )  ;
assign n34178 =  ( n101 ) & ( n32753 )  ;
assign n34179 =  ( n101 ) & ( n32755 )  ;
assign n34180 =  ( n101 ) & ( n32757 )  ;
assign n34181 =  ( n101 ) & ( n32759 )  ;
assign n34182 =  ( n101 ) & ( n32761 )  ;
assign n34183 =  ( n101 ) & ( n32763 )  ;
assign n34184 =  ( n101 ) & ( n32765 )  ;
assign n34185 =  ( n102 ) & ( n32735 )  ;
assign n34186 =  ( n102 ) & ( n32737 )  ;
assign n34187 =  ( n102 ) & ( n32739 )  ;
assign n34188 =  ( n102 ) & ( n32741 )  ;
assign n34189 =  ( n102 ) & ( n32743 )  ;
assign n34190 =  ( n102 ) & ( n32745 )  ;
assign n34191 =  ( n102 ) & ( n32747 )  ;
assign n34192 =  ( n102 ) & ( n32749 )  ;
assign n34193 =  ( n102 ) & ( n32751 )  ;
assign n34194 =  ( n102 ) & ( n32753 )  ;
assign n34195 =  ( n102 ) & ( n32755 )  ;
assign n34196 =  ( n102 ) & ( n32757 )  ;
assign n34197 =  ( n102 ) & ( n32759 )  ;
assign n34198 =  ( n102 ) & ( n32761 )  ;
assign n34199 =  ( n102 ) & ( n32763 )  ;
assign n34200 =  ( n102 ) & ( n32765 )  ;
assign n34201 =  ( n103 ) & ( n32735 )  ;
assign n34202 =  ( n103 ) & ( n32737 )  ;
assign n34203 =  ( n103 ) & ( n32739 )  ;
assign n34204 =  ( n103 ) & ( n32741 )  ;
assign n34205 =  ( n103 ) & ( n32743 )  ;
assign n34206 =  ( n103 ) & ( n32745 )  ;
assign n34207 =  ( n103 ) & ( n32747 )  ;
assign n34208 =  ( n103 ) & ( n32749 )  ;
assign n34209 =  ( n103 ) & ( n32751 )  ;
assign n34210 =  ( n103 ) & ( n32753 )  ;
assign n34211 =  ( n103 ) & ( n32755 )  ;
assign n34212 =  ( n103 ) & ( n32757 )  ;
assign n34213 =  ( n103 ) & ( n32759 )  ;
assign n34214 =  ( n103 ) & ( n32761 )  ;
assign n34215 =  ( n103 ) & ( n32763 )  ;
assign n34216 =  ( n103 ) & ( n32765 )  ;
assign n34217 =  ( n104 ) & ( n32735 )  ;
assign n34218 =  ( n104 ) & ( n32737 )  ;
assign n34219 =  ( n104 ) & ( n32739 )  ;
assign n34220 =  ( n104 ) & ( n32741 )  ;
assign n34221 =  ( n104 ) & ( n32743 )  ;
assign n34222 =  ( n104 ) & ( n32745 )  ;
assign n34223 =  ( n104 ) & ( n32747 )  ;
assign n34224 =  ( n104 ) & ( n32749 )  ;
assign n34225 =  ( n104 ) & ( n32751 )  ;
assign n34226 =  ( n104 ) & ( n32753 )  ;
assign n34227 =  ( n104 ) & ( n32755 )  ;
assign n34228 =  ( n104 ) & ( n32757 )  ;
assign n34229 =  ( n104 ) & ( n32759 )  ;
assign n34230 =  ( n104 ) & ( n32761 )  ;
assign n34231 =  ( n104 ) & ( n32763 )  ;
assign n34232 =  ( n104 ) & ( n32765 )  ;
assign n34233 =  ( n105 ) & ( n32735 )  ;
assign n34234 =  ( n105 ) & ( n32737 )  ;
assign n34235 =  ( n105 ) & ( n32739 )  ;
assign n34236 =  ( n105 ) & ( n32741 )  ;
assign n34237 =  ( n105 ) & ( n32743 )  ;
assign n34238 =  ( n105 ) & ( n32745 )  ;
assign n34239 =  ( n105 ) & ( n32747 )  ;
assign n34240 =  ( n105 ) & ( n32749 )  ;
assign n34241 =  ( n105 ) & ( n32751 )  ;
assign n34242 =  ( n105 ) & ( n32753 )  ;
assign n34243 =  ( n105 ) & ( n32755 )  ;
assign n34244 =  ( n105 ) & ( n32757 )  ;
assign n34245 =  ( n105 ) & ( n32759 )  ;
assign n34246 =  ( n105 ) & ( n32761 )  ;
assign n34247 =  ( n105 ) & ( n32763 )  ;
assign n34248 =  ( n105 ) & ( n32765 )  ;
assign n34249 =  ( n106 ) & ( n32735 )  ;
assign n34250 =  ( n106 ) & ( n32737 )  ;
assign n34251 =  ( n106 ) & ( n32739 )  ;
assign n34252 =  ( n106 ) & ( n32741 )  ;
assign n34253 =  ( n106 ) & ( n32743 )  ;
assign n34254 =  ( n106 ) & ( n32745 )  ;
assign n34255 =  ( n106 ) & ( n32747 )  ;
assign n34256 =  ( n106 ) & ( n32749 )  ;
assign n34257 =  ( n106 ) & ( n32751 )  ;
assign n34258 =  ( n106 ) & ( n32753 )  ;
assign n34259 =  ( n106 ) & ( n32755 )  ;
assign n34260 =  ( n106 ) & ( n32757 )  ;
assign n34261 =  ( n106 ) & ( n32759 )  ;
assign n34262 =  ( n106 ) & ( n32761 )  ;
assign n34263 =  ( n106 ) & ( n32763 )  ;
assign n34264 =  ( n106 ) & ( n32765 )  ;
assign n34265 =  ( n107 ) & ( n32735 )  ;
assign n34266 =  ( n107 ) & ( n32737 )  ;
assign n34267 =  ( n107 ) & ( n32739 )  ;
assign n34268 =  ( n107 ) & ( n32741 )  ;
assign n34269 =  ( n107 ) & ( n32743 )  ;
assign n34270 =  ( n107 ) & ( n32745 )  ;
assign n34271 =  ( n107 ) & ( n32747 )  ;
assign n34272 =  ( n107 ) & ( n32749 )  ;
assign n34273 =  ( n107 ) & ( n32751 )  ;
assign n34274 =  ( n107 ) & ( n32753 )  ;
assign n34275 =  ( n107 ) & ( n32755 )  ;
assign n34276 =  ( n107 ) & ( n32757 )  ;
assign n34277 =  ( n107 ) & ( n32759 )  ;
assign n34278 =  ( n107 ) & ( n32761 )  ;
assign n34279 =  ( n107 ) & ( n32763 )  ;
assign n34280 =  ( n107 ) & ( n32765 )  ;
assign n34281 =  ( n108 ) & ( n32735 )  ;
assign n34282 =  ( n108 ) & ( n32737 )  ;
assign n34283 =  ( n108 ) & ( n32739 )  ;
assign n34284 =  ( n108 ) & ( n32741 )  ;
assign n34285 =  ( n108 ) & ( n32743 )  ;
assign n34286 =  ( n108 ) & ( n32745 )  ;
assign n34287 =  ( n108 ) & ( n32747 )  ;
assign n34288 =  ( n108 ) & ( n32749 )  ;
assign n34289 =  ( n108 ) & ( n32751 )  ;
assign n34290 =  ( n108 ) & ( n32753 )  ;
assign n34291 =  ( n108 ) & ( n32755 )  ;
assign n34292 =  ( n108 ) & ( n32757 )  ;
assign n34293 =  ( n108 ) & ( n32759 )  ;
assign n34294 =  ( n108 ) & ( n32761 )  ;
assign n34295 =  ( n108 ) & ( n32763 )  ;
assign n34296 =  ( n108 ) & ( n32765 )  ;
assign n34297 =  ( n34296 ) ? ( VREG_0_0 ) : ( VREG_0_0 ) ;
assign n34298 =  ( n34295 ) ? ( VREG_0_1 ) : ( n34297 ) ;
assign n34299 =  ( n34294 ) ? ( VREG_0_2 ) : ( n34298 ) ;
assign n34300 =  ( n34293 ) ? ( VREG_0_3 ) : ( n34299 ) ;
assign n34301 =  ( n34292 ) ? ( VREG_0_4 ) : ( n34300 ) ;
assign n34302 =  ( n34291 ) ? ( VREG_0_5 ) : ( n34301 ) ;
assign n34303 =  ( n34290 ) ? ( VREG_0_6 ) : ( n34302 ) ;
assign n34304 =  ( n34289 ) ? ( VREG_0_7 ) : ( n34303 ) ;
assign n34305 =  ( n34288 ) ? ( VREG_0_8 ) : ( n34304 ) ;
assign n34306 =  ( n34287 ) ? ( VREG_0_9 ) : ( n34305 ) ;
assign n34307 =  ( n34286 ) ? ( VREG_0_10 ) : ( n34306 ) ;
assign n34308 =  ( n34285 ) ? ( VREG_0_11 ) : ( n34307 ) ;
assign n34309 =  ( n34284 ) ? ( VREG_0_12 ) : ( n34308 ) ;
assign n34310 =  ( n34283 ) ? ( VREG_0_13 ) : ( n34309 ) ;
assign n34311 =  ( n34282 ) ? ( VREG_0_14 ) : ( n34310 ) ;
assign n34312 =  ( n34281 ) ? ( VREG_0_15 ) : ( n34311 ) ;
assign n34313 =  ( n34280 ) ? ( VREG_1_0 ) : ( n34312 ) ;
assign n34314 =  ( n34279 ) ? ( VREG_1_1 ) : ( n34313 ) ;
assign n34315 =  ( n34278 ) ? ( VREG_1_2 ) : ( n34314 ) ;
assign n34316 =  ( n34277 ) ? ( VREG_1_3 ) : ( n34315 ) ;
assign n34317 =  ( n34276 ) ? ( VREG_1_4 ) : ( n34316 ) ;
assign n34318 =  ( n34275 ) ? ( VREG_1_5 ) : ( n34317 ) ;
assign n34319 =  ( n34274 ) ? ( VREG_1_6 ) : ( n34318 ) ;
assign n34320 =  ( n34273 ) ? ( VREG_1_7 ) : ( n34319 ) ;
assign n34321 =  ( n34272 ) ? ( VREG_1_8 ) : ( n34320 ) ;
assign n34322 =  ( n34271 ) ? ( VREG_1_9 ) : ( n34321 ) ;
assign n34323 =  ( n34270 ) ? ( VREG_1_10 ) : ( n34322 ) ;
assign n34324 =  ( n34269 ) ? ( VREG_1_11 ) : ( n34323 ) ;
assign n34325 =  ( n34268 ) ? ( VREG_1_12 ) : ( n34324 ) ;
assign n34326 =  ( n34267 ) ? ( VREG_1_13 ) : ( n34325 ) ;
assign n34327 =  ( n34266 ) ? ( VREG_1_14 ) : ( n34326 ) ;
assign n34328 =  ( n34265 ) ? ( VREG_1_15 ) : ( n34327 ) ;
assign n34329 =  ( n34264 ) ? ( VREG_2_0 ) : ( n34328 ) ;
assign n34330 =  ( n34263 ) ? ( VREG_2_1 ) : ( n34329 ) ;
assign n34331 =  ( n34262 ) ? ( VREG_2_2 ) : ( n34330 ) ;
assign n34332 =  ( n34261 ) ? ( VREG_2_3 ) : ( n34331 ) ;
assign n34333 =  ( n34260 ) ? ( VREG_2_4 ) : ( n34332 ) ;
assign n34334 =  ( n34259 ) ? ( VREG_2_5 ) : ( n34333 ) ;
assign n34335 =  ( n34258 ) ? ( VREG_2_6 ) : ( n34334 ) ;
assign n34336 =  ( n34257 ) ? ( VREG_2_7 ) : ( n34335 ) ;
assign n34337 =  ( n34256 ) ? ( VREG_2_8 ) : ( n34336 ) ;
assign n34338 =  ( n34255 ) ? ( VREG_2_9 ) : ( n34337 ) ;
assign n34339 =  ( n34254 ) ? ( VREG_2_10 ) : ( n34338 ) ;
assign n34340 =  ( n34253 ) ? ( VREG_2_11 ) : ( n34339 ) ;
assign n34341 =  ( n34252 ) ? ( VREG_2_12 ) : ( n34340 ) ;
assign n34342 =  ( n34251 ) ? ( VREG_2_13 ) : ( n34341 ) ;
assign n34343 =  ( n34250 ) ? ( VREG_2_14 ) : ( n34342 ) ;
assign n34344 =  ( n34249 ) ? ( VREG_2_15 ) : ( n34343 ) ;
assign n34345 =  ( n34248 ) ? ( VREG_3_0 ) : ( n34344 ) ;
assign n34346 =  ( n34247 ) ? ( VREG_3_1 ) : ( n34345 ) ;
assign n34347 =  ( n34246 ) ? ( VREG_3_2 ) : ( n34346 ) ;
assign n34348 =  ( n34245 ) ? ( VREG_3_3 ) : ( n34347 ) ;
assign n34349 =  ( n34244 ) ? ( VREG_3_4 ) : ( n34348 ) ;
assign n34350 =  ( n34243 ) ? ( VREG_3_5 ) : ( n34349 ) ;
assign n34351 =  ( n34242 ) ? ( VREG_3_6 ) : ( n34350 ) ;
assign n34352 =  ( n34241 ) ? ( VREG_3_7 ) : ( n34351 ) ;
assign n34353 =  ( n34240 ) ? ( VREG_3_8 ) : ( n34352 ) ;
assign n34354 =  ( n34239 ) ? ( VREG_3_9 ) : ( n34353 ) ;
assign n34355 =  ( n34238 ) ? ( VREG_3_10 ) : ( n34354 ) ;
assign n34356 =  ( n34237 ) ? ( VREG_3_11 ) : ( n34355 ) ;
assign n34357 =  ( n34236 ) ? ( VREG_3_12 ) : ( n34356 ) ;
assign n34358 =  ( n34235 ) ? ( VREG_3_13 ) : ( n34357 ) ;
assign n34359 =  ( n34234 ) ? ( VREG_3_14 ) : ( n34358 ) ;
assign n34360 =  ( n34233 ) ? ( VREG_3_15 ) : ( n34359 ) ;
assign n34361 =  ( n34232 ) ? ( VREG_4_0 ) : ( n34360 ) ;
assign n34362 =  ( n34231 ) ? ( VREG_4_1 ) : ( n34361 ) ;
assign n34363 =  ( n34230 ) ? ( VREG_4_2 ) : ( n34362 ) ;
assign n34364 =  ( n34229 ) ? ( VREG_4_3 ) : ( n34363 ) ;
assign n34365 =  ( n34228 ) ? ( VREG_4_4 ) : ( n34364 ) ;
assign n34366 =  ( n34227 ) ? ( VREG_4_5 ) : ( n34365 ) ;
assign n34367 =  ( n34226 ) ? ( VREG_4_6 ) : ( n34366 ) ;
assign n34368 =  ( n34225 ) ? ( VREG_4_7 ) : ( n34367 ) ;
assign n34369 =  ( n34224 ) ? ( VREG_4_8 ) : ( n34368 ) ;
assign n34370 =  ( n34223 ) ? ( VREG_4_9 ) : ( n34369 ) ;
assign n34371 =  ( n34222 ) ? ( VREG_4_10 ) : ( n34370 ) ;
assign n34372 =  ( n34221 ) ? ( VREG_4_11 ) : ( n34371 ) ;
assign n34373 =  ( n34220 ) ? ( VREG_4_12 ) : ( n34372 ) ;
assign n34374 =  ( n34219 ) ? ( VREG_4_13 ) : ( n34373 ) ;
assign n34375 =  ( n34218 ) ? ( VREG_4_14 ) : ( n34374 ) ;
assign n34376 =  ( n34217 ) ? ( VREG_4_15 ) : ( n34375 ) ;
assign n34377 =  ( n34216 ) ? ( VREG_5_0 ) : ( n34376 ) ;
assign n34378 =  ( n34215 ) ? ( VREG_5_1 ) : ( n34377 ) ;
assign n34379 =  ( n34214 ) ? ( VREG_5_2 ) : ( n34378 ) ;
assign n34380 =  ( n34213 ) ? ( VREG_5_3 ) : ( n34379 ) ;
assign n34381 =  ( n34212 ) ? ( VREG_5_4 ) : ( n34380 ) ;
assign n34382 =  ( n34211 ) ? ( VREG_5_5 ) : ( n34381 ) ;
assign n34383 =  ( n34210 ) ? ( VREG_5_6 ) : ( n34382 ) ;
assign n34384 =  ( n34209 ) ? ( VREG_5_7 ) : ( n34383 ) ;
assign n34385 =  ( n34208 ) ? ( VREG_5_8 ) : ( n34384 ) ;
assign n34386 =  ( n34207 ) ? ( VREG_5_9 ) : ( n34385 ) ;
assign n34387 =  ( n34206 ) ? ( VREG_5_10 ) : ( n34386 ) ;
assign n34388 =  ( n34205 ) ? ( VREG_5_11 ) : ( n34387 ) ;
assign n34389 =  ( n34204 ) ? ( VREG_5_12 ) : ( n34388 ) ;
assign n34390 =  ( n34203 ) ? ( VREG_5_13 ) : ( n34389 ) ;
assign n34391 =  ( n34202 ) ? ( VREG_5_14 ) : ( n34390 ) ;
assign n34392 =  ( n34201 ) ? ( VREG_5_15 ) : ( n34391 ) ;
assign n34393 =  ( n34200 ) ? ( VREG_6_0 ) : ( n34392 ) ;
assign n34394 =  ( n34199 ) ? ( VREG_6_1 ) : ( n34393 ) ;
assign n34395 =  ( n34198 ) ? ( VREG_6_2 ) : ( n34394 ) ;
assign n34396 =  ( n34197 ) ? ( VREG_6_3 ) : ( n34395 ) ;
assign n34397 =  ( n34196 ) ? ( VREG_6_4 ) : ( n34396 ) ;
assign n34398 =  ( n34195 ) ? ( VREG_6_5 ) : ( n34397 ) ;
assign n34399 =  ( n34194 ) ? ( VREG_6_6 ) : ( n34398 ) ;
assign n34400 =  ( n34193 ) ? ( VREG_6_7 ) : ( n34399 ) ;
assign n34401 =  ( n34192 ) ? ( VREG_6_8 ) : ( n34400 ) ;
assign n34402 =  ( n34191 ) ? ( VREG_6_9 ) : ( n34401 ) ;
assign n34403 =  ( n34190 ) ? ( VREG_6_10 ) : ( n34402 ) ;
assign n34404 =  ( n34189 ) ? ( VREG_6_11 ) : ( n34403 ) ;
assign n34405 =  ( n34188 ) ? ( VREG_6_12 ) : ( n34404 ) ;
assign n34406 =  ( n34187 ) ? ( VREG_6_13 ) : ( n34405 ) ;
assign n34407 =  ( n34186 ) ? ( VREG_6_14 ) : ( n34406 ) ;
assign n34408 =  ( n34185 ) ? ( VREG_6_15 ) : ( n34407 ) ;
assign n34409 =  ( n34184 ) ? ( VREG_7_0 ) : ( n34408 ) ;
assign n34410 =  ( n34183 ) ? ( VREG_7_1 ) : ( n34409 ) ;
assign n34411 =  ( n34182 ) ? ( VREG_7_2 ) : ( n34410 ) ;
assign n34412 =  ( n34181 ) ? ( VREG_7_3 ) : ( n34411 ) ;
assign n34413 =  ( n34180 ) ? ( VREG_7_4 ) : ( n34412 ) ;
assign n34414 =  ( n34179 ) ? ( VREG_7_5 ) : ( n34413 ) ;
assign n34415 =  ( n34178 ) ? ( VREG_7_6 ) : ( n34414 ) ;
assign n34416 =  ( n34177 ) ? ( VREG_7_7 ) : ( n34415 ) ;
assign n34417 =  ( n34176 ) ? ( VREG_7_8 ) : ( n34416 ) ;
assign n34418 =  ( n34175 ) ? ( VREG_7_9 ) : ( n34417 ) ;
assign n34419 =  ( n34174 ) ? ( VREG_7_10 ) : ( n34418 ) ;
assign n34420 =  ( n34173 ) ? ( VREG_7_11 ) : ( n34419 ) ;
assign n34421 =  ( n34172 ) ? ( VREG_7_12 ) : ( n34420 ) ;
assign n34422 =  ( n34171 ) ? ( VREG_7_13 ) : ( n34421 ) ;
assign n34423 =  ( n34170 ) ? ( VREG_7_14 ) : ( n34422 ) ;
assign n34424 =  ( n34169 ) ? ( VREG_7_15 ) : ( n34423 ) ;
assign n34425 =  ( n34168 ) ? ( VREG_8_0 ) : ( n34424 ) ;
assign n34426 =  ( n34167 ) ? ( VREG_8_1 ) : ( n34425 ) ;
assign n34427 =  ( n34166 ) ? ( VREG_8_2 ) : ( n34426 ) ;
assign n34428 =  ( n34165 ) ? ( VREG_8_3 ) : ( n34427 ) ;
assign n34429 =  ( n34164 ) ? ( VREG_8_4 ) : ( n34428 ) ;
assign n34430 =  ( n34163 ) ? ( VREG_8_5 ) : ( n34429 ) ;
assign n34431 =  ( n34162 ) ? ( VREG_8_6 ) : ( n34430 ) ;
assign n34432 =  ( n34161 ) ? ( VREG_8_7 ) : ( n34431 ) ;
assign n34433 =  ( n34160 ) ? ( VREG_8_8 ) : ( n34432 ) ;
assign n34434 =  ( n34159 ) ? ( VREG_8_9 ) : ( n34433 ) ;
assign n34435 =  ( n34158 ) ? ( VREG_8_10 ) : ( n34434 ) ;
assign n34436 =  ( n34157 ) ? ( VREG_8_11 ) : ( n34435 ) ;
assign n34437 =  ( n34156 ) ? ( VREG_8_12 ) : ( n34436 ) ;
assign n34438 =  ( n34155 ) ? ( VREG_8_13 ) : ( n34437 ) ;
assign n34439 =  ( n34154 ) ? ( VREG_8_14 ) : ( n34438 ) ;
assign n34440 =  ( n34153 ) ? ( VREG_8_15 ) : ( n34439 ) ;
assign n34441 =  ( n34152 ) ? ( VREG_9_0 ) : ( n34440 ) ;
assign n34442 =  ( n34151 ) ? ( VREG_9_1 ) : ( n34441 ) ;
assign n34443 =  ( n34150 ) ? ( VREG_9_2 ) : ( n34442 ) ;
assign n34444 =  ( n34149 ) ? ( VREG_9_3 ) : ( n34443 ) ;
assign n34445 =  ( n34148 ) ? ( VREG_9_4 ) : ( n34444 ) ;
assign n34446 =  ( n34147 ) ? ( VREG_9_5 ) : ( n34445 ) ;
assign n34447 =  ( n34146 ) ? ( VREG_9_6 ) : ( n34446 ) ;
assign n34448 =  ( n34145 ) ? ( VREG_9_7 ) : ( n34447 ) ;
assign n34449 =  ( n34144 ) ? ( VREG_9_8 ) : ( n34448 ) ;
assign n34450 =  ( n34143 ) ? ( VREG_9_9 ) : ( n34449 ) ;
assign n34451 =  ( n34142 ) ? ( VREG_9_10 ) : ( n34450 ) ;
assign n34452 =  ( n34141 ) ? ( VREG_9_11 ) : ( n34451 ) ;
assign n34453 =  ( n34140 ) ? ( VREG_9_12 ) : ( n34452 ) ;
assign n34454 =  ( n34139 ) ? ( VREG_9_13 ) : ( n34453 ) ;
assign n34455 =  ( n34138 ) ? ( VREG_9_14 ) : ( n34454 ) ;
assign n34456 =  ( n34137 ) ? ( VREG_9_15 ) : ( n34455 ) ;
assign n34457 =  ( n34136 ) ? ( VREG_10_0 ) : ( n34456 ) ;
assign n34458 =  ( n34135 ) ? ( VREG_10_1 ) : ( n34457 ) ;
assign n34459 =  ( n34134 ) ? ( VREG_10_2 ) : ( n34458 ) ;
assign n34460 =  ( n34133 ) ? ( VREG_10_3 ) : ( n34459 ) ;
assign n34461 =  ( n34132 ) ? ( VREG_10_4 ) : ( n34460 ) ;
assign n34462 =  ( n34131 ) ? ( VREG_10_5 ) : ( n34461 ) ;
assign n34463 =  ( n34130 ) ? ( VREG_10_6 ) : ( n34462 ) ;
assign n34464 =  ( n34129 ) ? ( VREG_10_7 ) : ( n34463 ) ;
assign n34465 =  ( n34128 ) ? ( VREG_10_8 ) : ( n34464 ) ;
assign n34466 =  ( n34127 ) ? ( VREG_10_9 ) : ( n34465 ) ;
assign n34467 =  ( n34126 ) ? ( VREG_10_10 ) : ( n34466 ) ;
assign n34468 =  ( n34125 ) ? ( VREG_10_11 ) : ( n34467 ) ;
assign n34469 =  ( n34124 ) ? ( VREG_10_12 ) : ( n34468 ) ;
assign n34470 =  ( n34123 ) ? ( VREG_10_13 ) : ( n34469 ) ;
assign n34471 =  ( n34122 ) ? ( VREG_10_14 ) : ( n34470 ) ;
assign n34472 =  ( n34121 ) ? ( VREG_10_15 ) : ( n34471 ) ;
assign n34473 =  ( n34120 ) ? ( VREG_11_0 ) : ( n34472 ) ;
assign n34474 =  ( n34119 ) ? ( VREG_11_1 ) : ( n34473 ) ;
assign n34475 =  ( n34118 ) ? ( VREG_11_2 ) : ( n34474 ) ;
assign n34476 =  ( n34117 ) ? ( VREG_11_3 ) : ( n34475 ) ;
assign n34477 =  ( n34116 ) ? ( VREG_11_4 ) : ( n34476 ) ;
assign n34478 =  ( n34115 ) ? ( VREG_11_5 ) : ( n34477 ) ;
assign n34479 =  ( n34114 ) ? ( VREG_11_6 ) : ( n34478 ) ;
assign n34480 =  ( n34113 ) ? ( VREG_11_7 ) : ( n34479 ) ;
assign n34481 =  ( n34112 ) ? ( VREG_11_8 ) : ( n34480 ) ;
assign n34482 =  ( n34111 ) ? ( VREG_11_9 ) : ( n34481 ) ;
assign n34483 =  ( n34110 ) ? ( VREG_11_10 ) : ( n34482 ) ;
assign n34484 =  ( n34109 ) ? ( VREG_11_11 ) : ( n34483 ) ;
assign n34485 =  ( n34108 ) ? ( VREG_11_12 ) : ( n34484 ) ;
assign n34486 =  ( n34107 ) ? ( VREG_11_13 ) : ( n34485 ) ;
assign n34487 =  ( n34106 ) ? ( VREG_11_14 ) : ( n34486 ) ;
assign n34488 =  ( n34105 ) ? ( VREG_11_15 ) : ( n34487 ) ;
assign n34489 =  ( n34104 ) ? ( VREG_12_0 ) : ( n34488 ) ;
assign n34490 =  ( n34103 ) ? ( VREG_12_1 ) : ( n34489 ) ;
assign n34491 =  ( n34102 ) ? ( VREG_12_2 ) : ( n34490 ) ;
assign n34492 =  ( n34101 ) ? ( VREG_12_3 ) : ( n34491 ) ;
assign n34493 =  ( n34100 ) ? ( VREG_12_4 ) : ( n34492 ) ;
assign n34494 =  ( n34099 ) ? ( VREG_12_5 ) : ( n34493 ) ;
assign n34495 =  ( n34098 ) ? ( VREG_12_6 ) : ( n34494 ) ;
assign n34496 =  ( n34097 ) ? ( VREG_12_7 ) : ( n34495 ) ;
assign n34497 =  ( n34096 ) ? ( VREG_12_8 ) : ( n34496 ) ;
assign n34498 =  ( n34095 ) ? ( VREG_12_9 ) : ( n34497 ) ;
assign n34499 =  ( n34094 ) ? ( VREG_12_10 ) : ( n34498 ) ;
assign n34500 =  ( n34093 ) ? ( VREG_12_11 ) : ( n34499 ) ;
assign n34501 =  ( n34092 ) ? ( VREG_12_12 ) : ( n34500 ) ;
assign n34502 =  ( n34091 ) ? ( VREG_12_13 ) : ( n34501 ) ;
assign n34503 =  ( n34090 ) ? ( VREG_12_14 ) : ( n34502 ) ;
assign n34504 =  ( n34089 ) ? ( VREG_12_15 ) : ( n34503 ) ;
assign n34505 =  ( n34088 ) ? ( VREG_13_0 ) : ( n34504 ) ;
assign n34506 =  ( n34087 ) ? ( VREG_13_1 ) : ( n34505 ) ;
assign n34507 =  ( n34086 ) ? ( VREG_13_2 ) : ( n34506 ) ;
assign n34508 =  ( n34085 ) ? ( VREG_13_3 ) : ( n34507 ) ;
assign n34509 =  ( n34084 ) ? ( VREG_13_4 ) : ( n34508 ) ;
assign n34510 =  ( n34083 ) ? ( VREG_13_5 ) : ( n34509 ) ;
assign n34511 =  ( n34082 ) ? ( VREG_13_6 ) : ( n34510 ) ;
assign n34512 =  ( n34081 ) ? ( VREG_13_7 ) : ( n34511 ) ;
assign n34513 =  ( n34080 ) ? ( VREG_13_8 ) : ( n34512 ) ;
assign n34514 =  ( n34079 ) ? ( VREG_13_9 ) : ( n34513 ) ;
assign n34515 =  ( n34078 ) ? ( VREG_13_10 ) : ( n34514 ) ;
assign n34516 =  ( n34077 ) ? ( VREG_13_11 ) : ( n34515 ) ;
assign n34517 =  ( n34076 ) ? ( VREG_13_12 ) : ( n34516 ) ;
assign n34518 =  ( n34075 ) ? ( VREG_13_13 ) : ( n34517 ) ;
assign n34519 =  ( n34074 ) ? ( VREG_13_14 ) : ( n34518 ) ;
assign n34520 =  ( n34073 ) ? ( VREG_13_15 ) : ( n34519 ) ;
assign n34521 =  ( n34072 ) ? ( VREG_14_0 ) : ( n34520 ) ;
assign n34522 =  ( n34071 ) ? ( VREG_14_1 ) : ( n34521 ) ;
assign n34523 =  ( n34070 ) ? ( VREG_14_2 ) : ( n34522 ) ;
assign n34524 =  ( n34069 ) ? ( VREG_14_3 ) : ( n34523 ) ;
assign n34525 =  ( n34068 ) ? ( VREG_14_4 ) : ( n34524 ) ;
assign n34526 =  ( n34067 ) ? ( VREG_14_5 ) : ( n34525 ) ;
assign n34527 =  ( n34066 ) ? ( VREG_14_6 ) : ( n34526 ) ;
assign n34528 =  ( n34065 ) ? ( VREG_14_7 ) : ( n34527 ) ;
assign n34529 =  ( n34064 ) ? ( VREG_14_8 ) : ( n34528 ) ;
assign n34530 =  ( n34063 ) ? ( VREG_14_9 ) : ( n34529 ) ;
assign n34531 =  ( n34062 ) ? ( VREG_14_10 ) : ( n34530 ) ;
assign n34532 =  ( n34061 ) ? ( VREG_14_11 ) : ( n34531 ) ;
assign n34533 =  ( n34060 ) ? ( VREG_14_12 ) : ( n34532 ) ;
assign n34534 =  ( n34059 ) ? ( VREG_14_13 ) : ( n34533 ) ;
assign n34535 =  ( n34058 ) ? ( VREG_14_14 ) : ( n34534 ) ;
assign n34536 =  ( n34057 ) ? ( VREG_14_15 ) : ( n34535 ) ;
assign n34537 =  ( n34056 ) ? ( VREG_15_0 ) : ( n34536 ) ;
assign n34538 =  ( n34055 ) ? ( VREG_15_1 ) : ( n34537 ) ;
assign n34539 =  ( n34054 ) ? ( VREG_15_2 ) : ( n34538 ) ;
assign n34540 =  ( n34053 ) ? ( VREG_15_3 ) : ( n34539 ) ;
assign n34541 =  ( n34052 ) ? ( VREG_15_4 ) : ( n34540 ) ;
assign n34542 =  ( n34051 ) ? ( VREG_15_5 ) : ( n34541 ) ;
assign n34543 =  ( n34050 ) ? ( VREG_15_6 ) : ( n34542 ) ;
assign n34544 =  ( n34049 ) ? ( VREG_15_7 ) : ( n34543 ) ;
assign n34545 =  ( n34048 ) ? ( VREG_15_8 ) : ( n34544 ) ;
assign n34546 =  ( n34047 ) ? ( VREG_15_9 ) : ( n34545 ) ;
assign n34547 =  ( n34046 ) ? ( VREG_15_10 ) : ( n34546 ) ;
assign n34548 =  ( n34045 ) ? ( VREG_15_11 ) : ( n34547 ) ;
assign n34549 =  ( n34044 ) ? ( VREG_15_12 ) : ( n34548 ) ;
assign n34550 =  ( n34043 ) ? ( VREG_15_13 ) : ( n34549 ) ;
assign n34551 =  ( n34042 ) ? ( VREG_15_14 ) : ( n34550 ) ;
assign n34552 =  ( n34041 ) ? ( VREG_15_15 ) : ( n34551 ) ;
assign n34553 =  ( n34040 ) ? ( VREG_16_0 ) : ( n34552 ) ;
assign n34554 =  ( n34039 ) ? ( VREG_16_1 ) : ( n34553 ) ;
assign n34555 =  ( n34038 ) ? ( VREG_16_2 ) : ( n34554 ) ;
assign n34556 =  ( n34037 ) ? ( VREG_16_3 ) : ( n34555 ) ;
assign n34557 =  ( n34036 ) ? ( VREG_16_4 ) : ( n34556 ) ;
assign n34558 =  ( n34035 ) ? ( VREG_16_5 ) : ( n34557 ) ;
assign n34559 =  ( n34034 ) ? ( VREG_16_6 ) : ( n34558 ) ;
assign n34560 =  ( n34033 ) ? ( VREG_16_7 ) : ( n34559 ) ;
assign n34561 =  ( n34032 ) ? ( VREG_16_8 ) : ( n34560 ) ;
assign n34562 =  ( n34031 ) ? ( VREG_16_9 ) : ( n34561 ) ;
assign n34563 =  ( n34030 ) ? ( VREG_16_10 ) : ( n34562 ) ;
assign n34564 =  ( n34029 ) ? ( VREG_16_11 ) : ( n34563 ) ;
assign n34565 =  ( n34028 ) ? ( VREG_16_12 ) : ( n34564 ) ;
assign n34566 =  ( n34027 ) ? ( VREG_16_13 ) : ( n34565 ) ;
assign n34567 =  ( n34026 ) ? ( VREG_16_14 ) : ( n34566 ) ;
assign n34568 =  ( n34025 ) ? ( VREG_16_15 ) : ( n34567 ) ;
assign n34569 =  ( n34024 ) ? ( VREG_17_0 ) : ( n34568 ) ;
assign n34570 =  ( n34023 ) ? ( VREG_17_1 ) : ( n34569 ) ;
assign n34571 =  ( n34022 ) ? ( VREG_17_2 ) : ( n34570 ) ;
assign n34572 =  ( n34021 ) ? ( VREG_17_3 ) : ( n34571 ) ;
assign n34573 =  ( n34020 ) ? ( VREG_17_4 ) : ( n34572 ) ;
assign n34574 =  ( n34019 ) ? ( VREG_17_5 ) : ( n34573 ) ;
assign n34575 =  ( n34018 ) ? ( VREG_17_6 ) : ( n34574 ) ;
assign n34576 =  ( n34017 ) ? ( VREG_17_7 ) : ( n34575 ) ;
assign n34577 =  ( n34016 ) ? ( VREG_17_8 ) : ( n34576 ) ;
assign n34578 =  ( n34015 ) ? ( VREG_17_9 ) : ( n34577 ) ;
assign n34579 =  ( n34014 ) ? ( VREG_17_10 ) : ( n34578 ) ;
assign n34580 =  ( n34013 ) ? ( VREG_17_11 ) : ( n34579 ) ;
assign n34581 =  ( n34012 ) ? ( VREG_17_12 ) : ( n34580 ) ;
assign n34582 =  ( n34011 ) ? ( VREG_17_13 ) : ( n34581 ) ;
assign n34583 =  ( n34010 ) ? ( VREG_17_14 ) : ( n34582 ) ;
assign n34584 =  ( n34009 ) ? ( VREG_17_15 ) : ( n34583 ) ;
assign n34585 =  ( n34008 ) ? ( VREG_18_0 ) : ( n34584 ) ;
assign n34586 =  ( n34007 ) ? ( VREG_18_1 ) : ( n34585 ) ;
assign n34587 =  ( n34006 ) ? ( VREG_18_2 ) : ( n34586 ) ;
assign n34588 =  ( n34005 ) ? ( VREG_18_3 ) : ( n34587 ) ;
assign n34589 =  ( n34004 ) ? ( VREG_18_4 ) : ( n34588 ) ;
assign n34590 =  ( n34003 ) ? ( VREG_18_5 ) : ( n34589 ) ;
assign n34591 =  ( n34002 ) ? ( VREG_18_6 ) : ( n34590 ) ;
assign n34592 =  ( n34001 ) ? ( VREG_18_7 ) : ( n34591 ) ;
assign n34593 =  ( n34000 ) ? ( VREG_18_8 ) : ( n34592 ) ;
assign n34594 =  ( n33999 ) ? ( VREG_18_9 ) : ( n34593 ) ;
assign n34595 =  ( n33998 ) ? ( VREG_18_10 ) : ( n34594 ) ;
assign n34596 =  ( n33997 ) ? ( VREG_18_11 ) : ( n34595 ) ;
assign n34597 =  ( n33996 ) ? ( VREG_18_12 ) : ( n34596 ) ;
assign n34598 =  ( n33995 ) ? ( VREG_18_13 ) : ( n34597 ) ;
assign n34599 =  ( n33994 ) ? ( VREG_18_14 ) : ( n34598 ) ;
assign n34600 =  ( n33993 ) ? ( VREG_18_15 ) : ( n34599 ) ;
assign n34601 =  ( n33992 ) ? ( VREG_19_0 ) : ( n34600 ) ;
assign n34602 =  ( n33991 ) ? ( VREG_19_1 ) : ( n34601 ) ;
assign n34603 =  ( n33990 ) ? ( VREG_19_2 ) : ( n34602 ) ;
assign n34604 =  ( n33989 ) ? ( VREG_19_3 ) : ( n34603 ) ;
assign n34605 =  ( n33988 ) ? ( VREG_19_4 ) : ( n34604 ) ;
assign n34606 =  ( n33987 ) ? ( VREG_19_5 ) : ( n34605 ) ;
assign n34607 =  ( n33986 ) ? ( VREG_19_6 ) : ( n34606 ) ;
assign n34608 =  ( n33985 ) ? ( VREG_19_7 ) : ( n34607 ) ;
assign n34609 =  ( n33984 ) ? ( VREG_19_8 ) : ( n34608 ) ;
assign n34610 =  ( n33983 ) ? ( VREG_19_9 ) : ( n34609 ) ;
assign n34611 =  ( n33982 ) ? ( VREG_19_10 ) : ( n34610 ) ;
assign n34612 =  ( n33981 ) ? ( VREG_19_11 ) : ( n34611 ) ;
assign n34613 =  ( n33980 ) ? ( VREG_19_12 ) : ( n34612 ) ;
assign n34614 =  ( n33979 ) ? ( VREG_19_13 ) : ( n34613 ) ;
assign n34615 =  ( n33978 ) ? ( VREG_19_14 ) : ( n34614 ) ;
assign n34616 =  ( n33977 ) ? ( VREG_19_15 ) : ( n34615 ) ;
assign n34617 =  ( n33976 ) ? ( VREG_20_0 ) : ( n34616 ) ;
assign n34618 =  ( n33975 ) ? ( VREG_20_1 ) : ( n34617 ) ;
assign n34619 =  ( n33974 ) ? ( VREG_20_2 ) : ( n34618 ) ;
assign n34620 =  ( n33973 ) ? ( VREG_20_3 ) : ( n34619 ) ;
assign n34621 =  ( n33972 ) ? ( VREG_20_4 ) : ( n34620 ) ;
assign n34622 =  ( n33971 ) ? ( VREG_20_5 ) : ( n34621 ) ;
assign n34623 =  ( n33970 ) ? ( VREG_20_6 ) : ( n34622 ) ;
assign n34624 =  ( n33969 ) ? ( VREG_20_7 ) : ( n34623 ) ;
assign n34625 =  ( n33968 ) ? ( VREG_20_8 ) : ( n34624 ) ;
assign n34626 =  ( n33967 ) ? ( VREG_20_9 ) : ( n34625 ) ;
assign n34627 =  ( n33966 ) ? ( VREG_20_10 ) : ( n34626 ) ;
assign n34628 =  ( n33965 ) ? ( VREG_20_11 ) : ( n34627 ) ;
assign n34629 =  ( n33964 ) ? ( VREG_20_12 ) : ( n34628 ) ;
assign n34630 =  ( n33963 ) ? ( VREG_20_13 ) : ( n34629 ) ;
assign n34631 =  ( n33962 ) ? ( VREG_20_14 ) : ( n34630 ) ;
assign n34632 =  ( n33961 ) ? ( VREG_20_15 ) : ( n34631 ) ;
assign n34633 =  ( n33960 ) ? ( VREG_21_0 ) : ( n34632 ) ;
assign n34634 =  ( n33959 ) ? ( VREG_21_1 ) : ( n34633 ) ;
assign n34635 =  ( n33958 ) ? ( VREG_21_2 ) : ( n34634 ) ;
assign n34636 =  ( n33957 ) ? ( VREG_21_3 ) : ( n34635 ) ;
assign n34637 =  ( n33956 ) ? ( VREG_21_4 ) : ( n34636 ) ;
assign n34638 =  ( n33955 ) ? ( VREG_21_5 ) : ( n34637 ) ;
assign n34639 =  ( n33954 ) ? ( VREG_21_6 ) : ( n34638 ) ;
assign n34640 =  ( n33953 ) ? ( VREG_21_7 ) : ( n34639 ) ;
assign n34641 =  ( n33952 ) ? ( VREG_21_8 ) : ( n34640 ) ;
assign n34642 =  ( n33951 ) ? ( VREG_21_9 ) : ( n34641 ) ;
assign n34643 =  ( n33950 ) ? ( VREG_21_10 ) : ( n34642 ) ;
assign n34644 =  ( n33949 ) ? ( VREG_21_11 ) : ( n34643 ) ;
assign n34645 =  ( n33948 ) ? ( VREG_21_12 ) : ( n34644 ) ;
assign n34646 =  ( n33947 ) ? ( VREG_21_13 ) : ( n34645 ) ;
assign n34647 =  ( n33946 ) ? ( VREG_21_14 ) : ( n34646 ) ;
assign n34648 =  ( n33945 ) ? ( VREG_21_15 ) : ( n34647 ) ;
assign n34649 =  ( n33944 ) ? ( VREG_22_0 ) : ( n34648 ) ;
assign n34650 =  ( n33943 ) ? ( VREG_22_1 ) : ( n34649 ) ;
assign n34651 =  ( n33942 ) ? ( VREG_22_2 ) : ( n34650 ) ;
assign n34652 =  ( n33941 ) ? ( VREG_22_3 ) : ( n34651 ) ;
assign n34653 =  ( n33940 ) ? ( VREG_22_4 ) : ( n34652 ) ;
assign n34654 =  ( n33939 ) ? ( VREG_22_5 ) : ( n34653 ) ;
assign n34655 =  ( n33938 ) ? ( VREG_22_6 ) : ( n34654 ) ;
assign n34656 =  ( n33937 ) ? ( VREG_22_7 ) : ( n34655 ) ;
assign n34657 =  ( n33936 ) ? ( VREG_22_8 ) : ( n34656 ) ;
assign n34658 =  ( n33935 ) ? ( VREG_22_9 ) : ( n34657 ) ;
assign n34659 =  ( n33934 ) ? ( VREG_22_10 ) : ( n34658 ) ;
assign n34660 =  ( n33933 ) ? ( VREG_22_11 ) : ( n34659 ) ;
assign n34661 =  ( n33932 ) ? ( VREG_22_12 ) : ( n34660 ) ;
assign n34662 =  ( n33931 ) ? ( VREG_22_13 ) : ( n34661 ) ;
assign n34663 =  ( n33930 ) ? ( VREG_22_14 ) : ( n34662 ) ;
assign n34664 =  ( n33929 ) ? ( VREG_22_15 ) : ( n34663 ) ;
assign n34665 =  ( n33928 ) ? ( VREG_23_0 ) : ( n34664 ) ;
assign n34666 =  ( n33927 ) ? ( VREG_23_1 ) : ( n34665 ) ;
assign n34667 =  ( n33926 ) ? ( VREG_23_2 ) : ( n34666 ) ;
assign n34668 =  ( n33925 ) ? ( VREG_23_3 ) : ( n34667 ) ;
assign n34669 =  ( n33924 ) ? ( VREG_23_4 ) : ( n34668 ) ;
assign n34670 =  ( n33923 ) ? ( VREG_23_5 ) : ( n34669 ) ;
assign n34671 =  ( n33922 ) ? ( VREG_23_6 ) : ( n34670 ) ;
assign n34672 =  ( n33921 ) ? ( VREG_23_7 ) : ( n34671 ) ;
assign n34673 =  ( n33920 ) ? ( VREG_23_8 ) : ( n34672 ) ;
assign n34674 =  ( n33919 ) ? ( VREG_23_9 ) : ( n34673 ) ;
assign n34675 =  ( n33918 ) ? ( VREG_23_10 ) : ( n34674 ) ;
assign n34676 =  ( n33917 ) ? ( VREG_23_11 ) : ( n34675 ) ;
assign n34677 =  ( n33916 ) ? ( VREG_23_12 ) : ( n34676 ) ;
assign n34678 =  ( n33915 ) ? ( VREG_23_13 ) : ( n34677 ) ;
assign n34679 =  ( n33914 ) ? ( VREG_23_14 ) : ( n34678 ) ;
assign n34680 =  ( n33913 ) ? ( VREG_23_15 ) : ( n34679 ) ;
assign n34681 =  ( n33912 ) ? ( VREG_24_0 ) : ( n34680 ) ;
assign n34682 =  ( n33911 ) ? ( VREG_24_1 ) : ( n34681 ) ;
assign n34683 =  ( n33910 ) ? ( VREG_24_2 ) : ( n34682 ) ;
assign n34684 =  ( n33909 ) ? ( VREG_24_3 ) : ( n34683 ) ;
assign n34685 =  ( n33908 ) ? ( VREG_24_4 ) : ( n34684 ) ;
assign n34686 =  ( n33907 ) ? ( VREG_24_5 ) : ( n34685 ) ;
assign n34687 =  ( n33906 ) ? ( VREG_24_6 ) : ( n34686 ) ;
assign n34688 =  ( n33905 ) ? ( VREG_24_7 ) : ( n34687 ) ;
assign n34689 =  ( n33904 ) ? ( VREG_24_8 ) : ( n34688 ) ;
assign n34690 =  ( n33903 ) ? ( VREG_24_9 ) : ( n34689 ) ;
assign n34691 =  ( n33902 ) ? ( VREG_24_10 ) : ( n34690 ) ;
assign n34692 =  ( n33901 ) ? ( VREG_24_11 ) : ( n34691 ) ;
assign n34693 =  ( n33900 ) ? ( VREG_24_12 ) : ( n34692 ) ;
assign n34694 =  ( n33899 ) ? ( VREG_24_13 ) : ( n34693 ) ;
assign n34695 =  ( n33898 ) ? ( VREG_24_14 ) : ( n34694 ) ;
assign n34696 =  ( n33897 ) ? ( VREG_24_15 ) : ( n34695 ) ;
assign n34697 =  ( n33896 ) ? ( VREG_25_0 ) : ( n34696 ) ;
assign n34698 =  ( n33895 ) ? ( VREG_25_1 ) : ( n34697 ) ;
assign n34699 =  ( n33894 ) ? ( VREG_25_2 ) : ( n34698 ) ;
assign n34700 =  ( n33893 ) ? ( VREG_25_3 ) : ( n34699 ) ;
assign n34701 =  ( n33892 ) ? ( VREG_25_4 ) : ( n34700 ) ;
assign n34702 =  ( n33891 ) ? ( VREG_25_5 ) : ( n34701 ) ;
assign n34703 =  ( n33890 ) ? ( VREG_25_6 ) : ( n34702 ) ;
assign n34704 =  ( n33889 ) ? ( VREG_25_7 ) : ( n34703 ) ;
assign n34705 =  ( n33888 ) ? ( VREG_25_8 ) : ( n34704 ) ;
assign n34706 =  ( n33887 ) ? ( VREG_25_9 ) : ( n34705 ) ;
assign n34707 =  ( n33886 ) ? ( VREG_25_10 ) : ( n34706 ) ;
assign n34708 =  ( n33885 ) ? ( VREG_25_11 ) : ( n34707 ) ;
assign n34709 =  ( n33884 ) ? ( VREG_25_12 ) : ( n34708 ) ;
assign n34710 =  ( n33883 ) ? ( VREG_25_13 ) : ( n34709 ) ;
assign n34711 =  ( n33882 ) ? ( VREG_25_14 ) : ( n34710 ) ;
assign n34712 =  ( n33881 ) ? ( VREG_25_15 ) : ( n34711 ) ;
assign n34713 =  ( n33880 ) ? ( VREG_26_0 ) : ( n34712 ) ;
assign n34714 =  ( n33879 ) ? ( VREG_26_1 ) : ( n34713 ) ;
assign n34715 =  ( n33878 ) ? ( VREG_26_2 ) : ( n34714 ) ;
assign n34716 =  ( n33877 ) ? ( VREG_26_3 ) : ( n34715 ) ;
assign n34717 =  ( n33876 ) ? ( VREG_26_4 ) : ( n34716 ) ;
assign n34718 =  ( n33875 ) ? ( VREG_26_5 ) : ( n34717 ) ;
assign n34719 =  ( n33874 ) ? ( VREG_26_6 ) : ( n34718 ) ;
assign n34720 =  ( n33873 ) ? ( VREG_26_7 ) : ( n34719 ) ;
assign n34721 =  ( n33872 ) ? ( VREG_26_8 ) : ( n34720 ) ;
assign n34722 =  ( n33871 ) ? ( VREG_26_9 ) : ( n34721 ) ;
assign n34723 =  ( n33870 ) ? ( VREG_26_10 ) : ( n34722 ) ;
assign n34724 =  ( n33869 ) ? ( VREG_26_11 ) : ( n34723 ) ;
assign n34725 =  ( n33868 ) ? ( VREG_26_12 ) : ( n34724 ) ;
assign n34726 =  ( n33867 ) ? ( VREG_26_13 ) : ( n34725 ) ;
assign n34727 =  ( n33866 ) ? ( VREG_26_14 ) : ( n34726 ) ;
assign n34728 =  ( n33865 ) ? ( VREG_26_15 ) : ( n34727 ) ;
assign n34729 =  ( n33864 ) ? ( VREG_27_0 ) : ( n34728 ) ;
assign n34730 =  ( n33863 ) ? ( VREG_27_1 ) : ( n34729 ) ;
assign n34731 =  ( n33862 ) ? ( VREG_27_2 ) : ( n34730 ) ;
assign n34732 =  ( n33861 ) ? ( VREG_27_3 ) : ( n34731 ) ;
assign n34733 =  ( n33860 ) ? ( VREG_27_4 ) : ( n34732 ) ;
assign n34734 =  ( n33859 ) ? ( VREG_27_5 ) : ( n34733 ) ;
assign n34735 =  ( n33858 ) ? ( VREG_27_6 ) : ( n34734 ) ;
assign n34736 =  ( n33857 ) ? ( VREG_27_7 ) : ( n34735 ) ;
assign n34737 =  ( n33856 ) ? ( VREG_27_8 ) : ( n34736 ) ;
assign n34738 =  ( n33855 ) ? ( VREG_27_9 ) : ( n34737 ) ;
assign n34739 =  ( n33854 ) ? ( VREG_27_10 ) : ( n34738 ) ;
assign n34740 =  ( n33853 ) ? ( VREG_27_11 ) : ( n34739 ) ;
assign n34741 =  ( n33852 ) ? ( VREG_27_12 ) : ( n34740 ) ;
assign n34742 =  ( n33851 ) ? ( VREG_27_13 ) : ( n34741 ) ;
assign n34743 =  ( n33850 ) ? ( VREG_27_14 ) : ( n34742 ) ;
assign n34744 =  ( n33849 ) ? ( VREG_27_15 ) : ( n34743 ) ;
assign n34745 =  ( n33848 ) ? ( VREG_28_0 ) : ( n34744 ) ;
assign n34746 =  ( n33847 ) ? ( VREG_28_1 ) : ( n34745 ) ;
assign n34747 =  ( n33846 ) ? ( VREG_28_2 ) : ( n34746 ) ;
assign n34748 =  ( n33845 ) ? ( VREG_28_3 ) : ( n34747 ) ;
assign n34749 =  ( n33844 ) ? ( VREG_28_4 ) : ( n34748 ) ;
assign n34750 =  ( n33843 ) ? ( VREG_28_5 ) : ( n34749 ) ;
assign n34751 =  ( n33842 ) ? ( VREG_28_6 ) : ( n34750 ) ;
assign n34752 =  ( n33841 ) ? ( VREG_28_7 ) : ( n34751 ) ;
assign n34753 =  ( n33840 ) ? ( VREG_28_8 ) : ( n34752 ) ;
assign n34754 =  ( n33839 ) ? ( VREG_28_9 ) : ( n34753 ) ;
assign n34755 =  ( n33838 ) ? ( VREG_28_10 ) : ( n34754 ) ;
assign n34756 =  ( n33837 ) ? ( VREG_28_11 ) : ( n34755 ) ;
assign n34757 =  ( n33836 ) ? ( VREG_28_12 ) : ( n34756 ) ;
assign n34758 =  ( n33835 ) ? ( VREG_28_13 ) : ( n34757 ) ;
assign n34759 =  ( n33834 ) ? ( VREG_28_14 ) : ( n34758 ) ;
assign n34760 =  ( n33833 ) ? ( VREG_28_15 ) : ( n34759 ) ;
assign n34761 =  ( n33832 ) ? ( VREG_29_0 ) : ( n34760 ) ;
assign n34762 =  ( n33831 ) ? ( VREG_29_1 ) : ( n34761 ) ;
assign n34763 =  ( n33830 ) ? ( VREG_29_2 ) : ( n34762 ) ;
assign n34764 =  ( n33829 ) ? ( VREG_29_3 ) : ( n34763 ) ;
assign n34765 =  ( n33828 ) ? ( VREG_29_4 ) : ( n34764 ) ;
assign n34766 =  ( n33827 ) ? ( VREG_29_5 ) : ( n34765 ) ;
assign n34767 =  ( n33826 ) ? ( VREG_29_6 ) : ( n34766 ) ;
assign n34768 =  ( n33825 ) ? ( VREG_29_7 ) : ( n34767 ) ;
assign n34769 =  ( n33824 ) ? ( VREG_29_8 ) : ( n34768 ) ;
assign n34770 =  ( n33823 ) ? ( VREG_29_9 ) : ( n34769 ) ;
assign n34771 =  ( n33822 ) ? ( VREG_29_10 ) : ( n34770 ) ;
assign n34772 =  ( n33821 ) ? ( VREG_29_11 ) : ( n34771 ) ;
assign n34773 =  ( n33820 ) ? ( VREG_29_12 ) : ( n34772 ) ;
assign n34774 =  ( n33819 ) ? ( VREG_29_13 ) : ( n34773 ) ;
assign n34775 =  ( n33818 ) ? ( VREG_29_14 ) : ( n34774 ) ;
assign n34776 =  ( n33817 ) ? ( VREG_29_15 ) : ( n34775 ) ;
assign n34777 =  ( n33816 ) ? ( VREG_30_0 ) : ( n34776 ) ;
assign n34778 =  ( n33815 ) ? ( VREG_30_1 ) : ( n34777 ) ;
assign n34779 =  ( n33814 ) ? ( VREG_30_2 ) : ( n34778 ) ;
assign n34780 =  ( n33813 ) ? ( VREG_30_3 ) : ( n34779 ) ;
assign n34781 =  ( n33812 ) ? ( VREG_30_4 ) : ( n34780 ) ;
assign n34782 =  ( n33811 ) ? ( VREG_30_5 ) : ( n34781 ) ;
assign n34783 =  ( n33810 ) ? ( VREG_30_6 ) : ( n34782 ) ;
assign n34784 =  ( n33809 ) ? ( VREG_30_7 ) : ( n34783 ) ;
assign n34785 =  ( n33808 ) ? ( VREG_30_8 ) : ( n34784 ) ;
assign n34786 =  ( n33807 ) ? ( VREG_30_9 ) : ( n34785 ) ;
assign n34787 =  ( n33806 ) ? ( VREG_30_10 ) : ( n34786 ) ;
assign n34788 =  ( n33805 ) ? ( VREG_30_11 ) : ( n34787 ) ;
assign n34789 =  ( n33804 ) ? ( VREG_30_12 ) : ( n34788 ) ;
assign n34790 =  ( n33803 ) ? ( VREG_30_13 ) : ( n34789 ) ;
assign n34791 =  ( n33802 ) ? ( VREG_30_14 ) : ( n34790 ) ;
assign n34792 =  ( n33801 ) ? ( VREG_30_15 ) : ( n34791 ) ;
assign n34793 =  ( n33800 ) ? ( VREG_31_0 ) : ( n34792 ) ;
assign n34794 =  ( n33799 ) ? ( VREG_31_1 ) : ( n34793 ) ;
assign n34795 =  ( n33798 ) ? ( VREG_31_2 ) : ( n34794 ) ;
assign n34796 =  ( n33797 ) ? ( VREG_31_3 ) : ( n34795 ) ;
assign n34797 =  ( n33796 ) ? ( VREG_31_4 ) : ( n34796 ) ;
assign n34798 =  ( n33795 ) ? ( VREG_31_5 ) : ( n34797 ) ;
assign n34799 =  ( n33794 ) ? ( VREG_31_6 ) : ( n34798 ) ;
assign n34800 =  ( n33793 ) ? ( VREG_31_7 ) : ( n34799 ) ;
assign n34801 =  ( n33792 ) ? ( VREG_31_8 ) : ( n34800 ) ;
assign n34802 =  ( n33791 ) ? ( VREG_31_9 ) : ( n34801 ) ;
assign n34803 =  ( n33790 ) ? ( VREG_31_10 ) : ( n34802 ) ;
assign n34804 =  ( n33789 ) ? ( VREG_31_11 ) : ( n34803 ) ;
assign n34805 =  ( n33788 ) ? ( VREG_31_12 ) : ( n34804 ) ;
assign n34806 =  ( n33787 ) ? ( VREG_31_13 ) : ( n34805 ) ;
assign n34807 =  ( n33786 ) ? ( VREG_31_14 ) : ( n34806 ) ;
assign n34808 =  ( n33785 ) ? ( VREG_31_15 ) : ( n34807 ) ;
assign n34809 =  ( n33774 ) + ( n34808 )  ;
assign n34810 =  ( n33774 ) - ( n34808 )  ;
assign n34811 =  ( n33774 ) & ( n34808 )  ;
assign n34812 =  ( n33774 ) | ( n34808 )  ;
assign n34813 =  ( ( n33774 ) * ( n34808 ))  ;
assign n34814 =  ( n148 ) ? ( n34813 ) : ( VREG_0_9 ) ;
assign n34815 =  ( n146 ) ? ( n34812 ) : ( n34814 ) ;
assign n34816 =  ( n144 ) ? ( n34811 ) : ( n34815 ) ;
assign n34817 =  ( n142 ) ? ( n34810 ) : ( n34816 ) ;
assign n34818 =  ( n10 ) ? ( n34809 ) : ( n34817 ) ;
assign n34819 = n3030[9:9] ;
assign n34820 =  ( n34819 ) == ( 1'd0 )  ;
assign n34821 =  ( n34820 ) ? ( VREG_0_9 ) : ( n33784 ) ;
assign n34822 =  ( n34820 ) ? ( VREG_0_9 ) : ( n34818 ) ;
assign n34823 =  ( n3034 ) ? ( n34822 ) : ( VREG_0_9 ) ;
assign n34824 =  ( n2965 ) ? ( n34821 ) : ( n34823 ) ;
assign n34825 =  ( n1930 ) ? ( n34818 ) : ( n34824 ) ;
assign n34826 =  ( n879 ) ? ( n33784 ) : ( n34825 ) ;
assign n34827 =  ( n33774 ) + ( n164 )  ;
assign n34828 =  ( n33774 ) - ( n164 )  ;
assign n34829 =  ( n33774 ) & ( n164 )  ;
assign n34830 =  ( n33774 ) | ( n164 )  ;
assign n34831 =  ( ( n33774 ) * ( n164 ))  ;
assign n34832 =  ( n172 ) ? ( n34831 ) : ( VREG_0_9 ) ;
assign n34833 =  ( n170 ) ? ( n34830 ) : ( n34832 ) ;
assign n34834 =  ( n168 ) ? ( n34829 ) : ( n34833 ) ;
assign n34835 =  ( n166 ) ? ( n34828 ) : ( n34834 ) ;
assign n34836 =  ( n162 ) ? ( n34827 ) : ( n34835 ) ;
assign n34837 =  ( n33774 ) + ( n180 )  ;
assign n34838 =  ( n33774 ) - ( n180 )  ;
assign n34839 =  ( n33774 ) & ( n180 )  ;
assign n34840 =  ( n33774 ) | ( n180 )  ;
assign n34841 =  ( ( n33774 ) * ( n180 ))  ;
assign n34842 =  ( n172 ) ? ( n34841 ) : ( VREG_0_9 ) ;
assign n34843 =  ( n170 ) ? ( n34840 ) : ( n34842 ) ;
assign n34844 =  ( n168 ) ? ( n34839 ) : ( n34843 ) ;
assign n34845 =  ( n166 ) ? ( n34838 ) : ( n34844 ) ;
assign n34846 =  ( n162 ) ? ( n34837 ) : ( n34845 ) ;
assign n34847 =  ( n34820 ) ? ( VREG_0_9 ) : ( n34846 ) ;
assign n34848 =  ( n3051 ) ? ( n34847 ) : ( VREG_0_9 ) ;
assign n34849 =  ( n3040 ) ? ( n34836 ) : ( n34848 ) ;
assign n34850 =  ( n192 ) ? ( VREG_0_9 ) : ( VREG_0_9 ) ;
assign n34851 =  ( n157 ) ? ( n34849 ) : ( n34850 ) ;
assign n34852 =  ( n6 ) ? ( n34826 ) : ( n34851 ) ;
assign n34853 =  ( n4 ) ? ( n34852 ) : ( VREG_0_9 ) ;
assign n34854 =  ( n148 ) ? ( n1924 ) : ( VREG_10_0 ) ;
assign n34855 =  ( n146 ) ? ( n1923 ) : ( n34854 ) ;
assign n34856 =  ( n144 ) ? ( n1922 ) : ( n34855 ) ;
assign n34857 =  ( n142 ) ? ( n1921 ) : ( n34856 ) ;
assign n34858 =  ( n10 ) ? ( n1920 ) : ( n34857 ) ;
assign n34859 =  ( n148 ) ? ( n2959 ) : ( VREG_10_0 ) ;
assign n34860 =  ( n146 ) ? ( n2958 ) : ( n34859 ) ;
assign n34861 =  ( n144 ) ? ( n2957 ) : ( n34860 ) ;
assign n34862 =  ( n142 ) ? ( n2956 ) : ( n34861 ) ;
assign n34863 =  ( n10 ) ? ( n2955 ) : ( n34862 ) ;
assign n34864 =  ( n3032 ) ? ( VREG_10_0 ) : ( n34858 ) ;
assign n34865 =  ( n3032 ) ? ( VREG_10_0 ) : ( n34863 ) ;
assign n34866 =  ( n3034 ) ? ( n34865 ) : ( VREG_10_0 ) ;
assign n34867 =  ( n2965 ) ? ( n34864 ) : ( n34866 ) ;
assign n34868 =  ( n1930 ) ? ( n34863 ) : ( n34867 ) ;
assign n34869 =  ( n879 ) ? ( n34858 ) : ( n34868 ) ;
assign n34870 =  ( n172 ) ? ( n3045 ) : ( VREG_10_0 ) ;
assign n34871 =  ( n170 ) ? ( n3044 ) : ( n34870 ) ;
assign n34872 =  ( n168 ) ? ( n3043 ) : ( n34871 ) ;
assign n34873 =  ( n166 ) ? ( n3042 ) : ( n34872 ) ;
assign n34874 =  ( n162 ) ? ( n3041 ) : ( n34873 ) ;
assign n34875 =  ( n172 ) ? ( n3056 ) : ( VREG_10_0 ) ;
assign n34876 =  ( n170 ) ? ( n3055 ) : ( n34875 ) ;
assign n34877 =  ( n168 ) ? ( n3054 ) : ( n34876 ) ;
assign n34878 =  ( n166 ) ? ( n3053 ) : ( n34877 ) ;
assign n34879 =  ( n162 ) ? ( n3052 ) : ( n34878 ) ;
assign n34880 =  ( n3032 ) ? ( VREG_10_0 ) : ( n34879 ) ;
assign n34881 =  ( n3051 ) ? ( n34880 ) : ( VREG_10_0 ) ;
assign n34882 =  ( n3040 ) ? ( n34874 ) : ( n34881 ) ;
assign n34883 =  ( n192 ) ? ( VREG_10_0 ) : ( VREG_10_0 ) ;
assign n34884 =  ( n157 ) ? ( n34882 ) : ( n34883 ) ;
assign n34885 =  ( n6 ) ? ( n34869 ) : ( n34884 ) ;
assign n34886 =  ( n219 ) ? ( n34885 ) : ( VREG_10_0 ) ;
assign n34887 =  ( n148 ) ? ( n4113 ) : ( VREG_10_1 ) ;
assign n34888 =  ( n146 ) ? ( n4112 ) : ( n34887 ) ;
assign n34889 =  ( n144 ) ? ( n4111 ) : ( n34888 ) ;
assign n34890 =  ( n142 ) ? ( n4110 ) : ( n34889 ) ;
assign n34891 =  ( n10 ) ? ( n4109 ) : ( n34890 ) ;
assign n34892 =  ( n148 ) ? ( n5147 ) : ( VREG_10_1 ) ;
assign n34893 =  ( n146 ) ? ( n5146 ) : ( n34892 ) ;
assign n34894 =  ( n144 ) ? ( n5145 ) : ( n34893 ) ;
assign n34895 =  ( n142 ) ? ( n5144 ) : ( n34894 ) ;
assign n34896 =  ( n10 ) ? ( n5143 ) : ( n34895 ) ;
assign n34897 =  ( n5154 ) ? ( VREG_10_1 ) : ( n34891 ) ;
assign n34898 =  ( n5154 ) ? ( VREG_10_1 ) : ( n34896 ) ;
assign n34899 =  ( n3034 ) ? ( n34898 ) : ( VREG_10_1 ) ;
assign n34900 =  ( n2965 ) ? ( n34897 ) : ( n34899 ) ;
assign n34901 =  ( n1930 ) ? ( n34896 ) : ( n34900 ) ;
assign n34902 =  ( n879 ) ? ( n34891 ) : ( n34901 ) ;
assign n34903 =  ( n172 ) ? ( n5165 ) : ( VREG_10_1 ) ;
assign n34904 =  ( n170 ) ? ( n5164 ) : ( n34903 ) ;
assign n34905 =  ( n168 ) ? ( n5163 ) : ( n34904 ) ;
assign n34906 =  ( n166 ) ? ( n5162 ) : ( n34905 ) ;
assign n34907 =  ( n162 ) ? ( n5161 ) : ( n34906 ) ;
assign n34908 =  ( n172 ) ? ( n5175 ) : ( VREG_10_1 ) ;
assign n34909 =  ( n170 ) ? ( n5174 ) : ( n34908 ) ;
assign n34910 =  ( n168 ) ? ( n5173 ) : ( n34909 ) ;
assign n34911 =  ( n166 ) ? ( n5172 ) : ( n34910 ) ;
assign n34912 =  ( n162 ) ? ( n5171 ) : ( n34911 ) ;
assign n34913 =  ( n5154 ) ? ( VREG_10_1 ) : ( n34912 ) ;
assign n34914 =  ( n3051 ) ? ( n34913 ) : ( VREG_10_1 ) ;
assign n34915 =  ( n3040 ) ? ( n34907 ) : ( n34914 ) ;
assign n34916 =  ( n192 ) ? ( VREG_10_1 ) : ( VREG_10_1 ) ;
assign n34917 =  ( n157 ) ? ( n34915 ) : ( n34916 ) ;
assign n34918 =  ( n6 ) ? ( n34902 ) : ( n34917 ) ;
assign n34919 =  ( n219 ) ? ( n34918 ) : ( VREG_10_1 ) ;
assign n34920 =  ( n148 ) ? ( n6232 ) : ( VREG_10_10 ) ;
assign n34921 =  ( n146 ) ? ( n6231 ) : ( n34920 ) ;
assign n34922 =  ( n144 ) ? ( n6230 ) : ( n34921 ) ;
assign n34923 =  ( n142 ) ? ( n6229 ) : ( n34922 ) ;
assign n34924 =  ( n10 ) ? ( n6228 ) : ( n34923 ) ;
assign n34925 =  ( n148 ) ? ( n7266 ) : ( VREG_10_10 ) ;
assign n34926 =  ( n146 ) ? ( n7265 ) : ( n34925 ) ;
assign n34927 =  ( n144 ) ? ( n7264 ) : ( n34926 ) ;
assign n34928 =  ( n142 ) ? ( n7263 ) : ( n34927 ) ;
assign n34929 =  ( n10 ) ? ( n7262 ) : ( n34928 ) ;
assign n34930 =  ( n7273 ) ? ( VREG_10_10 ) : ( n34924 ) ;
assign n34931 =  ( n7273 ) ? ( VREG_10_10 ) : ( n34929 ) ;
assign n34932 =  ( n3034 ) ? ( n34931 ) : ( VREG_10_10 ) ;
assign n34933 =  ( n2965 ) ? ( n34930 ) : ( n34932 ) ;
assign n34934 =  ( n1930 ) ? ( n34929 ) : ( n34933 ) ;
assign n34935 =  ( n879 ) ? ( n34924 ) : ( n34934 ) ;
assign n34936 =  ( n172 ) ? ( n7284 ) : ( VREG_10_10 ) ;
assign n34937 =  ( n170 ) ? ( n7283 ) : ( n34936 ) ;
assign n34938 =  ( n168 ) ? ( n7282 ) : ( n34937 ) ;
assign n34939 =  ( n166 ) ? ( n7281 ) : ( n34938 ) ;
assign n34940 =  ( n162 ) ? ( n7280 ) : ( n34939 ) ;
assign n34941 =  ( n172 ) ? ( n7294 ) : ( VREG_10_10 ) ;
assign n34942 =  ( n170 ) ? ( n7293 ) : ( n34941 ) ;
assign n34943 =  ( n168 ) ? ( n7292 ) : ( n34942 ) ;
assign n34944 =  ( n166 ) ? ( n7291 ) : ( n34943 ) ;
assign n34945 =  ( n162 ) ? ( n7290 ) : ( n34944 ) ;
assign n34946 =  ( n7273 ) ? ( VREG_10_10 ) : ( n34945 ) ;
assign n34947 =  ( n3051 ) ? ( n34946 ) : ( VREG_10_10 ) ;
assign n34948 =  ( n3040 ) ? ( n34940 ) : ( n34947 ) ;
assign n34949 =  ( n192 ) ? ( VREG_10_10 ) : ( VREG_10_10 ) ;
assign n34950 =  ( n157 ) ? ( n34948 ) : ( n34949 ) ;
assign n34951 =  ( n6 ) ? ( n34935 ) : ( n34950 ) ;
assign n34952 =  ( n219 ) ? ( n34951 ) : ( VREG_10_10 ) ;
assign n34953 =  ( n148 ) ? ( n8351 ) : ( VREG_10_11 ) ;
assign n34954 =  ( n146 ) ? ( n8350 ) : ( n34953 ) ;
assign n34955 =  ( n144 ) ? ( n8349 ) : ( n34954 ) ;
assign n34956 =  ( n142 ) ? ( n8348 ) : ( n34955 ) ;
assign n34957 =  ( n10 ) ? ( n8347 ) : ( n34956 ) ;
assign n34958 =  ( n148 ) ? ( n9385 ) : ( VREG_10_11 ) ;
assign n34959 =  ( n146 ) ? ( n9384 ) : ( n34958 ) ;
assign n34960 =  ( n144 ) ? ( n9383 ) : ( n34959 ) ;
assign n34961 =  ( n142 ) ? ( n9382 ) : ( n34960 ) ;
assign n34962 =  ( n10 ) ? ( n9381 ) : ( n34961 ) ;
assign n34963 =  ( n9392 ) ? ( VREG_10_11 ) : ( n34957 ) ;
assign n34964 =  ( n9392 ) ? ( VREG_10_11 ) : ( n34962 ) ;
assign n34965 =  ( n3034 ) ? ( n34964 ) : ( VREG_10_11 ) ;
assign n34966 =  ( n2965 ) ? ( n34963 ) : ( n34965 ) ;
assign n34967 =  ( n1930 ) ? ( n34962 ) : ( n34966 ) ;
assign n34968 =  ( n879 ) ? ( n34957 ) : ( n34967 ) ;
assign n34969 =  ( n172 ) ? ( n9403 ) : ( VREG_10_11 ) ;
assign n34970 =  ( n170 ) ? ( n9402 ) : ( n34969 ) ;
assign n34971 =  ( n168 ) ? ( n9401 ) : ( n34970 ) ;
assign n34972 =  ( n166 ) ? ( n9400 ) : ( n34971 ) ;
assign n34973 =  ( n162 ) ? ( n9399 ) : ( n34972 ) ;
assign n34974 =  ( n172 ) ? ( n9413 ) : ( VREG_10_11 ) ;
assign n34975 =  ( n170 ) ? ( n9412 ) : ( n34974 ) ;
assign n34976 =  ( n168 ) ? ( n9411 ) : ( n34975 ) ;
assign n34977 =  ( n166 ) ? ( n9410 ) : ( n34976 ) ;
assign n34978 =  ( n162 ) ? ( n9409 ) : ( n34977 ) ;
assign n34979 =  ( n9392 ) ? ( VREG_10_11 ) : ( n34978 ) ;
assign n34980 =  ( n3051 ) ? ( n34979 ) : ( VREG_10_11 ) ;
assign n34981 =  ( n3040 ) ? ( n34973 ) : ( n34980 ) ;
assign n34982 =  ( n192 ) ? ( VREG_10_11 ) : ( VREG_10_11 ) ;
assign n34983 =  ( n157 ) ? ( n34981 ) : ( n34982 ) ;
assign n34984 =  ( n6 ) ? ( n34968 ) : ( n34983 ) ;
assign n34985 =  ( n219 ) ? ( n34984 ) : ( VREG_10_11 ) ;
assign n34986 =  ( n148 ) ? ( n10470 ) : ( VREG_10_12 ) ;
assign n34987 =  ( n146 ) ? ( n10469 ) : ( n34986 ) ;
assign n34988 =  ( n144 ) ? ( n10468 ) : ( n34987 ) ;
assign n34989 =  ( n142 ) ? ( n10467 ) : ( n34988 ) ;
assign n34990 =  ( n10 ) ? ( n10466 ) : ( n34989 ) ;
assign n34991 =  ( n148 ) ? ( n11504 ) : ( VREG_10_12 ) ;
assign n34992 =  ( n146 ) ? ( n11503 ) : ( n34991 ) ;
assign n34993 =  ( n144 ) ? ( n11502 ) : ( n34992 ) ;
assign n34994 =  ( n142 ) ? ( n11501 ) : ( n34993 ) ;
assign n34995 =  ( n10 ) ? ( n11500 ) : ( n34994 ) ;
assign n34996 =  ( n11511 ) ? ( VREG_10_12 ) : ( n34990 ) ;
assign n34997 =  ( n11511 ) ? ( VREG_10_12 ) : ( n34995 ) ;
assign n34998 =  ( n3034 ) ? ( n34997 ) : ( VREG_10_12 ) ;
assign n34999 =  ( n2965 ) ? ( n34996 ) : ( n34998 ) ;
assign n35000 =  ( n1930 ) ? ( n34995 ) : ( n34999 ) ;
assign n35001 =  ( n879 ) ? ( n34990 ) : ( n35000 ) ;
assign n35002 =  ( n172 ) ? ( n11522 ) : ( VREG_10_12 ) ;
assign n35003 =  ( n170 ) ? ( n11521 ) : ( n35002 ) ;
assign n35004 =  ( n168 ) ? ( n11520 ) : ( n35003 ) ;
assign n35005 =  ( n166 ) ? ( n11519 ) : ( n35004 ) ;
assign n35006 =  ( n162 ) ? ( n11518 ) : ( n35005 ) ;
assign n35007 =  ( n172 ) ? ( n11532 ) : ( VREG_10_12 ) ;
assign n35008 =  ( n170 ) ? ( n11531 ) : ( n35007 ) ;
assign n35009 =  ( n168 ) ? ( n11530 ) : ( n35008 ) ;
assign n35010 =  ( n166 ) ? ( n11529 ) : ( n35009 ) ;
assign n35011 =  ( n162 ) ? ( n11528 ) : ( n35010 ) ;
assign n35012 =  ( n11511 ) ? ( VREG_10_12 ) : ( n35011 ) ;
assign n35013 =  ( n3051 ) ? ( n35012 ) : ( VREG_10_12 ) ;
assign n35014 =  ( n3040 ) ? ( n35006 ) : ( n35013 ) ;
assign n35015 =  ( n192 ) ? ( VREG_10_12 ) : ( VREG_10_12 ) ;
assign n35016 =  ( n157 ) ? ( n35014 ) : ( n35015 ) ;
assign n35017 =  ( n6 ) ? ( n35001 ) : ( n35016 ) ;
assign n35018 =  ( n219 ) ? ( n35017 ) : ( VREG_10_12 ) ;
assign n35019 =  ( n148 ) ? ( n12589 ) : ( VREG_10_13 ) ;
assign n35020 =  ( n146 ) ? ( n12588 ) : ( n35019 ) ;
assign n35021 =  ( n144 ) ? ( n12587 ) : ( n35020 ) ;
assign n35022 =  ( n142 ) ? ( n12586 ) : ( n35021 ) ;
assign n35023 =  ( n10 ) ? ( n12585 ) : ( n35022 ) ;
assign n35024 =  ( n148 ) ? ( n13623 ) : ( VREG_10_13 ) ;
assign n35025 =  ( n146 ) ? ( n13622 ) : ( n35024 ) ;
assign n35026 =  ( n144 ) ? ( n13621 ) : ( n35025 ) ;
assign n35027 =  ( n142 ) ? ( n13620 ) : ( n35026 ) ;
assign n35028 =  ( n10 ) ? ( n13619 ) : ( n35027 ) ;
assign n35029 =  ( n13630 ) ? ( VREG_10_13 ) : ( n35023 ) ;
assign n35030 =  ( n13630 ) ? ( VREG_10_13 ) : ( n35028 ) ;
assign n35031 =  ( n3034 ) ? ( n35030 ) : ( VREG_10_13 ) ;
assign n35032 =  ( n2965 ) ? ( n35029 ) : ( n35031 ) ;
assign n35033 =  ( n1930 ) ? ( n35028 ) : ( n35032 ) ;
assign n35034 =  ( n879 ) ? ( n35023 ) : ( n35033 ) ;
assign n35035 =  ( n172 ) ? ( n13641 ) : ( VREG_10_13 ) ;
assign n35036 =  ( n170 ) ? ( n13640 ) : ( n35035 ) ;
assign n35037 =  ( n168 ) ? ( n13639 ) : ( n35036 ) ;
assign n35038 =  ( n166 ) ? ( n13638 ) : ( n35037 ) ;
assign n35039 =  ( n162 ) ? ( n13637 ) : ( n35038 ) ;
assign n35040 =  ( n172 ) ? ( n13651 ) : ( VREG_10_13 ) ;
assign n35041 =  ( n170 ) ? ( n13650 ) : ( n35040 ) ;
assign n35042 =  ( n168 ) ? ( n13649 ) : ( n35041 ) ;
assign n35043 =  ( n166 ) ? ( n13648 ) : ( n35042 ) ;
assign n35044 =  ( n162 ) ? ( n13647 ) : ( n35043 ) ;
assign n35045 =  ( n13630 ) ? ( VREG_10_13 ) : ( n35044 ) ;
assign n35046 =  ( n3051 ) ? ( n35045 ) : ( VREG_10_13 ) ;
assign n35047 =  ( n3040 ) ? ( n35039 ) : ( n35046 ) ;
assign n35048 =  ( n192 ) ? ( VREG_10_13 ) : ( VREG_10_13 ) ;
assign n35049 =  ( n157 ) ? ( n35047 ) : ( n35048 ) ;
assign n35050 =  ( n6 ) ? ( n35034 ) : ( n35049 ) ;
assign n35051 =  ( n219 ) ? ( n35050 ) : ( VREG_10_13 ) ;
assign n35052 =  ( n148 ) ? ( n14708 ) : ( VREG_10_14 ) ;
assign n35053 =  ( n146 ) ? ( n14707 ) : ( n35052 ) ;
assign n35054 =  ( n144 ) ? ( n14706 ) : ( n35053 ) ;
assign n35055 =  ( n142 ) ? ( n14705 ) : ( n35054 ) ;
assign n35056 =  ( n10 ) ? ( n14704 ) : ( n35055 ) ;
assign n35057 =  ( n148 ) ? ( n15742 ) : ( VREG_10_14 ) ;
assign n35058 =  ( n146 ) ? ( n15741 ) : ( n35057 ) ;
assign n35059 =  ( n144 ) ? ( n15740 ) : ( n35058 ) ;
assign n35060 =  ( n142 ) ? ( n15739 ) : ( n35059 ) ;
assign n35061 =  ( n10 ) ? ( n15738 ) : ( n35060 ) ;
assign n35062 =  ( n15749 ) ? ( VREG_10_14 ) : ( n35056 ) ;
assign n35063 =  ( n15749 ) ? ( VREG_10_14 ) : ( n35061 ) ;
assign n35064 =  ( n3034 ) ? ( n35063 ) : ( VREG_10_14 ) ;
assign n35065 =  ( n2965 ) ? ( n35062 ) : ( n35064 ) ;
assign n35066 =  ( n1930 ) ? ( n35061 ) : ( n35065 ) ;
assign n35067 =  ( n879 ) ? ( n35056 ) : ( n35066 ) ;
assign n35068 =  ( n172 ) ? ( n15760 ) : ( VREG_10_14 ) ;
assign n35069 =  ( n170 ) ? ( n15759 ) : ( n35068 ) ;
assign n35070 =  ( n168 ) ? ( n15758 ) : ( n35069 ) ;
assign n35071 =  ( n166 ) ? ( n15757 ) : ( n35070 ) ;
assign n35072 =  ( n162 ) ? ( n15756 ) : ( n35071 ) ;
assign n35073 =  ( n172 ) ? ( n15770 ) : ( VREG_10_14 ) ;
assign n35074 =  ( n170 ) ? ( n15769 ) : ( n35073 ) ;
assign n35075 =  ( n168 ) ? ( n15768 ) : ( n35074 ) ;
assign n35076 =  ( n166 ) ? ( n15767 ) : ( n35075 ) ;
assign n35077 =  ( n162 ) ? ( n15766 ) : ( n35076 ) ;
assign n35078 =  ( n15749 ) ? ( VREG_10_14 ) : ( n35077 ) ;
assign n35079 =  ( n3051 ) ? ( n35078 ) : ( VREG_10_14 ) ;
assign n35080 =  ( n3040 ) ? ( n35072 ) : ( n35079 ) ;
assign n35081 =  ( n192 ) ? ( VREG_10_14 ) : ( VREG_10_14 ) ;
assign n35082 =  ( n157 ) ? ( n35080 ) : ( n35081 ) ;
assign n35083 =  ( n6 ) ? ( n35067 ) : ( n35082 ) ;
assign n35084 =  ( n219 ) ? ( n35083 ) : ( VREG_10_14 ) ;
assign n35085 =  ( n148 ) ? ( n16827 ) : ( VREG_10_15 ) ;
assign n35086 =  ( n146 ) ? ( n16826 ) : ( n35085 ) ;
assign n35087 =  ( n144 ) ? ( n16825 ) : ( n35086 ) ;
assign n35088 =  ( n142 ) ? ( n16824 ) : ( n35087 ) ;
assign n35089 =  ( n10 ) ? ( n16823 ) : ( n35088 ) ;
assign n35090 =  ( n148 ) ? ( n17861 ) : ( VREG_10_15 ) ;
assign n35091 =  ( n146 ) ? ( n17860 ) : ( n35090 ) ;
assign n35092 =  ( n144 ) ? ( n17859 ) : ( n35091 ) ;
assign n35093 =  ( n142 ) ? ( n17858 ) : ( n35092 ) ;
assign n35094 =  ( n10 ) ? ( n17857 ) : ( n35093 ) ;
assign n35095 =  ( n17868 ) ? ( VREG_10_15 ) : ( n35089 ) ;
assign n35096 =  ( n17868 ) ? ( VREG_10_15 ) : ( n35094 ) ;
assign n35097 =  ( n3034 ) ? ( n35096 ) : ( VREG_10_15 ) ;
assign n35098 =  ( n2965 ) ? ( n35095 ) : ( n35097 ) ;
assign n35099 =  ( n1930 ) ? ( n35094 ) : ( n35098 ) ;
assign n35100 =  ( n879 ) ? ( n35089 ) : ( n35099 ) ;
assign n35101 =  ( n172 ) ? ( n17879 ) : ( VREG_10_15 ) ;
assign n35102 =  ( n170 ) ? ( n17878 ) : ( n35101 ) ;
assign n35103 =  ( n168 ) ? ( n17877 ) : ( n35102 ) ;
assign n35104 =  ( n166 ) ? ( n17876 ) : ( n35103 ) ;
assign n35105 =  ( n162 ) ? ( n17875 ) : ( n35104 ) ;
assign n35106 =  ( n172 ) ? ( n17889 ) : ( VREG_10_15 ) ;
assign n35107 =  ( n170 ) ? ( n17888 ) : ( n35106 ) ;
assign n35108 =  ( n168 ) ? ( n17887 ) : ( n35107 ) ;
assign n35109 =  ( n166 ) ? ( n17886 ) : ( n35108 ) ;
assign n35110 =  ( n162 ) ? ( n17885 ) : ( n35109 ) ;
assign n35111 =  ( n17868 ) ? ( VREG_10_15 ) : ( n35110 ) ;
assign n35112 =  ( n3051 ) ? ( n35111 ) : ( VREG_10_15 ) ;
assign n35113 =  ( n3040 ) ? ( n35105 ) : ( n35112 ) ;
assign n35114 =  ( n192 ) ? ( VREG_10_15 ) : ( VREG_10_15 ) ;
assign n35115 =  ( n157 ) ? ( n35113 ) : ( n35114 ) ;
assign n35116 =  ( n6 ) ? ( n35100 ) : ( n35115 ) ;
assign n35117 =  ( n219 ) ? ( n35116 ) : ( VREG_10_15 ) ;
assign n35118 =  ( n148 ) ? ( n18946 ) : ( VREG_10_2 ) ;
assign n35119 =  ( n146 ) ? ( n18945 ) : ( n35118 ) ;
assign n35120 =  ( n144 ) ? ( n18944 ) : ( n35119 ) ;
assign n35121 =  ( n142 ) ? ( n18943 ) : ( n35120 ) ;
assign n35122 =  ( n10 ) ? ( n18942 ) : ( n35121 ) ;
assign n35123 =  ( n148 ) ? ( n19980 ) : ( VREG_10_2 ) ;
assign n35124 =  ( n146 ) ? ( n19979 ) : ( n35123 ) ;
assign n35125 =  ( n144 ) ? ( n19978 ) : ( n35124 ) ;
assign n35126 =  ( n142 ) ? ( n19977 ) : ( n35125 ) ;
assign n35127 =  ( n10 ) ? ( n19976 ) : ( n35126 ) ;
assign n35128 =  ( n19987 ) ? ( VREG_10_2 ) : ( n35122 ) ;
assign n35129 =  ( n19987 ) ? ( VREG_10_2 ) : ( n35127 ) ;
assign n35130 =  ( n3034 ) ? ( n35129 ) : ( VREG_10_2 ) ;
assign n35131 =  ( n2965 ) ? ( n35128 ) : ( n35130 ) ;
assign n35132 =  ( n1930 ) ? ( n35127 ) : ( n35131 ) ;
assign n35133 =  ( n879 ) ? ( n35122 ) : ( n35132 ) ;
assign n35134 =  ( n172 ) ? ( n19998 ) : ( VREG_10_2 ) ;
assign n35135 =  ( n170 ) ? ( n19997 ) : ( n35134 ) ;
assign n35136 =  ( n168 ) ? ( n19996 ) : ( n35135 ) ;
assign n35137 =  ( n166 ) ? ( n19995 ) : ( n35136 ) ;
assign n35138 =  ( n162 ) ? ( n19994 ) : ( n35137 ) ;
assign n35139 =  ( n172 ) ? ( n20008 ) : ( VREG_10_2 ) ;
assign n35140 =  ( n170 ) ? ( n20007 ) : ( n35139 ) ;
assign n35141 =  ( n168 ) ? ( n20006 ) : ( n35140 ) ;
assign n35142 =  ( n166 ) ? ( n20005 ) : ( n35141 ) ;
assign n35143 =  ( n162 ) ? ( n20004 ) : ( n35142 ) ;
assign n35144 =  ( n19987 ) ? ( VREG_10_2 ) : ( n35143 ) ;
assign n35145 =  ( n3051 ) ? ( n35144 ) : ( VREG_10_2 ) ;
assign n35146 =  ( n3040 ) ? ( n35138 ) : ( n35145 ) ;
assign n35147 =  ( n192 ) ? ( VREG_10_2 ) : ( VREG_10_2 ) ;
assign n35148 =  ( n157 ) ? ( n35146 ) : ( n35147 ) ;
assign n35149 =  ( n6 ) ? ( n35133 ) : ( n35148 ) ;
assign n35150 =  ( n219 ) ? ( n35149 ) : ( VREG_10_2 ) ;
assign n35151 =  ( n148 ) ? ( n21065 ) : ( VREG_10_3 ) ;
assign n35152 =  ( n146 ) ? ( n21064 ) : ( n35151 ) ;
assign n35153 =  ( n144 ) ? ( n21063 ) : ( n35152 ) ;
assign n35154 =  ( n142 ) ? ( n21062 ) : ( n35153 ) ;
assign n35155 =  ( n10 ) ? ( n21061 ) : ( n35154 ) ;
assign n35156 =  ( n148 ) ? ( n22099 ) : ( VREG_10_3 ) ;
assign n35157 =  ( n146 ) ? ( n22098 ) : ( n35156 ) ;
assign n35158 =  ( n144 ) ? ( n22097 ) : ( n35157 ) ;
assign n35159 =  ( n142 ) ? ( n22096 ) : ( n35158 ) ;
assign n35160 =  ( n10 ) ? ( n22095 ) : ( n35159 ) ;
assign n35161 =  ( n22106 ) ? ( VREG_10_3 ) : ( n35155 ) ;
assign n35162 =  ( n22106 ) ? ( VREG_10_3 ) : ( n35160 ) ;
assign n35163 =  ( n3034 ) ? ( n35162 ) : ( VREG_10_3 ) ;
assign n35164 =  ( n2965 ) ? ( n35161 ) : ( n35163 ) ;
assign n35165 =  ( n1930 ) ? ( n35160 ) : ( n35164 ) ;
assign n35166 =  ( n879 ) ? ( n35155 ) : ( n35165 ) ;
assign n35167 =  ( n172 ) ? ( n22117 ) : ( VREG_10_3 ) ;
assign n35168 =  ( n170 ) ? ( n22116 ) : ( n35167 ) ;
assign n35169 =  ( n168 ) ? ( n22115 ) : ( n35168 ) ;
assign n35170 =  ( n166 ) ? ( n22114 ) : ( n35169 ) ;
assign n35171 =  ( n162 ) ? ( n22113 ) : ( n35170 ) ;
assign n35172 =  ( n172 ) ? ( n22127 ) : ( VREG_10_3 ) ;
assign n35173 =  ( n170 ) ? ( n22126 ) : ( n35172 ) ;
assign n35174 =  ( n168 ) ? ( n22125 ) : ( n35173 ) ;
assign n35175 =  ( n166 ) ? ( n22124 ) : ( n35174 ) ;
assign n35176 =  ( n162 ) ? ( n22123 ) : ( n35175 ) ;
assign n35177 =  ( n22106 ) ? ( VREG_10_3 ) : ( n35176 ) ;
assign n35178 =  ( n3051 ) ? ( n35177 ) : ( VREG_10_3 ) ;
assign n35179 =  ( n3040 ) ? ( n35171 ) : ( n35178 ) ;
assign n35180 =  ( n192 ) ? ( VREG_10_3 ) : ( VREG_10_3 ) ;
assign n35181 =  ( n157 ) ? ( n35179 ) : ( n35180 ) ;
assign n35182 =  ( n6 ) ? ( n35166 ) : ( n35181 ) ;
assign n35183 =  ( n219 ) ? ( n35182 ) : ( VREG_10_3 ) ;
assign n35184 =  ( n148 ) ? ( n23184 ) : ( VREG_10_4 ) ;
assign n35185 =  ( n146 ) ? ( n23183 ) : ( n35184 ) ;
assign n35186 =  ( n144 ) ? ( n23182 ) : ( n35185 ) ;
assign n35187 =  ( n142 ) ? ( n23181 ) : ( n35186 ) ;
assign n35188 =  ( n10 ) ? ( n23180 ) : ( n35187 ) ;
assign n35189 =  ( n148 ) ? ( n24218 ) : ( VREG_10_4 ) ;
assign n35190 =  ( n146 ) ? ( n24217 ) : ( n35189 ) ;
assign n35191 =  ( n144 ) ? ( n24216 ) : ( n35190 ) ;
assign n35192 =  ( n142 ) ? ( n24215 ) : ( n35191 ) ;
assign n35193 =  ( n10 ) ? ( n24214 ) : ( n35192 ) ;
assign n35194 =  ( n24225 ) ? ( VREG_10_4 ) : ( n35188 ) ;
assign n35195 =  ( n24225 ) ? ( VREG_10_4 ) : ( n35193 ) ;
assign n35196 =  ( n3034 ) ? ( n35195 ) : ( VREG_10_4 ) ;
assign n35197 =  ( n2965 ) ? ( n35194 ) : ( n35196 ) ;
assign n35198 =  ( n1930 ) ? ( n35193 ) : ( n35197 ) ;
assign n35199 =  ( n879 ) ? ( n35188 ) : ( n35198 ) ;
assign n35200 =  ( n172 ) ? ( n24236 ) : ( VREG_10_4 ) ;
assign n35201 =  ( n170 ) ? ( n24235 ) : ( n35200 ) ;
assign n35202 =  ( n168 ) ? ( n24234 ) : ( n35201 ) ;
assign n35203 =  ( n166 ) ? ( n24233 ) : ( n35202 ) ;
assign n35204 =  ( n162 ) ? ( n24232 ) : ( n35203 ) ;
assign n35205 =  ( n172 ) ? ( n24246 ) : ( VREG_10_4 ) ;
assign n35206 =  ( n170 ) ? ( n24245 ) : ( n35205 ) ;
assign n35207 =  ( n168 ) ? ( n24244 ) : ( n35206 ) ;
assign n35208 =  ( n166 ) ? ( n24243 ) : ( n35207 ) ;
assign n35209 =  ( n162 ) ? ( n24242 ) : ( n35208 ) ;
assign n35210 =  ( n24225 ) ? ( VREG_10_4 ) : ( n35209 ) ;
assign n35211 =  ( n3051 ) ? ( n35210 ) : ( VREG_10_4 ) ;
assign n35212 =  ( n3040 ) ? ( n35204 ) : ( n35211 ) ;
assign n35213 =  ( n192 ) ? ( VREG_10_4 ) : ( VREG_10_4 ) ;
assign n35214 =  ( n157 ) ? ( n35212 ) : ( n35213 ) ;
assign n35215 =  ( n6 ) ? ( n35199 ) : ( n35214 ) ;
assign n35216 =  ( n219 ) ? ( n35215 ) : ( VREG_10_4 ) ;
assign n35217 =  ( n148 ) ? ( n25303 ) : ( VREG_10_5 ) ;
assign n35218 =  ( n146 ) ? ( n25302 ) : ( n35217 ) ;
assign n35219 =  ( n144 ) ? ( n25301 ) : ( n35218 ) ;
assign n35220 =  ( n142 ) ? ( n25300 ) : ( n35219 ) ;
assign n35221 =  ( n10 ) ? ( n25299 ) : ( n35220 ) ;
assign n35222 =  ( n148 ) ? ( n26337 ) : ( VREG_10_5 ) ;
assign n35223 =  ( n146 ) ? ( n26336 ) : ( n35222 ) ;
assign n35224 =  ( n144 ) ? ( n26335 ) : ( n35223 ) ;
assign n35225 =  ( n142 ) ? ( n26334 ) : ( n35224 ) ;
assign n35226 =  ( n10 ) ? ( n26333 ) : ( n35225 ) ;
assign n35227 =  ( n26344 ) ? ( VREG_10_5 ) : ( n35221 ) ;
assign n35228 =  ( n26344 ) ? ( VREG_10_5 ) : ( n35226 ) ;
assign n35229 =  ( n3034 ) ? ( n35228 ) : ( VREG_10_5 ) ;
assign n35230 =  ( n2965 ) ? ( n35227 ) : ( n35229 ) ;
assign n35231 =  ( n1930 ) ? ( n35226 ) : ( n35230 ) ;
assign n35232 =  ( n879 ) ? ( n35221 ) : ( n35231 ) ;
assign n35233 =  ( n172 ) ? ( n26355 ) : ( VREG_10_5 ) ;
assign n35234 =  ( n170 ) ? ( n26354 ) : ( n35233 ) ;
assign n35235 =  ( n168 ) ? ( n26353 ) : ( n35234 ) ;
assign n35236 =  ( n166 ) ? ( n26352 ) : ( n35235 ) ;
assign n35237 =  ( n162 ) ? ( n26351 ) : ( n35236 ) ;
assign n35238 =  ( n172 ) ? ( n26365 ) : ( VREG_10_5 ) ;
assign n35239 =  ( n170 ) ? ( n26364 ) : ( n35238 ) ;
assign n35240 =  ( n168 ) ? ( n26363 ) : ( n35239 ) ;
assign n35241 =  ( n166 ) ? ( n26362 ) : ( n35240 ) ;
assign n35242 =  ( n162 ) ? ( n26361 ) : ( n35241 ) ;
assign n35243 =  ( n26344 ) ? ( VREG_10_5 ) : ( n35242 ) ;
assign n35244 =  ( n3051 ) ? ( n35243 ) : ( VREG_10_5 ) ;
assign n35245 =  ( n3040 ) ? ( n35237 ) : ( n35244 ) ;
assign n35246 =  ( n192 ) ? ( VREG_10_5 ) : ( VREG_10_5 ) ;
assign n35247 =  ( n157 ) ? ( n35245 ) : ( n35246 ) ;
assign n35248 =  ( n6 ) ? ( n35232 ) : ( n35247 ) ;
assign n35249 =  ( n219 ) ? ( n35248 ) : ( VREG_10_5 ) ;
assign n35250 =  ( n148 ) ? ( n27422 ) : ( VREG_10_6 ) ;
assign n35251 =  ( n146 ) ? ( n27421 ) : ( n35250 ) ;
assign n35252 =  ( n144 ) ? ( n27420 ) : ( n35251 ) ;
assign n35253 =  ( n142 ) ? ( n27419 ) : ( n35252 ) ;
assign n35254 =  ( n10 ) ? ( n27418 ) : ( n35253 ) ;
assign n35255 =  ( n148 ) ? ( n28456 ) : ( VREG_10_6 ) ;
assign n35256 =  ( n146 ) ? ( n28455 ) : ( n35255 ) ;
assign n35257 =  ( n144 ) ? ( n28454 ) : ( n35256 ) ;
assign n35258 =  ( n142 ) ? ( n28453 ) : ( n35257 ) ;
assign n35259 =  ( n10 ) ? ( n28452 ) : ( n35258 ) ;
assign n35260 =  ( n28463 ) ? ( VREG_10_6 ) : ( n35254 ) ;
assign n35261 =  ( n28463 ) ? ( VREG_10_6 ) : ( n35259 ) ;
assign n35262 =  ( n3034 ) ? ( n35261 ) : ( VREG_10_6 ) ;
assign n35263 =  ( n2965 ) ? ( n35260 ) : ( n35262 ) ;
assign n35264 =  ( n1930 ) ? ( n35259 ) : ( n35263 ) ;
assign n35265 =  ( n879 ) ? ( n35254 ) : ( n35264 ) ;
assign n35266 =  ( n172 ) ? ( n28474 ) : ( VREG_10_6 ) ;
assign n35267 =  ( n170 ) ? ( n28473 ) : ( n35266 ) ;
assign n35268 =  ( n168 ) ? ( n28472 ) : ( n35267 ) ;
assign n35269 =  ( n166 ) ? ( n28471 ) : ( n35268 ) ;
assign n35270 =  ( n162 ) ? ( n28470 ) : ( n35269 ) ;
assign n35271 =  ( n172 ) ? ( n28484 ) : ( VREG_10_6 ) ;
assign n35272 =  ( n170 ) ? ( n28483 ) : ( n35271 ) ;
assign n35273 =  ( n168 ) ? ( n28482 ) : ( n35272 ) ;
assign n35274 =  ( n166 ) ? ( n28481 ) : ( n35273 ) ;
assign n35275 =  ( n162 ) ? ( n28480 ) : ( n35274 ) ;
assign n35276 =  ( n28463 ) ? ( VREG_10_6 ) : ( n35275 ) ;
assign n35277 =  ( n3051 ) ? ( n35276 ) : ( VREG_10_6 ) ;
assign n35278 =  ( n3040 ) ? ( n35270 ) : ( n35277 ) ;
assign n35279 =  ( n192 ) ? ( VREG_10_6 ) : ( VREG_10_6 ) ;
assign n35280 =  ( n157 ) ? ( n35278 ) : ( n35279 ) ;
assign n35281 =  ( n6 ) ? ( n35265 ) : ( n35280 ) ;
assign n35282 =  ( n219 ) ? ( n35281 ) : ( VREG_10_6 ) ;
assign n35283 =  ( n148 ) ? ( n29541 ) : ( VREG_10_7 ) ;
assign n35284 =  ( n146 ) ? ( n29540 ) : ( n35283 ) ;
assign n35285 =  ( n144 ) ? ( n29539 ) : ( n35284 ) ;
assign n35286 =  ( n142 ) ? ( n29538 ) : ( n35285 ) ;
assign n35287 =  ( n10 ) ? ( n29537 ) : ( n35286 ) ;
assign n35288 =  ( n148 ) ? ( n30575 ) : ( VREG_10_7 ) ;
assign n35289 =  ( n146 ) ? ( n30574 ) : ( n35288 ) ;
assign n35290 =  ( n144 ) ? ( n30573 ) : ( n35289 ) ;
assign n35291 =  ( n142 ) ? ( n30572 ) : ( n35290 ) ;
assign n35292 =  ( n10 ) ? ( n30571 ) : ( n35291 ) ;
assign n35293 =  ( n30582 ) ? ( VREG_10_7 ) : ( n35287 ) ;
assign n35294 =  ( n30582 ) ? ( VREG_10_7 ) : ( n35292 ) ;
assign n35295 =  ( n3034 ) ? ( n35294 ) : ( VREG_10_7 ) ;
assign n35296 =  ( n2965 ) ? ( n35293 ) : ( n35295 ) ;
assign n35297 =  ( n1930 ) ? ( n35292 ) : ( n35296 ) ;
assign n35298 =  ( n879 ) ? ( n35287 ) : ( n35297 ) ;
assign n35299 =  ( n172 ) ? ( n30593 ) : ( VREG_10_7 ) ;
assign n35300 =  ( n170 ) ? ( n30592 ) : ( n35299 ) ;
assign n35301 =  ( n168 ) ? ( n30591 ) : ( n35300 ) ;
assign n35302 =  ( n166 ) ? ( n30590 ) : ( n35301 ) ;
assign n35303 =  ( n162 ) ? ( n30589 ) : ( n35302 ) ;
assign n35304 =  ( n172 ) ? ( n30603 ) : ( VREG_10_7 ) ;
assign n35305 =  ( n170 ) ? ( n30602 ) : ( n35304 ) ;
assign n35306 =  ( n168 ) ? ( n30601 ) : ( n35305 ) ;
assign n35307 =  ( n166 ) ? ( n30600 ) : ( n35306 ) ;
assign n35308 =  ( n162 ) ? ( n30599 ) : ( n35307 ) ;
assign n35309 =  ( n30582 ) ? ( VREG_10_7 ) : ( n35308 ) ;
assign n35310 =  ( n3051 ) ? ( n35309 ) : ( VREG_10_7 ) ;
assign n35311 =  ( n3040 ) ? ( n35303 ) : ( n35310 ) ;
assign n35312 =  ( n192 ) ? ( VREG_10_7 ) : ( VREG_10_7 ) ;
assign n35313 =  ( n157 ) ? ( n35311 ) : ( n35312 ) ;
assign n35314 =  ( n6 ) ? ( n35298 ) : ( n35313 ) ;
assign n35315 =  ( n219 ) ? ( n35314 ) : ( VREG_10_7 ) ;
assign n35316 =  ( n148 ) ? ( n31660 ) : ( VREG_10_8 ) ;
assign n35317 =  ( n146 ) ? ( n31659 ) : ( n35316 ) ;
assign n35318 =  ( n144 ) ? ( n31658 ) : ( n35317 ) ;
assign n35319 =  ( n142 ) ? ( n31657 ) : ( n35318 ) ;
assign n35320 =  ( n10 ) ? ( n31656 ) : ( n35319 ) ;
assign n35321 =  ( n148 ) ? ( n32694 ) : ( VREG_10_8 ) ;
assign n35322 =  ( n146 ) ? ( n32693 ) : ( n35321 ) ;
assign n35323 =  ( n144 ) ? ( n32692 ) : ( n35322 ) ;
assign n35324 =  ( n142 ) ? ( n32691 ) : ( n35323 ) ;
assign n35325 =  ( n10 ) ? ( n32690 ) : ( n35324 ) ;
assign n35326 =  ( n32701 ) ? ( VREG_10_8 ) : ( n35320 ) ;
assign n35327 =  ( n32701 ) ? ( VREG_10_8 ) : ( n35325 ) ;
assign n35328 =  ( n3034 ) ? ( n35327 ) : ( VREG_10_8 ) ;
assign n35329 =  ( n2965 ) ? ( n35326 ) : ( n35328 ) ;
assign n35330 =  ( n1930 ) ? ( n35325 ) : ( n35329 ) ;
assign n35331 =  ( n879 ) ? ( n35320 ) : ( n35330 ) ;
assign n35332 =  ( n172 ) ? ( n32712 ) : ( VREG_10_8 ) ;
assign n35333 =  ( n170 ) ? ( n32711 ) : ( n35332 ) ;
assign n35334 =  ( n168 ) ? ( n32710 ) : ( n35333 ) ;
assign n35335 =  ( n166 ) ? ( n32709 ) : ( n35334 ) ;
assign n35336 =  ( n162 ) ? ( n32708 ) : ( n35335 ) ;
assign n35337 =  ( n172 ) ? ( n32722 ) : ( VREG_10_8 ) ;
assign n35338 =  ( n170 ) ? ( n32721 ) : ( n35337 ) ;
assign n35339 =  ( n168 ) ? ( n32720 ) : ( n35338 ) ;
assign n35340 =  ( n166 ) ? ( n32719 ) : ( n35339 ) ;
assign n35341 =  ( n162 ) ? ( n32718 ) : ( n35340 ) ;
assign n35342 =  ( n32701 ) ? ( VREG_10_8 ) : ( n35341 ) ;
assign n35343 =  ( n3051 ) ? ( n35342 ) : ( VREG_10_8 ) ;
assign n35344 =  ( n3040 ) ? ( n35336 ) : ( n35343 ) ;
assign n35345 =  ( n192 ) ? ( VREG_10_8 ) : ( VREG_10_8 ) ;
assign n35346 =  ( n157 ) ? ( n35344 ) : ( n35345 ) ;
assign n35347 =  ( n6 ) ? ( n35331 ) : ( n35346 ) ;
assign n35348 =  ( n219 ) ? ( n35347 ) : ( VREG_10_8 ) ;
assign n35349 =  ( n148 ) ? ( n33779 ) : ( VREG_10_9 ) ;
assign n35350 =  ( n146 ) ? ( n33778 ) : ( n35349 ) ;
assign n35351 =  ( n144 ) ? ( n33777 ) : ( n35350 ) ;
assign n35352 =  ( n142 ) ? ( n33776 ) : ( n35351 ) ;
assign n35353 =  ( n10 ) ? ( n33775 ) : ( n35352 ) ;
assign n35354 =  ( n148 ) ? ( n34813 ) : ( VREG_10_9 ) ;
assign n35355 =  ( n146 ) ? ( n34812 ) : ( n35354 ) ;
assign n35356 =  ( n144 ) ? ( n34811 ) : ( n35355 ) ;
assign n35357 =  ( n142 ) ? ( n34810 ) : ( n35356 ) ;
assign n35358 =  ( n10 ) ? ( n34809 ) : ( n35357 ) ;
assign n35359 =  ( n34820 ) ? ( VREG_10_9 ) : ( n35353 ) ;
assign n35360 =  ( n34820 ) ? ( VREG_10_9 ) : ( n35358 ) ;
assign n35361 =  ( n3034 ) ? ( n35360 ) : ( VREG_10_9 ) ;
assign n35362 =  ( n2965 ) ? ( n35359 ) : ( n35361 ) ;
assign n35363 =  ( n1930 ) ? ( n35358 ) : ( n35362 ) ;
assign n35364 =  ( n879 ) ? ( n35353 ) : ( n35363 ) ;
assign n35365 =  ( n172 ) ? ( n34831 ) : ( VREG_10_9 ) ;
assign n35366 =  ( n170 ) ? ( n34830 ) : ( n35365 ) ;
assign n35367 =  ( n168 ) ? ( n34829 ) : ( n35366 ) ;
assign n35368 =  ( n166 ) ? ( n34828 ) : ( n35367 ) ;
assign n35369 =  ( n162 ) ? ( n34827 ) : ( n35368 ) ;
assign n35370 =  ( n172 ) ? ( n34841 ) : ( VREG_10_9 ) ;
assign n35371 =  ( n170 ) ? ( n34840 ) : ( n35370 ) ;
assign n35372 =  ( n168 ) ? ( n34839 ) : ( n35371 ) ;
assign n35373 =  ( n166 ) ? ( n34838 ) : ( n35372 ) ;
assign n35374 =  ( n162 ) ? ( n34837 ) : ( n35373 ) ;
assign n35375 =  ( n34820 ) ? ( VREG_10_9 ) : ( n35374 ) ;
assign n35376 =  ( n3051 ) ? ( n35375 ) : ( VREG_10_9 ) ;
assign n35377 =  ( n3040 ) ? ( n35369 ) : ( n35376 ) ;
assign n35378 =  ( n192 ) ? ( VREG_10_9 ) : ( VREG_10_9 ) ;
assign n35379 =  ( n157 ) ? ( n35377 ) : ( n35378 ) ;
assign n35380 =  ( n6 ) ? ( n35364 ) : ( n35379 ) ;
assign n35381 =  ( n219 ) ? ( n35380 ) : ( VREG_10_9 ) ;
assign n35382 =  ( n148 ) ? ( n1924 ) : ( VREG_11_0 ) ;
assign n35383 =  ( n146 ) ? ( n1923 ) : ( n35382 ) ;
assign n35384 =  ( n144 ) ? ( n1922 ) : ( n35383 ) ;
assign n35385 =  ( n142 ) ? ( n1921 ) : ( n35384 ) ;
assign n35386 =  ( n10 ) ? ( n1920 ) : ( n35385 ) ;
assign n35387 =  ( n148 ) ? ( n2959 ) : ( VREG_11_0 ) ;
assign n35388 =  ( n146 ) ? ( n2958 ) : ( n35387 ) ;
assign n35389 =  ( n144 ) ? ( n2957 ) : ( n35388 ) ;
assign n35390 =  ( n142 ) ? ( n2956 ) : ( n35389 ) ;
assign n35391 =  ( n10 ) ? ( n2955 ) : ( n35390 ) ;
assign n35392 =  ( n3032 ) ? ( VREG_11_0 ) : ( n35386 ) ;
assign n35393 =  ( n3032 ) ? ( VREG_11_0 ) : ( n35391 ) ;
assign n35394 =  ( n3034 ) ? ( n35393 ) : ( VREG_11_0 ) ;
assign n35395 =  ( n2965 ) ? ( n35392 ) : ( n35394 ) ;
assign n35396 =  ( n1930 ) ? ( n35391 ) : ( n35395 ) ;
assign n35397 =  ( n879 ) ? ( n35386 ) : ( n35396 ) ;
assign n35398 =  ( n172 ) ? ( n3045 ) : ( VREG_11_0 ) ;
assign n35399 =  ( n170 ) ? ( n3044 ) : ( n35398 ) ;
assign n35400 =  ( n168 ) ? ( n3043 ) : ( n35399 ) ;
assign n35401 =  ( n166 ) ? ( n3042 ) : ( n35400 ) ;
assign n35402 =  ( n162 ) ? ( n3041 ) : ( n35401 ) ;
assign n35403 =  ( n172 ) ? ( n3056 ) : ( VREG_11_0 ) ;
assign n35404 =  ( n170 ) ? ( n3055 ) : ( n35403 ) ;
assign n35405 =  ( n168 ) ? ( n3054 ) : ( n35404 ) ;
assign n35406 =  ( n166 ) ? ( n3053 ) : ( n35405 ) ;
assign n35407 =  ( n162 ) ? ( n3052 ) : ( n35406 ) ;
assign n35408 =  ( n3032 ) ? ( VREG_11_0 ) : ( n35407 ) ;
assign n35409 =  ( n3051 ) ? ( n35408 ) : ( VREG_11_0 ) ;
assign n35410 =  ( n3040 ) ? ( n35402 ) : ( n35409 ) ;
assign n35411 =  ( n192 ) ? ( VREG_11_0 ) : ( VREG_11_0 ) ;
assign n35412 =  ( n157 ) ? ( n35410 ) : ( n35411 ) ;
assign n35413 =  ( n6 ) ? ( n35397 ) : ( n35412 ) ;
assign n35414 =  ( n241 ) ? ( n35413 ) : ( VREG_11_0 ) ;
assign n35415 =  ( n148 ) ? ( n4113 ) : ( VREG_11_1 ) ;
assign n35416 =  ( n146 ) ? ( n4112 ) : ( n35415 ) ;
assign n35417 =  ( n144 ) ? ( n4111 ) : ( n35416 ) ;
assign n35418 =  ( n142 ) ? ( n4110 ) : ( n35417 ) ;
assign n35419 =  ( n10 ) ? ( n4109 ) : ( n35418 ) ;
assign n35420 =  ( n148 ) ? ( n5147 ) : ( VREG_11_1 ) ;
assign n35421 =  ( n146 ) ? ( n5146 ) : ( n35420 ) ;
assign n35422 =  ( n144 ) ? ( n5145 ) : ( n35421 ) ;
assign n35423 =  ( n142 ) ? ( n5144 ) : ( n35422 ) ;
assign n35424 =  ( n10 ) ? ( n5143 ) : ( n35423 ) ;
assign n35425 =  ( n5154 ) ? ( VREG_11_1 ) : ( n35419 ) ;
assign n35426 =  ( n5154 ) ? ( VREG_11_1 ) : ( n35424 ) ;
assign n35427 =  ( n3034 ) ? ( n35426 ) : ( VREG_11_1 ) ;
assign n35428 =  ( n2965 ) ? ( n35425 ) : ( n35427 ) ;
assign n35429 =  ( n1930 ) ? ( n35424 ) : ( n35428 ) ;
assign n35430 =  ( n879 ) ? ( n35419 ) : ( n35429 ) ;
assign n35431 =  ( n172 ) ? ( n5165 ) : ( VREG_11_1 ) ;
assign n35432 =  ( n170 ) ? ( n5164 ) : ( n35431 ) ;
assign n35433 =  ( n168 ) ? ( n5163 ) : ( n35432 ) ;
assign n35434 =  ( n166 ) ? ( n5162 ) : ( n35433 ) ;
assign n35435 =  ( n162 ) ? ( n5161 ) : ( n35434 ) ;
assign n35436 =  ( n172 ) ? ( n5175 ) : ( VREG_11_1 ) ;
assign n35437 =  ( n170 ) ? ( n5174 ) : ( n35436 ) ;
assign n35438 =  ( n168 ) ? ( n5173 ) : ( n35437 ) ;
assign n35439 =  ( n166 ) ? ( n5172 ) : ( n35438 ) ;
assign n35440 =  ( n162 ) ? ( n5171 ) : ( n35439 ) ;
assign n35441 =  ( n5154 ) ? ( VREG_11_1 ) : ( n35440 ) ;
assign n35442 =  ( n3051 ) ? ( n35441 ) : ( VREG_11_1 ) ;
assign n35443 =  ( n3040 ) ? ( n35435 ) : ( n35442 ) ;
assign n35444 =  ( n192 ) ? ( VREG_11_1 ) : ( VREG_11_1 ) ;
assign n35445 =  ( n157 ) ? ( n35443 ) : ( n35444 ) ;
assign n35446 =  ( n6 ) ? ( n35430 ) : ( n35445 ) ;
assign n35447 =  ( n241 ) ? ( n35446 ) : ( VREG_11_1 ) ;
assign n35448 =  ( n148 ) ? ( n6232 ) : ( VREG_11_10 ) ;
assign n35449 =  ( n146 ) ? ( n6231 ) : ( n35448 ) ;
assign n35450 =  ( n144 ) ? ( n6230 ) : ( n35449 ) ;
assign n35451 =  ( n142 ) ? ( n6229 ) : ( n35450 ) ;
assign n35452 =  ( n10 ) ? ( n6228 ) : ( n35451 ) ;
assign n35453 =  ( n148 ) ? ( n7266 ) : ( VREG_11_10 ) ;
assign n35454 =  ( n146 ) ? ( n7265 ) : ( n35453 ) ;
assign n35455 =  ( n144 ) ? ( n7264 ) : ( n35454 ) ;
assign n35456 =  ( n142 ) ? ( n7263 ) : ( n35455 ) ;
assign n35457 =  ( n10 ) ? ( n7262 ) : ( n35456 ) ;
assign n35458 =  ( n7273 ) ? ( VREG_11_10 ) : ( n35452 ) ;
assign n35459 =  ( n7273 ) ? ( VREG_11_10 ) : ( n35457 ) ;
assign n35460 =  ( n3034 ) ? ( n35459 ) : ( VREG_11_10 ) ;
assign n35461 =  ( n2965 ) ? ( n35458 ) : ( n35460 ) ;
assign n35462 =  ( n1930 ) ? ( n35457 ) : ( n35461 ) ;
assign n35463 =  ( n879 ) ? ( n35452 ) : ( n35462 ) ;
assign n35464 =  ( n172 ) ? ( n7284 ) : ( VREG_11_10 ) ;
assign n35465 =  ( n170 ) ? ( n7283 ) : ( n35464 ) ;
assign n35466 =  ( n168 ) ? ( n7282 ) : ( n35465 ) ;
assign n35467 =  ( n166 ) ? ( n7281 ) : ( n35466 ) ;
assign n35468 =  ( n162 ) ? ( n7280 ) : ( n35467 ) ;
assign n35469 =  ( n172 ) ? ( n7294 ) : ( VREG_11_10 ) ;
assign n35470 =  ( n170 ) ? ( n7293 ) : ( n35469 ) ;
assign n35471 =  ( n168 ) ? ( n7292 ) : ( n35470 ) ;
assign n35472 =  ( n166 ) ? ( n7291 ) : ( n35471 ) ;
assign n35473 =  ( n162 ) ? ( n7290 ) : ( n35472 ) ;
assign n35474 =  ( n7273 ) ? ( VREG_11_10 ) : ( n35473 ) ;
assign n35475 =  ( n3051 ) ? ( n35474 ) : ( VREG_11_10 ) ;
assign n35476 =  ( n3040 ) ? ( n35468 ) : ( n35475 ) ;
assign n35477 =  ( n192 ) ? ( VREG_11_10 ) : ( VREG_11_10 ) ;
assign n35478 =  ( n157 ) ? ( n35476 ) : ( n35477 ) ;
assign n35479 =  ( n6 ) ? ( n35463 ) : ( n35478 ) ;
assign n35480 =  ( n241 ) ? ( n35479 ) : ( VREG_11_10 ) ;
assign n35481 =  ( n148 ) ? ( n8351 ) : ( VREG_11_11 ) ;
assign n35482 =  ( n146 ) ? ( n8350 ) : ( n35481 ) ;
assign n35483 =  ( n144 ) ? ( n8349 ) : ( n35482 ) ;
assign n35484 =  ( n142 ) ? ( n8348 ) : ( n35483 ) ;
assign n35485 =  ( n10 ) ? ( n8347 ) : ( n35484 ) ;
assign n35486 =  ( n148 ) ? ( n9385 ) : ( VREG_11_11 ) ;
assign n35487 =  ( n146 ) ? ( n9384 ) : ( n35486 ) ;
assign n35488 =  ( n144 ) ? ( n9383 ) : ( n35487 ) ;
assign n35489 =  ( n142 ) ? ( n9382 ) : ( n35488 ) ;
assign n35490 =  ( n10 ) ? ( n9381 ) : ( n35489 ) ;
assign n35491 =  ( n9392 ) ? ( VREG_11_11 ) : ( n35485 ) ;
assign n35492 =  ( n9392 ) ? ( VREG_11_11 ) : ( n35490 ) ;
assign n35493 =  ( n3034 ) ? ( n35492 ) : ( VREG_11_11 ) ;
assign n35494 =  ( n2965 ) ? ( n35491 ) : ( n35493 ) ;
assign n35495 =  ( n1930 ) ? ( n35490 ) : ( n35494 ) ;
assign n35496 =  ( n879 ) ? ( n35485 ) : ( n35495 ) ;
assign n35497 =  ( n172 ) ? ( n9403 ) : ( VREG_11_11 ) ;
assign n35498 =  ( n170 ) ? ( n9402 ) : ( n35497 ) ;
assign n35499 =  ( n168 ) ? ( n9401 ) : ( n35498 ) ;
assign n35500 =  ( n166 ) ? ( n9400 ) : ( n35499 ) ;
assign n35501 =  ( n162 ) ? ( n9399 ) : ( n35500 ) ;
assign n35502 =  ( n172 ) ? ( n9413 ) : ( VREG_11_11 ) ;
assign n35503 =  ( n170 ) ? ( n9412 ) : ( n35502 ) ;
assign n35504 =  ( n168 ) ? ( n9411 ) : ( n35503 ) ;
assign n35505 =  ( n166 ) ? ( n9410 ) : ( n35504 ) ;
assign n35506 =  ( n162 ) ? ( n9409 ) : ( n35505 ) ;
assign n35507 =  ( n9392 ) ? ( VREG_11_11 ) : ( n35506 ) ;
assign n35508 =  ( n3051 ) ? ( n35507 ) : ( VREG_11_11 ) ;
assign n35509 =  ( n3040 ) ? ( n35501 ) : ( n35508 ) ;
assign n35510 =  ( n192 ) ? ( VREG_11_11 ) : ( VREG_11_11 ) ;
assign n35511 =  ( n157 ) ? ( n35509 ) : ( n35510 ) ;
assign n35512 =  ( n6 ) ? ( n35496 ) : ( n35511 ) ;
assign n35513 =  ( n241 ) ? ( n35512 ) : ( VREG_11_11 ) ;
assign n35514 =  ( n148 ) ? ( n10470 ) : ( VREG_11_12 ) ;
assign n35515 =  ( n146 ) ? ( n10469 ) : ( n35514 ) ;
assign n35516 =  ( n144 ) ? ( n10468 ) : ( n35515 ) ;
assign n35517 =  ( n142 ) ? ( n10467 ) : ( n35516 ) ;
assign n35518 =  ( n10 ) ? ( n10466 ) : ( n35517 ) ;
assign n35519 =  ( n148 ) ? ( n11504 ) : ( VREG_11_12 ) ;
assign n35520 =  ( n146 ) ? ( n11503 ) : ( n35519 ) ;
assign n35521 =  ( n144 ) ? ( n11502 ) : ( n35520 ) ;
assign n35522 =  ( n142 ) ? ( n11501 ) : ( n35521 ) ;
assign n35523 =  ( n10 ) ? ( n11500 ) : ( n35522 ) ;
assign n35524 =  ( n11511 ) ? ( VREG_11_12 ) : ( n35518 ) ;
assign n35525 =  ( n11511 ) ? ( VREG_11_12 ) : ( n35523 ) ;
assign n35526 =  ( n3034 ) ? ( n35525 ) : ( VREG_11_12 ) ;
assign n35527 =  ( n2965 ) ? ( n35524 ) : ( n35526 ) ;
assign n35528 =  ( n1930 ) ? ( n35523 ) : ( n35527 ) ;
assign n35529 =  ( n879 ) ? ( n35518 ) : ( n35528 ) ;
assign n35530 =  ( n172 ) ? ( n11522 ) : ( VREG_11_12 ) ;
assign n35531 =  ( n170 ) ? ( n11521 ) : ( n35530 ) ;
assign n35532 =  ( n168 ) ? ( n11520 ) : ( n35531 ) ;
assign n35533 =  ( n166 ) ? ( n11519 ) : ( n35532 ) ;
assign n35534 =  ( n162 ) ? ( n11518 ) : ( n35533 ) ;
assign n35535 =  ( n172 ) ? ( n11532 ) : ( VREG_11_12 ) ;
assign n35536 =  ( n170 ) ? ( n11531 ) : ( n35535 ) ;
assign n35537 =  ( n168 ) ? ( n11530 ) : ( n35536 ) ;
assign n35538 =  ( n166 ) ? ( n11529 ) : ( n35537 ) ;
assign n35539 =  ( n162 ) ? ( n11528 ) : ( n35538 ) ;
assign n35540 =  ( n11511 ) ? ( VREG_11_12 ) : ( n35539 ) ;
assign n35541 =  ( n3051 ) ? ( n35540 ) : ( VREG_11_12 ) ;
assign n35542 =  ( n3040 ) ? ( n35534 ) : ( n35541 ) ;
assign n35543 =  ( n192 ) ? ( VREG_11_12 ) : ( VREG_11_12 ) ;
assign n35544 =  ( n157 ) ? ( n35542 ) : ( n35543 ) ;
assign n35545 =  ( n6 ) ? ( n35529 ) : ( n35544 ) ;
assign n35546 =  ( n241 ) ? ( n35545 ) : ( VREG_11_12 ) ;
assign n35547 =  ( n148 ) ? ( n12589 ) : ( VREG_11_13 ) ;
assign n35548 =  ( n146 ) ? ( n12588 ) : ( n35547 ) ;
assign n35549 =  ( n144 ) ? ( n12587 ) : ( n35548 ) ;
assign n35550 =  ( n142 ) ? ( n12586 ) : ( n35549 ) ;
assign n35551 =  ( n10 ) ? ( n12585 ) : ( n35550 ) ;
assign n35552 =  ( n148 ) ? ( n13623 ) : ( VREG_11_13 ) ;
assign n35553 =  ( n146 ) ? ( n13622 ) : ( n35552 ) ;
assign n35554 =  ( n144 ) ? ( n13621 ) : ( n35553 ) ;
assign n35555 =  ( n142 ) ? ( n13620 ) : ( n35554 ) ;
assign n35556 =  ( n10 ) ? ( n13619 ) : ( n35555 ) ;
assign n35557 =  ( n13630 ) ? ( VREG_11_13 ) : ( n35551 ) ;
assign n35558 =  ( n13630 ) ? ( VREG_11_13 ) : ( n35556 ) ;
assign n35559 =  ( n3034 ) ? ( n35558 ) : ( VREG_11_13 ) ;
assign n35560 =  ( n2965 ) ? ( n35557 ) : ( n35559 ) ;
assign n35561 =  ( n1930 ) ? ( n35556 ) : ( n35560 ) ;
assign n35562 =  ( n879 ) ? ( n35551 ) : ( n35561 ) ;
assign n35563 =  ( n172 ) ? ( n13641 ) : ( VREG_11_13 ) ;
assign n35564 =  ( n170 ) ? ( n13640 ) : ( n35563 ) ;
assign n35565 =  ( n168 ) ? ( n13639 ) : ( n35564 ) ;
assign n35566 =  ( n166 ) ? ( n13638 ) : ( n35565 ) ;
assign n35567 =  ( n162 ) ? ( n13637 ) : ( n35566 ) ;
assign n35568 =  ( n172 ) ? ( n13651 ) : ( VREG_11_13 ) ;
assign n35569 =  ( n170 ) ? ( n13650 ) : ( n35568 ) ;
assign n35570 =  ( n168 ) ? ( n13649 ) : ( n35569 ) ;
assign n35571 =  ( n166 ) ? ( n13648 ) : ( n35570 ) ;
assign n35572 =  ( n162 ) ? ( n13647 ) : ( n35571 ) ;
assign n35573 =  ( n13630 ) ? ( VREG_11_13 ) : ( n35572 ) ;
assign n35574 =  ( n3051 ) ? ( n35573 ) : ( VREG_11_13 ) ;
assign n35575 =  ( n3040 ) ? ( n35567 ) : ( n35574 ) ;
assign n35576 =  ( n192 ) ? ( VREG_11_13 ) : ( VREG_11_13 ) ;
assign n35577 =  ( n157 ) ? ( n35575 ) : ( n35576 ) ;
assign n35578 =  ( n6 ) ? ( n35562 ) : ( n35577 ) ;
assign n35579 =  ( n241 ) ? ( n35578 ) : ( VREG_11_13 ) ;
assign n35580 =  ( n148 ) ? ( n14708 ) : ( VREG_11_14 ) ;
assign n35581 =  ( n146 ) ? ( n14707 ) : ( n35580 ) ;
assign n35582 =  ( n144 ) ? ( n14706 ) : ( n35581 ) ;
assign n35583 =  ( n142 ) ? ( n14705 ) : ( n35582 ) ;
assign n35584 =  ( n10 ) ? ( n14704 ) : ( n35583 ) ;
assign n35585 =  ( n148 ) ? ( n15742 ) : ( VREG_11_14 ) ;
assign n35586 =  ( n146 ) ? ( n15741 ) : ( n35585 ) ;
assign n35587 =  ( n144 ) ? ( n15740 ) : ( n35586 ) ;
assign n35588 =  ( n142 ) ? ( n15739 ) : ( n35587 ) ;
assign n35589 =  ( n10 ) ? ( n15738 ) : ( n35588 ) ;
assign n35590 =  ( n15749 ) ? ( VREG_11_14 ) : ( n35584 ) ;
assign n35591 =  ( n15749 ) ? ( VREG_11_14 ) : ( n35589 ) ;
assign n35592 =  ( n3034 ) ? ( n35591 ) : ( VREG_11_14 ) ;
assign n35593 =  ( n2965 ) ? ( n35590 ) : ( n35592 ) ;
assign n35594 =  ( n1930 ) ? ( n35589 ) : ( n35593 ) ;
assign n35595 =  ( n879 ) ? ( n35584 ) : ( n35594 ) ;
assign n35596 =  ( n172 ) ? ( n15760 ) : ( VREG_11_14 ) ;
assign n35597 =  ( n170 ) ? ( n15759 ) : ( n35596 ) ;
assign n35598 =  ( n168 ) ? ( n15758 ) : ( n35597 ) ;
assign n35599 =  ( n166 ) ? ( n15757 ) : ( n35598 ) ;
assign n35600 =  ( n162 ) ? ( n15756 ) : ( n35599 ) ;
assign n35601 =  ( n172 ) ? ( n15770 ) : ( VREG_11_14 ) ;
assign n35602 =  ( n170 ) ? ( n15769 ) : ( n35601 ) ;
assign n35603 =  ( n168 ) ? ( n15768 ) : ( n35602 ) ;
assign n35604 =  ( n166 ) ? ( n15767 ) : ( n35603 ) ;
assign n35605 =  ( n162 ) ? ( n15766 ) : ( n35604 ) ;
assign n35606 =  ( n15749 ) ? ( VREG_11_14 ) : ( n35605 ) ;
assign n35607 =  ( n3051 ) ? ( n35606 ) : ( VREG_11_14 ) ;
assign n35608 =  ( n3040 ) ? ( n35600 ) : ( n35607 ) ;
assign n35609 =  ( n192 ) ? ( VREG_11_14 ) : ( VREG_11_14 ) ;
assign n35610 =  ( n157 ) ? ( n35608 ) : ( n35609 ) ;
assign n35611 =  ( n6 ) ? ( n35595 ) : ( n35610 ) ;
assign n35612 =  ( n241 ) ? ( n35611 ) : ( VREG_11_14 ) ;
assign n35613 =  ( n148 ) ? ( n16827 ) : ( VREG_11_15 ) ;
assign n35614 =  ( n146 ) ? ( n16826 ) : ( n35613 ) ;
assign n35615 =  ( n144 ) ? ( n16825 ) : ( n35614 ) ;
assign n35616 =  ( n142 ) ? ( n16824 ) : ( n35615 ) ;
assign n35617 =  ( n10 ) ? ( n16823 ) : ( n35616 ) ;
assign n35618 =  ( n148 ) ? ( n17861 ) : ( VREG_11_15 ) ;
assign n35619 =  ( n146 ) ? ( n17860 ) : ( n35618 ) ;
assign n35620 =  ( n144 ) ? ( n17859 ) : ( n35619 ) ;
assign n35621 =  ( n142 ) ? ( n17858 ) : ( n35620 ) ;
assign n35622 =  ( n10 ) ? ( n17857 ) : ( n35621 ) ;
assign n35623 =  ( n17868 ) ? ( VREG_11_15 ) : ( n35617 ) ;
assign n35624 =  ( n17868 ) ? ( VREG_11_15 ) : ( n35622 ) ;
assign n35625 =  ( n3034 ) ? ( n35624 ) : ( VREG_11_15 ) ;
assign n35626 =  ( n2965 ) ? ( n35623 ) : ( n35625 ) ;
assign n35627 =  ( n1930 ) ? ( n35622 ) : ( n35626 ) ;
assign n35628 =  ( n879 ) ? ( n35617 ) : ( n35627 ) ;
assign n35629 =  ( n172 ) ? ( n17879 ) : ( VREG_11_15 ) ;
assign n35630 =  ( n170 ) ? ( n17878 ) : ( n35629 ) ;
assign n35631 =  ( n168 ) ? ( n17877 ) : ( n35630 ) ;
assign n35632 =  ( n166 ) ? ( n17876 ) : ( n35631 ) ;
assign n35633 =  ( n162 ) ? ( n17875 ) : ( n35632 ) ;
assign n35634 =  ( n172 ) ? ( n17889 ) : ( VREG_11_15 ) ;
assign n35635 =  ( n170 ) ? ( n17888 ) : ( n35634 ) ;
assign n35636 =  ( n168 ) ? ( n17887 ) : ( n35635 ) ;
assign n35637 =  ( n166 ) ? ( n17886 ) : ( n35636 ) ;
assign n35638 =  ( n162 ) ? ( n17885 ) : ( n35637 ) ;
assign n35639 =  ( n17868 ) ? ( VREG_11_15 ) : ( n35638 ) ;
assign n35640 =  ( n3051 ) ? ( n35639 ) : ( VREG_11_15 ) ;
assign n35641 =  ( n3040 ) ? ( n35633 ) : ( n35640 ) ;
assign n35642 =  ( n192 ) ? ( VREG_11_15 ) : ( VREG_11_15 ) ;
assign n35643 =  ( n157 ) ? ( n35641 ) : ( n35642 ) ;
assign n35644 =  ( n6 ) ? ( n35628 ) : ( n35643 ) ;
assign n35645 =  ( n241 ) ? ( n35644 ) : ( VREG_11_15 ) ;
assign n35646 =  ( n148 ) ? ( n18946 ) : ( VREG_11_2 ) ;
assign n35647 =  ( n146 ) ? ( n18945 ) : ( n35646 ) ;
assign n35648 =  ( n144 ) ? ( n18944 ) : ( n35647 ) ;
assign n35649 =  ( n142 ) ? ( n18943 ) : ( n35648 ) ;
assign n35650 =  ( n10 ) ? ( n18942 ) : ( n35649 ) ;
assign n35651 =  ( n148 ) ? ( n19980 ) : ( VREG_11_2 ) ;
assign n35652 =  ( n146 ) ? ( n19979 ) : ( n35651 ) ;
assign n35653 =  ( n144 ) ? ( n19978 ) : ( n35652 ) ;
assign n35654 =  ( n142 ) ? ( n19977 ) : ( n35653 ) ;
assign n35655 =  ( n10 ) ? ( n19976 ) : ( n35654 ) ;
assign n35656 =  ( n19987 ) ? ( VREG_11_2 ) : ( n35650 ) ;
assign n35657 =  ( n19987 ) ? ( VREG_11_2 ) : ( n35655 ) ;
assign n35658 =  ( n3034 ) ? ( n35657 ) : ( VREG_11_2 ) ;
assign n35659 =  ( n2965 ) ? ( n35656 ) : ( n35658 ) ;
assign n35660 =  ( n1930 ) ? ( n35655 ) : ( n35659 ) ;
assign n35661 =  ( n879 ) ? ( n35650 ) : ( n35660 ) ;
assign n35662 =  ( n172 ) ? ( n19998 ) : ( VREG_11_2 ) ;
assign n35663 =  ( n170 ) ? ( n19997 ) : ( n35662 ) ;
assign n35664 =  ( n168 ) ? ( n19996 ) : ( n35663 ) ;
assign n35665 =  ( n166 ) ? ( n19995 ) : ( n35664 ) ;
assign n35666 =  ( n162 ) ? ( n19994 ) : ( n35665 ) ;
assign n35667 =  ( n172 ) ? ( n20008 ) : ( VREG_11_2 ) ;
assign n35668 =  ( n170 ) ? ( n20007 ) : ( n35667 ) ;
assign n35669 =  ( n168 ) ? ( n20006 ) : ( n35668 ) ;
assign n35670 =  ( n166 ) ? ( n20005 ) : ( n35669 ) ;
assign n35671 =  ( n162 ) ? ( n20004 ) : ( n35670 ) ;
assign n35672 =  ( n19987 ) ? ( VREG_11_2 ) : ( n35671 ) ;
assign n35673 =  ( n3051 ) ? ( n35672 ) : ( VREG_11_2 ) ;
assign n35674 =  ( n3040 ) ? ( n35666 ) : ( n35673 ) ;
assign n35675 =  ( n192 ) ? ( VREG_11_2 ) : ( VREG_11_2 ) ;
assign n35676 =  ( n157 ) ? ( n35674 ) : ( n35675 ) ;
assign n35677 =  ( n6 ) ? ( n35661 ) : ( n35676 ) ;
assign n35678 =  ( n241 ) ? ( n35677 ) : ( VREG_11_2 ) ;
assign n35679 =  ( n148 ) ? ( n21065 ) : ( VREG_11_3 ) ;
assign n35680 =  ( n146 ) ? ( n21064 ) : ( n35679 ) ;
assign n35681 =  ( n144 ) ? ( n21063 ) : ( n35680 ) ;
assign n35682 =  ( n142 ) ? ( n21062 ) : ( n35681 ) ;
assign n35683 =  ( n10 ) ? ( n21061 ) : ( n35682 ) ;
assign n35684 =  ( n148 ) ? ( n22099 ) : ( VREG_11_3 ) ;
assign n35685 =  ( n146 ) ? ( n22098 ) : ( n35684 ) ;
assign n35686 =  ( n144 ) ? ( n22097 ) : ( n35685 ) ;
assign n35687 =  ( n142 ) ? ( n22096 ) : ( n35686 ) ;
assign n35688 =  ( n10 ) ? ( n22095 ) : ( n35687 ) ;
assign n35689 =  ( n22106 ) ? ( VREG_11_3 ) : ( n35683 ) ;
assign n35690 =  ( n22106 ) ? ( VREG_11_3 ) : ( n35688 ) ;
assign n35691 =  ( n3034 ) ? ( n35690 ) : ( VREG_11_3 ) ;
assign n35692 =  ( n2965 ) ? ( n35689 ) : ( n35691 ) ;
assign n35693 =  ( n1930 ) ? ( n35688 ) : ( n35692 ) ;
assign n35694 =  ( n879 ) ? ( n35683 ) : ( n35693 ) ;
assign n35695 =  ( n172 ) ? ( n22117 ) : ( VREG_11_3 ) ;
assign n35696 =  ( n170 ) ? ( n22116 ) : ( n35695 ) ;
assign n35697 =  ( n168 ) ? ( n22115 ) : ( n35696 ) ;
assign n35698 =  ( n166 ) ? ( n22114 ) : ( n35697 ) ;
assign n35699 =  ( n162 ) ? ( n22113 ) : ( n35698 ) ;
assign n35700 =  ( n172 ) ? ( n22127 ) : ( VREG_11_3 ) ;
assign n35701 =  ( n170 ) ? ( n22126 ) : ( n35700 ) ;
assign n35702 =  ( n168 ) ? ( n22125 ) : ( n35701 ) ;
assign n35703 =  ( n166 ) ? ( n22124 ) : ( n35702 ) ;
assign n35704 =  ( n162 ) ? ( n22123 ) : ( n35703 ) ;
assign n35705 =  ( n22106 ) ? ( VREG_11_3 ) : ( n35704 ) ;
assign n35706 =  ( n3051 ) ? ( n35705 ) : ( VREG_11_3 ) ;
assign n35707 =  ( n3040 ) ? ( n35699 ) : ( n35706 ) ;
assign n35708 =  ( n192 ) ? ( VREG_11_3 ) : ( VREG_11_3 ) ;
assign n35709 =  ( n157 ) ? ( n35707 ) : ( n35708 ) ;
assign n35710 =  ( n6 ) ? ( n35694 ) : ( n35709 ) ;
assign n35711 =  ( n241 ) ? ( n35710 ) : ( VREG_11_3 ) ;
assign n35712 =  ( n148 ) ? ( n23184 ) : ( VREG_11_4 ) ;
assign n35713 =  ( n146 ) ? ( n23183 ) : ( n35712 ) ;
assign n35714 =  ( n144 ) ? ( n23182 ) : ( n35713 ) ;
assign n35715 =  ( n142 ) ? ( n23181 ) : ( n35714 ) ;
assign n35716 =  ( n10 ) ? ( n23180 ) : ( n35715 ) ;
assign n35717 =  ( n148 ) ? ( n24218 ) : ( VREG_11_4 ) ;
assign n35718 =  ( n146 ) ? ( n24217 ) : ( n35717 ) ;
assign n35719 =  ( n144 ) ? ( n24216 ) : ( n35718 ) ;
assign n35720 =  ( n142 ) ? ( n24215 ) : ( n35719 ) ;
assign n35721 =  ( n10 ) ? ( n24214 ) : ( n35720 ) ;
assign n35722 =  ( n24225 ) ? ( VREG_11_4 ) : ( n35716 ) ;
assign n35723 =  ( n24225 ) ? ( VREG_11_4 ) : ( n35721 ) ;
assign n35724 =  ( n3034 ) ? ( n35723 ) : ( VREG_11_4 ) ;
assign n35725 =  ( n2965 ) ? ( n35722 ) : ( n35724 ) ;
assign n35726 =  ( n1930 ) ? ( n35721 ) : ( n35725 ) ;
assign n35727 =  ( n879 ) ? ( n35716 ) : ( n35726 ) ;
assign n35728 =  ( n172 ) ? ( n24236 ) : ( VREG_11_4 ) ;
assign n35729 =  ( n170 ) ? ( n24235 ) : ( n35728 ) ;
assign n35730 =  ( n168 ) ? ( n24234 ) : ( n35729 ) ;
assign n35731 =  ( n166 ) ? ( n24233 ) : ( n35730 ) ;
assign n35732 =  ( n162 ) ? ( n24232 ) : ( n35731 ) ;
assign n35733 =  ( n172 ) ? ( n24246 ) : ( VREG_11_4 ) ;
assign n35734 =  ( n170 ) ? ( n24245 ) : ( n35733 ) ;
assign n35735 =  ( n168 ) ? ( n24244 ) : ( n35734 ) ;
assign n35736 =  ( n166 ) ? ( n24243 ) : ( n35735 ) ;
assign n35737 =  ( n162 ) ? ( n24242 ) : ( n35736 ) ;
assign n35738 =  ( n24225 ) ? ( VREG_11_4 ) : ( n35737 ) ;
assign n35739 =  ( n3051 ) ? ( n35738 ) : ( VREG_11_4 ) ;
assign n35740 =  ( n3040 ) ? ( n35732 ) : ( n35739 ) ;
assign n35741 =  ( n192 ) ? ( VREG_11_4 ) : ( VREG_11_4 ) ;
assign n35742 =  ( n157 ) ? ( n35740 ) : ( n35741 ) ;
assign n35743 =  ( n6 ) ? ( n35727 ) : ( n35742 ) ;
assign n35744 =  ( n241 ) ? ( n35743 ) : ( VREG_11_4 ) ;
assign n35745 =  ( n148 ) ? ( n25303 ) : ( VREG_11_5 ) ;
assign n35746 =  ( n146 ) ? ( n25302 ) : ( n35745 ) ;
assign n35747 =  ( n144 ) ? ( n25301 ) : ( n35746 ) ;
assign n35748 =  ( n142 ) ? ( n25300 ) : ( n35747 ) ;
assign n35749 =  ( n10 ) ? ( n25299 ) : ( n35748 ) ;
assign n35750 =  ( n148 ) ? ( n26337 ) : ( VREG_11_5 ) ;
assign n35751 =  ( n146 ) ? ( n26336 ) : ( n35750 ) ;
assign n35752 =  ( n144 ) ? ( n26335 ) : ( n35751 ) ;
assign n35753 =  ( n142 ) ? ( n26334 ) : ( n35752 ) ;
assign n35754 =  ( n10 ) ? ( n26333 ) : ( n35753 ) ;
assign n35755 =  ( n26344 ) ? ( VREG_11_5 ) : ( n35749 ) ;
assign n35756 =  ( n26344 ) ? ( VREG_11_5 ) : ( n35754 ) ;
assign n35757 =  ( n3034 ) ? ( n35756 ) : ( VREG_11_5 ) ;
assign n35758 =  ( n2965 ) ? ( n35755 ) : ( n35757 ) ;
assign n35759 =  ( n1930 ) ? ( n35754 ) : ( n35758 ) ;
assign n35760 =  ( n879 ) ? ( n35749 ) : ( n35759 ) ;
assign n35761 =  ( n172 ) ? ( n26355 ) : ( VREG_11_5 ) ;
assign n35762 =  ( n170 ) ? ( n26354 ) : ( n35761 ) ;
assign n35763 =  ( n168 ) ? ( n26353 ) : ( n35762 ) ;
assign n35764 =  ( n166 ) ? ( n26352 ) : ( n35763 ) ;
assign n35765 =  ( n162 ) ? ( n26351 ) : ( n35764 ) ;
assign n35766 =  ( n172 ) ? ( n26365 ) : ( VREG_11_5 ) ;
assign n35767 =  ( n170 ) ? ( n26364 ) : ( n35766 ) ;
assign n35768 =  ( n168 ) ? ( n26363 ) : ( n35767 ) ;
assign n35769 =  ( n166 ) ? ( n26362 ) : ( n35768 ) ;
assign n35770 =  ( n162 ) ? ( n26361 ) : ( n35769 ) ;
assign n35771 =  ( n26344 ) ? ( VREG_11_5 ) : ( n35770 ) ;
assign n35772 =  ( n3051 ) ? ( n35771 ) : ( VREG_11_5 ) ;
assign n35773 =  ( n3040 ) ? ( n35765 ) : ( n35772 ) ;
assign n35774 =  ( n192 ) ? ( VREG_11_5 ) : ( VREG_11_5 ) ;
assign n35775 =  ( n157 ) ? ( n35773 ) : ( n35774 ) ;
assign n35776 =  ( n6 ) ? ( n35760 ) : ( n35775 ) ;
assign n35777 =  ( n241 ) ? ( n35776 ) : ( VREG_11_5 ) ;
assign n35778 =  ( n148 ) ? ( n27422 ) : ( VREG_11_6 ) ;
assign n35779 =  ( n146 ) ? ( n27421 ) : ( n35778 ) ;
assign n35780 =  ( n144 ) ? ( n27420 ) : ( n35779 ) ;
assign n35781 =  ( n142 ) ? ( n27419 ) : ( n35780 ) ;
assign n35782 =  ( n10 ) ? ( n27418 ) : ( n35781 ) ;
assign n35783 =  ( n148 ) ? ( n28456 ) : ( VREG_11_6 ) ;
assign n35784 =  ( n146 ) ? ( n28455 ) : ( n35783 ) ;
assign n35785 =  ( n144 ) ? ( n28454 ) : ( n35784 ) ;
assign n35786 =  ( n142 ) ? ( n28453 ) : ( n35785 ) ;
assign n35787 =  ( n10 ) ? ( n28452 ) : ( n35786 ) ;
assign n35788 =  ( n28463 ) ? ( VREG_11_6 ) : ( n35782 ) ;
assign n35789 =  ( n28463 ) ? ( VREG_11_6 ) : ( n35787 ) ;
assign n35790 =  ( n3034 ) ? ( n35789 ) : ( VREG_11_6 ) ;
assign n35791 =  ( n2965 ) ? ( n35788 ) : ( n35790 ) ;
assign n35792 =  ( n1930 ) ? ( n35787 ) : ( n35791 ) ;
assign n35793 =  ( n879 ) ? ( n35782 ) : ( n35792 ) ;
assign n35794 =  ( n172 ) ? ( n28474 ) : ( VREG_11_6 ) ;
assign n35795 =  ( n170 ) ? ( n28473 ) : ( n35794 ) ;
assign n35796 =  ( n168 ) ? ( n28472 ) : ( n35795 ) ;
assign n35797 =  ( n166 ) ? ( n28471 ) : ( n35796 ) ;
assign n35798 =  ( n162 ) ? ( n28470 ) : ( n35797 ) ;
assign n35799 =  ( n172 ) ? ( n28484 ) : ( VREG_11_6 ) ;
assign n35800 =  ( n170 ) ? ( n28483 ) : ( n35799 ) ;
assign n35801 =  ( n168 ) ? ( n28482 ) : ( n35800 ) ;
assign n35802 =  ( n166 ) ? ( n28481 ) : ( n35801 ) ;
assign n35803 =  ( n162 ) ? ( n28480 ) : ( n35802 ) ;
assign n35804 =  ( n28463 ) ? ( VREG_11_6 ) : ( n35803 ) ;
assign n35805 =  ( n3051 ) ? ( n35804 ) : ( VREG_11_6 ) ;
assign n35806 =  ( n3040 ) ? ( n35798 ) : ( n35805 ) ;
assign n35807 =  ( n192 ) ? ( VREG_11_6 ) : ( VREG_11_6 ) ;
assign n35808 =  ( n157 ) ? ( n35806 ) : ( n35807 ) ;
assign n35809 =  ( n6 ) ? ( n35793 ) : ( n35808 ) ;
assign n35810 =  ( n241 ) ? ( n35809 ) : ( VREG_11_6 ) ;
assign n35811 =  ( n148 ) ? ( n29541 ) : ( VREG_11_7 ) ;
assign n35812 =  ( n146 ) ? ( n29540 ) : ( n35811 ) ;
assign n35813 =  ( n144 ) ? ( n29539 ) : ( n35812 ) ;
assign n35814 =  ( n142 ) ? ( n29538 ) : ( n35813 ) ;
assign n35815 =  ( n10 ) ? ( n29537 ) : ( n35814 ) ;
assign n35816 =  ( n148 ) ? ( n30575 ) : ( VREG_11_7 ) ;
assign n35817 =  ( n146 ) ? ( n30574 ) : ( n35816 ) ;
assign n35818 =  ( n144 ) ? ( n30573 ) : ( n35817 ) ;
assign n35819 =  ( n142 ) ? ( n30572 ) : ( n35818 ) ;
assign n35820 =  ( n10 ) ? ( n30571 ) : ( n35819 ) ;
assign n35821 =  ( n30582 ) ? ( VREG_11_7 ) : ( n35815 ) ;
assign n35822 =  ( n30582 ) ? ( VREG_11_7 ) : ( n35820 ) ;
assign n35823 =  ( n3034 ) ? ( n35822 ) : ( VREG_11_7 ) ;
assign n35824 =  ( n2965 ) ? ( n35821 ) : ( n35823 ) ;
assign n35825 =  ( n1930 ) ? ( n35820 ) : ( n35824 ) ;
assign n35826 =  ( n879 ) ? ( n35815 ) : ( n35825 ) ;
assign n35827 =  ( n172 ) ? ( n30593 ) : ( VREG_11_7 ) ;
assign n35828 =  ( n170 ) ? ( n30592 ) : ( n35827 ) ;
assign n35829 =  ( n168 ) ? ( n30591 ) : ( n35828 ) ;
assign n35830 =  ( n166 ) ? ( n30590 ) : ( n35829 ) ;
assign n35831 =  ( n162 ) ? ( n30589 ) : ( n35830 ) ;
assign n35832 =  ( n172 ) ? ( n30603 ) : ( VREG_11_7 ) ;
assign n35833 =  ( n170 ) ? ( n30602 ) : ( n35832 ) ;
assign n35834 =  ( n168 ) ? ( n30601 ) : ( n35833 ) ;
assign n35835 =  ( n166 ) ? ( n30600 ) : ( n35834 ) ;
assign n35836 =  ( n162 ) ? ( n30599 ) : ( n35835 ) ;
assign n35837 =  ( n30582 ) ? ( VREG_11_7 ) : ( n35836 ) ;
assign n35838 =  ( n3051 ) ? ( n35837 ) : ( VREG_11_7 ) ;
assign n35839 =  ( n3040 ) ? ( n35831 ) : ( n35838 ) ;
assign n35840 =  ( n192 ) ? ( VREG_11_7 ) : ( VREG_11_7 ) ;
assign n35841 =  ( n157 ) ? ( n35839 ) : ( n35840 ) ;
assign n35842 =  ( n6 ) ? ( n35826 ) : ( n35841 ) ;
assign n35843 =  ( n241 ) ? ( n35842 ) : ( VREG_11_7 ) ;
assign n35844 =  ( n148 ) ? ( n31660 ) : ( VREG_11_8 ) ;
assign n35845 =  ( n146 ) ? ( n31659 ) : ( n35844 ) ;
assign n35846 =  ( n144 ) ? ( n31658 ) : ( n35845 ) ;
assign n35847 =  ( n142 ) ? ( n31657 ) : ( n35846 ) ;
assign n35848 =  ( n10 ) ? ( n31656 ) : ( n35847 ) ;
assign n35849 =  ( n148 ) ? ( n32694 ) : ( VREG_11_8 ) ;
assign n35850 =  ( n146 ) ? ( n32693 ) : ( n35849 ) ;
assign n35851 =  ( n144 ) ? ( n32692 ) : ( n35850 ) ;
assign n35852 =  ( n142 ) ? ( n32691 ) : ( n35851 ) ;
assign n35853 =  ( n10 ) ? ( n32690 ) : ( n35852 ) ;
assign n35854 =  ( n32701 ) ? ( VREG_11_8 ) : ( n35848 ) ;
assign n35855 =  ( n32701 ) ? ( VREG_11_8 ) : ( n35853 ) ;
assign n35856 =  ( n3034 ) ? ( n35855 ) : ( VREG_11_8 ) ;
assign n35857 =  ( n2965 ) ? ( n35854 ) : ( n35856 ) ;
assign n35858 =  ( n1930 ) ? ( n35853 ) : ( n35857 ) ;
assign n35859 =  ( n879 ) ? ( n35848 ) : ( n35858 ) ;
assign n35860 =  ( n172 ) ? ( n32712 ) : ( VREG_11_8 ) ;
assign n35861 =  ( n170 ) ? ( n32711 ) : ( n35860 ) ;
assign n35862 =  ( n168 ) ? ( n32710 ) : ( n35861 ) ;
assign n35863 =  ( n166 ) ? ( n32709 ) : ( n35862 ) ;
assign n35864 =  ( n162 ) ? ( n32708 ) : ( n35863 ) ;
assign n35865 =  ( n172 ) ? ( n32722 ) : ( VREG_11_8 ) ;
assign n35866 =  ( n170 ) ? ( n32721 ) : ( n35865 ) ;
assign n35867 =  ( n168 ) ? ( n32720 ) : ( n35866 ) ;
assign n35868 =  ( n166 ) ? ( n32719 ) : ( n35867 ) ;
assign n35869 =  ( n162 ) ? ( n32718 ) : ( n35868 ) ;
assign n35870 =  ( n32701 ) ? ( VREG_11_8 ) : ( n35869 ) ;
assign n35871 =  ( n3051 ) ? ( n35870 ) : ( VREG_11_8 ) ;
assign n35872 =  ( n3040 ) ? ( n35864 ) : ( n35871 ) ;
assign n35873 =  ( n192 ) ? ( VREG_11_8 ) : ( VREG_11_8 ) ;
assign n35874 =  ( n157 ) ? ( n35872 ) : ( n35873 ) ;
assign n35875 =  ( n6 ) ? ( n35859 ) : ( n35874 ) ;
assign n35876 =  ( n241 ) ? ( n35875 ) : ( VREG_11_8 ) ;
assign n35877 =  ( n148 ) ? ( n33779 ) : ( VREG_11_9 ) ;
assign n35878 =  ( n146 ) ? ( n33778 ) : ( n35877 ) ;
assign n35879 =  ( n144 ) ? ( n33777 ) : ( n35878 ) ;
assign n35880 =  ( n142 ) ? ( n33776 ) : ( n35879 ) ;
assign n35881 =  ( n10 ) ? ( n33775 ) : ( n35880 ) ;
assign n35882 =  ( n148 ) ? ( n34813 ) : ( VREG_11_9 ) ;
assign n35883 =  ( n146 ) ? ( n34812 ) : ( n35882 ) ;
assign n35884 =  ( n144 ) ? ( n34811 ) : ( n35883 ) ;
assign n35885 =  ( n142 ) ? ( n34810 ) : ( n35884 ) ;
assign n35886 =  ( n10 ) ? ( n34809 ) : ( n35885 ) ;
assign n35887 =  ( n34820 ) ? ( VREG_11_9 ) : ( n35881 ) ;
assign n35888 =  ( n34820 ) ? ( VREG_11_9 ) : ( n35886 ) ;
assign n35889 =  ( n3034 ) ? ( n35888 ) : ( VREG_11_9 ) ;
assign n35890 =  ( n2965 ) ? ( n35887 ) : ( n35889 ) ;
assign n35891 =  ( n1930 ) ? ( n35886 ) : ( n35890 ) ;
assign n35892 =  ( n879 ) ? ( n35881 ) : ( n35891 ) ;
assign n35893 =  ( n172 ) ? ( n34831 ) : ( VREG_11_9 ) ;
assign n35894 =  ( n170 ) ? ( n34830 ) : ( n35893 ) ;
assign n35895 =  ( n168 ) ? ( n34829 ) : ( n35894 ) ;
assign n35896 =  ( n166 ) ? ( n34828 ) : ( n35895 ) ;
assign n35897 =  ( n162 ) ? ( n34827 ) : ( n35896 ) ;
assign n35898 =  ( n172 ) ? ( n34841 ) : ( VREG_11_9 ) ;
assign n35899 =  ( n170 ) ? ( n34840 ) : ( n35898 ) ;
assign n35900 =  ( n168 ) ? ( n34839 ) : ( n35899 ) ;
assign n35901 =  ( n166 ) ? ( n34838 ) : ( n35900 ) ;
assign n35902 =  ( n162 ) ? ( n34837 ) : ( n35901 ) ;
assign n35903 =  ( n34820 ) ? ( VREG_11_9 ) : ( n35902 ) ;
assign n35904 =  ( n3051 ) ? ( n35903 ) : ( VREG_11_9 ) ;
assign n35905 =  ( n3040 ) ? ( n35897 ) : ( n35904 ) ;
assign n35906 =  ( n192 ) ? ( VREG_11_9 ) : ( VREG_11_9 ) ;
assign n35907 =  ( n157 ) ? ( n35905 ) : ( n35906 ) ;
assign n35908 =  ( n6 ) ? ( n35892 ) : ( n35907 ) ;
assign n35909 =  ( n241 ) ? ( n35908 ) : ( VREG_11_9 ) ;
assign n35910 =  ( n148 ) ? ( n1924 ) : ( VREG_12_0 ) ;
assign n35911 =  ( n146 ) ? ( n1923 ) : ( n35910 ) ;
assign n35912 =  ( n144 ) ? ( n1922 ) : ( n35911 ) ;
assign n35913 =  ( n142 ) ? ( n1921 ) : ( n35912 ) ;
assign n35914 =  ( n10 ) ? ( n1920 ) : ( n35913 ) ;
assign n35915 =  ( n148 ) ? ( n2959 ) : ( VREG_12_0 ) ;
assign n35916 =  ( n146 ) ? ( n2958 ) : ( n35915 ) ;
assign n35917 =  ( n144 ) ? ( n2957 ) : ( n35916 ) ;
assign n35918 =  ( n142 ) ? ( n2956 ) : ( n35917 ) ;
assign n35919 =  ( n10 ) ? ( n2955 ) : ( n35918 ) ;
assign n35920 =  ( n3032 ) ? ( VREG_12_0 ) : ( n35914 ) ;
assign n35921 =  ( n3032 ) ? ( VREG_12_0 ) : ( n35919 ) ;
assign n35922 =  ( n3034 ) ? ( n35921 ) : ( VREG_12_0 ) ;
assign n35923 =  ( n2965 ) ? ( n35920 ) : ( n35922 ) ;
assign n35924 =  ( n1930 ) ? ( n35919 ) : ( n35923 ) ;
assign n35925 =  ( n879 ) ? ( n35914 ) : ( n35924 ) ;
assign n35926 =  ( n172 ) ? ( n3045 ) : ( VREG_12_0 ) ;
assign n35927 =  ( n170 ) ? ( n3044 ) : ( n35926 ) ;
assign n35928 =  ( n168 ) ? ( n3043 ) : ( n35927 ) ;
assign n35929 =  ( n166 ) ? ( n3042 ) : ( n35928 ) ;
assign n35930 =  ( n162 ) ? ( n3041 ) : ( n35929 ) ;
assign n35931 =  ( n172 ) ? ( n3056 ) : ( VREG_12_0 ) ;
assign n35932 =  ( n170 ) ? ( n3055 ) : ( n35931 ) ;
assign n35933 =  ( n168 ) ? ( n3054 ) : ( n35932 ) ;
assign n35934 =  ( n166 ) ? ( n3053 ) : ( n35933 ) ;
assign n35935 =  ( n162 ) ? ( n3052 ) : ( n35934 ) ;
assign n35936 =  ( n3032 ) ? ( VREG_12_0 ) : ( n35935 ) ;
assign n35937 =  ( n3051 ) ? ( n35936 ) : ( VREG_12_0 ) ;
assign n35938 =  ( n3040 ) ? ( n35930 ) : ( n35937 ) ;
assign n35939 =  ( n192 ) ? ( VREG_12_0 ) : ( VREG_12_0 ) ;
assign n35940 =  ( n157 ) ? ( n35938 ) : ( n35939 ) ;
assign n35941 =  ( n6 ) ? ( n35925 ) : ( n35940 ) ;
assign n35942 =  ( n263 ) ? ( n35941 ) : ( VREG_12_0 ) ;
assign n35943 =  ( n148 ) ? ( n4113 ) : ( VREG_12_1 ) ;
assign n35944 =  ( n146 ) ? ( n4112 ) : ( n35943 ) ;
assign n35945 =  ( n144 ) ? ( n4111 ) : ( n35944 ) ;
assign n35946 =  ( n142 ) ? ( n4110 ) : ( n35945 ) ;
assign n35947 =  ( n10 ) ? ( n4109 ) : ( n35946 ) ;
assign n35948 =  ( n148 ) ? ( n5147 ) : ( VREG_12_1 ) ;
assign n35949 =  ( n146 ) ? ( n5146 ) : ( n35948 ) ;
assign n35950 =  ( n144 ) ? ( n5145 ) : ( n35949 ) ;
assign n35951 =  ( n142 ) ? ( n5144 ) : ( n35950 ) ;
assign n35952 =  ( n10 ) ? ( n5143 ) : ( n35951 ) ;
assign n35953 =  ( n5154 ) ? ( VREG_12_1 ) : ( n35947 ) ;
assign n35954 =  ( n5154 ) ? ( VREG_12_1 ) : ( n35952 ) ;
assign n35955 =  ( n3034 ) ? ( n35954 ) : ( VREG_12_1 ) ;
assign n35956 =  ( n2965 ) ? ( n35953 ) : ( n35955 ) ;
assign n35957 =  ( n1930 ) ? ( n35952 ) : ( n35956 ) ;
assign n35958 =  ( n879 ) ? ( n35947 ) : ( n35957 ) ;
assign n35959 =  ( n172 ) ? ( n5165 ) : ( VREG_12_1 ) ;
assign n35960 =  ( n170 ) ? ( n5164 ) : ( n35959 ) ;
assign n35961 =  ( n168 ) ? ( n5163 ) : ( n35960 ) ;
assign n35962 =  ( n166 ) ? ( n5162 ) : ( n35961 ) ;
assign n35963 =  ( n162 ) ? ( n5161 ) : ( n35962 ) ;
assign n35964 =  ( n172 ) ? ( n5175 ) : ( VREG_12_1 ) ;
assign n35965 =  ( n170 ) ? ( n5174 ) : ( n35964 ) ;
assign n35966 =  ( n168 ) ? ( n5173 ) : ( n35965 ) ;
assign n35967 =  ( n166 ) ? ( n5172 ) : ( n35966 ) ;
assign n35968 =  ( n162 ) ? ( n5171 ) : ( n35967 ) ;
assign n35969 =  ( n5154 ) ? ( VREG_12_1 ) : ( n35968 ) ;
assign n35970 =  ( n3051 ) ? ( n35969 ) : ( VREG_12_1 ) ;
assign n35971 =  ( n3040 ) ? ( n35963 ) : ( n35970 ) ;
assign n35972 =  ( n192 ) ? ( VREG_12_1 ) : ( VREG_12_1 ) ;
assign n35973 =  ( n157 ) ? ( n35971 ) : ( n35972 ) ;
assign n35974 =  ( n6 ) ? ( n35958 ) : ( n35973 ) ;
assign n35975 =  ( n263 ) ? ( n35974 ) : ( VREG_12_1 ) ;
assign n35976 =  ( n148 ) ? ( n6232 ) : ( VREG_12_10 ) ;
assign n35977 =  ( n146 ) ? ( n6231 ) : ( n35976 ) ;
assign n35978 =  ( n144 ) ? ( n6230 ) : ( n35977 ) ;
assign n35979 =  ( n142 ) ? ( n6229 ) : ( n35978 ) ;
assign n35980 =  ( n10 ) ? ( n6228 ) : ( n35979 ) ;
assign n35981 =  ( n148 ) ? ( n7266 ) : ( VREG_12_10 ) ;
assign n35982 =  ( n146 ) ? ( n7265 ) : ( n35981 ) ;
assign n35983 =  ( n144 ) ? ( n7264 ) : ( n35982 ) ;
assign n35984 =  ( n142 ) ? ( n7263 ) : ( n35983 ) ;
assign n35985 =  ( n10 ) ? ( n7262 ) : ( n35984 ) ;
assign n35986 =  ( n7273 ) ? ( VREG_12_10 ) : ( n35980 ) ;
assign n35987 =  ( n7273 ) ? ( VREG_12_10 ) : ( n35985 ) ;
assign n35988 =  ( n3034 ) ? ( n35987 ) : ( VREG_12_10 ) ;
assign n35989 =  ( n2965 ) ? ( n35986 ) : ( n35988 ) ;
assign n35990 =  ( n1930 ) ? ( n35985 ) : ( n35989 ) ;
assign n35991 =  ( n879 ) ? ( n35980 ) : ( n35990 ) ;
assign n35992 =  ( n172 ) ? ( n7284 ) : ( VREG_12_10 ) ;
assign n35993 =  ( n170 ) ? ( n7283 ) : ( n35992 ) ;
assign n35994 =  ( n168 ) ? ( n7282 ) : ( n35993 ) ;
assign n35995 =  ( n166 ) ? ( n7281 ) : ( n35994 ) ;
assign n35996 =  ( n162 ) ? ( n7280 ) : ( n35995 ) ;
assign n35997 =  ( n172 ) ? ( n7294 ) : ( VREG_12_10 ) ;
assign n35998 =  ( n170 ) ? ( n7293 ) : ( n35997 ) ;
assign n35999 =  ( n168 ) ? ( n7292 ) : ( n35998 ) ;
assign n36000 =  ( n166 ) ? ( n7291 ) : ( n35999 ) ;
assign n36001 =  ( n162 ) ? ( n7290 ) : ( n36000 ) ;
assign n36002 =  ( n7273 ) ? ( VREG_12_10 ) : ( n36001 ) ;
assign n36003 =  ( n3051 ) ? ( n36002 ) : ( VREG_12_10 ) ;
assign n36004 =  ( n3040 ) ? ( n35996 ) : ( n36003 ) ;
assign n36005 =  ( n192 ) ? ( VREG_12_10 ) : ( VREG_12_10 ) ;
assign n36006 =  ( n157 ) ? ( n36004 ) : ( n36005 ) ;
assign n36007 =  ( n6 ) ? ( n35991 ) : ( n36006 ) ;
assign n36008 =  ( n263 ) ? ( n36007 ) : ( VREG_12_10 ) ;
assign n36009 =  ( n148 ) ? ( n8351 ) : ( VREG_12_11 ) ;
assign n36010 =  ( n146 ) ? ( n8350 ) : ( n36009 ) ;
assign n36011 =  ( n144 ) ? ( n8349 ) : ( n36010 ) ;
assign n36012 =  ( n142 ) ? ( n8348 ) : ( n36011 ) ;
assign n36013 =  ( n10 ) ? ( n8347 ) : ( n36012 ) ;
assign n36014 =  ( n148 ) ? ( n9385 ) : ( VREG_12_11 ) ;
assign n36015 =  ( n146 ) ? ( n9384 ) : ( n36014 ) ;
assign n36016 =  ( n144 ) ? ( n9383 ) : ( n36015 ) ;
assign n36017 =  ( n142 ) ? ( n9382 ) : ( n36016 ) ;
assign n36018 =  ( n10 ) ? ( n9381 ) : ( n36017 ) ;
assign n36019 =  ( n9392 ) ? ( VREG_12_11 ) : ( n36013 ) ;
assign n36020 =  ( n9392 ) ? ( VREG_12_11 ) : ( n36018 ) ;
assign n36021 =  ( n3034 ) ? ( n36020 ) : ( VREG_12_11 ) ;
assign n36022 =  ( n2965 ) ? ( n36019 ) : ( n36021 ) ;
assign n36023 =  ( n1930 ) ? ( n36018 ) : ( n36022 ) ;
assign n36024 =  ( n879 ) ? ( n36013 ) : ( n36023 ) ;
assign n36025 =  ( n172 ) ? ( n9403 ) : ( VREG_12_11 ) ;
assign n36026 =  ( n170 ) ? ( n9402 ) : ( n36025 ) ;
assign n36027 =  ( n168 ) ? ( n9401 ) : ( n36026 ) ;
assign n36028 =  ( n166 ) ? ( n9400 ) : ( n36027 ) ;
assign n36029 =  ( n162 ) ? ( n9399 ) : ( n36028 ) ;
assign n36030 =  ( n172 ) ? ( n9413 ) : ( VREG_12_11 ) ;
assign n36031 =  ( n170 ) ? ( n9412 ) : ( n36030 ) ;
assign n36032 =  ( n168 ) ? ( n9411 ) : ( n36031 ) ;
assign n36033 =  ( n166 ) ? ( n9410 ) : ( n36032 ) ;
assign n36034 =  ( n162 ) ? ( n9409 ) : ( n36033 ) ;
assign n36035 =  ( n9392 ) ? ( VREG_12_11 ) : ( n36034 ) ;
assign n36036 =  ( n3051 ) ? ( n36035 ) : ( VREG_12_11 ) ;
assign n36037 =  ( n3040 ) ? ( n36029 ) : ( n36036 ) ;
assign n36038 =  ( n192 ) ? ( VREG_12_11 ) : ( VREG_12_11 ) ;
assign n36039 =  ( n157 ) ? ( n36037 ) : ( n36038 ) ;
assign n36040 =  ( n6 ) ? ( n36024 ) : ( n36039 ) ;
assign n36041 =  ( n263 ) ? ( n36040 ) : ( VREG_12_11 ) ;
assign n36042 =  ( n148 ) ? ( n10470 ) : ( VREG_12_12 ) ;
assign n36043 =  ( n146 ) ? ( n10469 ) : ( n36042 ) ;
assign n36044 =  ( n144 ) ? ( n10468 ) : ( n36043 ) ;
assign n36045 =  ( n142 ) ? ( n10467 ) : ( n36044 ) ;
assign n36046 =  ( n10 ) ? ( n10466 ) : ( n36045 ) ;
assign n36047 =  ( n148 ) ? ( n11504 ) : ( VREG_12_12 ) ;
assign n36048 =  ( n146 ) ? ( n11503 ) : ( n36047 ) ;
assign n36049 =  ( n144 ) ? ( n11502 ) : ( n36048 ) ;
assign n36050 =  ( n142 ) ? ( n11501 ) : ( n36049 ) ;
assign n36051 =  ( n10 ) ? ( n11500 ) : ( n36050 ) ;
assign n36052 =  ( n11511 ) ? ( VREG_12_12 ) : ( n36046 ) ;
assign n36053 =  ( n11511 ) ? ( VREG_12_12 ) : ( n36051 ) ;
assign n36054 =  ( n3034 ) ? ( n36053 ) : ( VREG_12_12 ) ;
assign n36055 =  ( n2965 ) ? ( n36052 ) : ( n36054 ) ;
assign n36056 =  ( n1930 ) ? ( n36051 ) : ( n36055 ) ;
assign n36057 =  ( n879 ) ? ( n36046 ) : ( n36056 ) ;
assign n36058 =  ( n172 ) ? ( n11522 ) : ( VREG_12_12 ) ;
assign n36059 =  ( n170 ) ? ( n11521 ) : ( n36058 ) ;
assign n36060 =  ( n168 ) ? ( n11520 ) : ( n36059 ) ;
assign n36061 =  ( n166 ) ? ( n11519 ) : ( n36060 ) ;
assign n36062 =  ( n162 ) ? ( n11518 ) : ( n36061 ) ;
assign n36063 =  ( n172 ) ? ( n11532 ) : ( VREG_12_12 ) ;
assign n36064 =  ( n170 ) ? ( n11531 ) : ( n36063 ) ;
assign n36065 =  ( n168 ) ? ( n11530 ) : ( n36064 ) ;
assign n36066 =  ( n166 ) ? ( n11529 ) : ( n36065 ) ;
assign n36067 =  ( n162 ) ? ( n11528 ) : ( n36066 ) ;
assign n36068 =  ( n11511 ) ? ( VREG_12_12 ) : ( n36067 ) ;
assign n36069 =  ( n3051 ) ? ( n36068 ) : ( VREG_12_12 ) ;
assign n36070 =  ( n3040 ) ? ( n36062 ) : ( n36069 ) ;
assign n36071 =  ( n192 ) ? ( VREG_12_12 ) : ( VREG_12_12 ) ;
assign n36072 =  ( n157 ) ? ( n36070 ) : ( n36071 ) ;
assign n36073 =  ( n6 ) ? ( n36057 ) : ( n36072 ) ;
assign n36074 =  ( n263 ) ? ( n36073 ) : ( VREG_12_12 ) ;
assign n36075 =  ( n148 ) ? ( n12589 ) : ( VREG_12_13 ) ;
assign n36076 =  ( n146 ) ? ( n12588 ) : ( n36075 ) ;
assign n36077 =  ( n144 ) ? ( n12587 ) : ( n36076 ) ;
assign n36078 =  ( n142 ) ? ( n12586 ) : ( n36077 ) ;
assign n36079 =  ( n10 ) ? ( n12585 ) : ( n36078 ) ;
assign n36080 =  ( n148 ) ? ( n13623 ) : ( VREG_12_13 ) ;
assign n36081 =  ( n146 ) ? ( n13622 ) : ( n36080 ) ;
assign n36082 =  ( n144 ) ? ( n13621 ) : ( n36081 ) ;
assign n36083 =  ( n142 ) ? ( n13620 ) : ( n36082 ) ;
assign n36084 =  ( n10 ) ? ( n13619 ) : ( n36083 ) ;
assign n36085 =  ( n13630 ) ? ( VREG_12_13 ) : ( n36079 ) ;
assign n36086 =  ( n13630 ) ? ( VREG_12_13 ) : ( n36084 ) ;
assign n36087 =  ( n3034 ) ? ( n36086 ) : ( VREG_12_13 ) ;
assign n36088 =  ( n2965 ) ? ( n36085 ) : ( n36087 ) ;
assign n36089 =  ( n1930 ) ? ( n36084 ) : ( n36088 ) ;
assign n36090 =  ( n879 ) ? ( n36079 ) : ( n36089 ) ;
assign n36091 =  ( n172 ) ? ( n13641 ) : ( VREG_12_13 ) ;
assign n36092 =  ( n170 ) ? ( n13640 ) : ( n36091 ) ;
assign n36093 =  ( n168 ) ? ( n13639 ) : ( n36092 ) ;
assign n36094 =  ( n166 ) ? ( n13638 ) : ( n36093 ) ;
assign n36095 =  ( n162 ) ? ( n13637 ) : ( n36094 ) ;
assign n36096 =  ( n172 ) ? ( n13651 ) : ( VREG_12_13 ) ;
assign n36097 =  ( n170 ) ? ( n13650 ) : ( n36096 ) ;
assign n36098 =  ( n168 ) ? ( n13649 ) : ( n36097 ) ;
assign n36099 =  ( n166 ) ? ( n13648 ) : ( n36098 ) ;
assign n36100 =  ( n162 ) ? ( n13647 ) : ( n36099 ) ;
assign n36101 =  ( n13630 ) ? ( VREG_12_13 ) : ( n36100 ) ;
assign n36102 =  ( n3051 ) ? ( n36101 ) : ( VREG_12_13 ) ;
assign n36103 =  ( n3040 ) ? ( n36095 ) : ( n36102 ) ;
assign n36104 =  ( n192 ) ? ( VREG_12_13 ) : ( VREG_12_13 ) ;
assign n36105 =  ( n157 ) ? ( n36103 ) : ( n36104 ) ;
assign n36106 =  ( n6 ) ? ( n36090 ) : ( n36105 ) ;
assign n36107 =  ( n263 ) ? ( n36106 ) : ( VREG_12_13 ) ;
assign n36108 =  ( n148 ) ? ( n14708 ) : ( VREG_12_14 ) ;
assign n36109 =  ( n146 ) ? ( n14707 ) : ( n36108 ) ;
assign n36110 =  ( n144 ) ? ( n14706 ) : ( n36109 ) ;
assign n36111 =  ( n142 ) ? ( n14705 ) : ( n36110 ) ;
assign n36112 =  ( n10 ) ? ( n14704 ) : ( n36111 ) ;
assign n36113 =  ( n148 ) ? ( n15742 ) : ( VREG_12_14 ) ;
assign n36114 =  ( n146 ) ? ( n15741 ) : ( n36113 ) ;
assign n36115 =  ( n144 ) ? ( n15740 ) : ( n36114 ) ;
assign n36116 =  ( n142 ) ? ( n15739 ) : ( n36115 ) ;
assign n36117 =  ( n10 ) ? ( n15738 ) : ( n36116 ) ;
assign n36118 =  ( n15749 ) ? ( VREG_12_14 ) : ( n36112 ) ;
assign n36119 =  ( n15749 ) ? ( VREG_12_14 ) : ( n36117 ) ;
assign n36120 =  ( n3034 ) ? ( n36119 ) : ( VREG_12_14 ) ;
assign n36121 =  ( n2965 ) ? ( n36118 ) : ( n36120 ) ;
assign n36122 =  ( n1930 ) ? ( n36117 ) : ( n36121 ) ;
assign n36123 =  ( n879 ) ? ( n36112 ) : ( n36122 ) ;
assign n36124 =  ( n172 ) ? ( n15760 ) : ( VREG_12_14 ) ;
assign n36125 =  ( n170 ) ? ( n15759 ) : ( n36124 ) ;
assign n36126 =  ( n168 ) ? ( n15758 ) : ( n36125 ) ;
assign n36127 =  ( n166 ) ? ( n15757 ) : ( n36126 ) ;
assign n36128 =  ( n162 ) ? ( n15756 ) : ( n36127 ) ;
assign n36129 =  ( n172 ) ? ( n15770 ) : ( VREG_12_14 ) ;
assign n36130 =  ( n170 ) ? ( n15769 ) : ( n36129 ) ;
assign n36131 =  ( n168 ) ? ( n15768 ) : ( n36130 ) ;
assign n36132 =  ( n166 ) ? ( n15767 ) : ( n36131 ) ;
assign n36133 =  ( n162 ) ? ( n15766 ) : ( n36132 ) ;
assign n36134 =  ( n15749 ) ? ( VREG_12_14 ) : ( n36133 ) ;
assign n36135 =  ( n3051 ) ? ( n36134 ) : ( VREG_12_14 ) ;
assign n36136 =  ( n3040 ) ? ( n36128 ) : ( n36135 ) ;
assign n36137 =  ( n192 ) ? ( VREG_12_14 ) : ( VREG_12_14 ) ;
assign n36138 =  ( n157 ) ? ( n36136 ) : ( n36137 ) ;
assign n36139 =  ( n6 ) ? ( n36123 ) : ( n36138 ) ;
assign n36140 =  ( n263 ) ? ( n36139 ) : ( VREG_12_14 ) ;
assign n36141 =  ( n148 ) ? ( n16827 ) : ( VREG_12_15 ) ;
assign n36142 =  ( n146 ) ? ( n16826 ) : ( n36141 ) ;
assign n36143 =  ( n144 ) ? ( n16825 ) : ( n36142 ) ;
assign n36144 =  ( n142 ) ? ( n16824 ) : ( n36143 ) ;
assign n36145 =  ( n10 ) ? ( n16823 ) : ( n36144 ) ;
assign n36146 =  ( n148 ) ? ( n17861 ) : ( VREG_12_15 ) ;
assign n36147 =  ( n146 ) ? ( n17860 ) : ( n36146 ) ;
assign n36148 =  ( n144 ) ? ( n17859 ) : ( n36147 ) ;
assign n36149 =  ( n142 ) ? ( n17858 ) : ( n36148 ) ;
assign n36150 =  ( n10 ) ? ( n17857 ) : ( n36149 ) ;
assign n36151 =  ( n17868 ) ? ( VREG_12_15 ) : ( n36145 ) ;
assign n36152 =  ( n17868 ) ? ( VREG_12_15 ) : ( n36150 ) ;
assign n36153 =  ( n3034 ) ? ( n36152 ) : ( VREG_12_15 ) ;
assign n36154 =  ( n2965 ) ? ( n36151 ) : ( n36153 ) ;
assign n36155 =  ( n1930 ) ? ( n36150 ) : ( n36154 ) ;
assign n36156 =  ( n879 ) ? ( n36145 ) : ( n36155 ) ;
assign n36157 =  ( n172 ) ? ( n17879 ) : ( VREG_12_15 ) ;
assign n36158 =  ( n170 ) ? ( n17878 ) : ( n36157 ) ;
assign n36159 =  ( n168 ) ? ( n17877 ) : ( n36158 ) ;
assign n36160 =  ( n166 ) ? ( n17876 ) : ( n36159 ) ;
assign n36161 =  ( n162 ) ? ( n17875 ) : ( n36160 ) ;
assign n36162 =  ( n172 ) ? ( n17889 ) : ( VREG_12_15 ) ;
assign n36163 =  ( n170 ) ? ( n17888 ) : ( n36162 ) ;
assign n36164 =  ( n168 ) ? ( n17887 ) : ( n36163 ) ;
assign n36165 =  ( n166 ) ? ( n17886 ) : ( n36164 ) ;
assign n36166 =  ( n162 ) ? ( n17885 ) : ( n36165 ) ;
assign n36167 =  ( n17868 ) ? ( VREG_12_15 ) : ( n36166 ) ;
assign n36168 =  ( n3051 ) ? ( n36167 ) : ( VREG_12_15 ) ;
assign n36169 =  ( n3040 ) ? ( n36161 ) : ( n36168 ) ;
assign n36170 =  ( n192 ) ? ( VREG_12_15 ) : ( VREG_12_15 ) ;
assign n36171 =  ( n157 ) ? ( n36169 ) : ( n36170 ) ;
assign n36172 =  ( n6 ) ? ( n36156 ) : ( n36171 ) ;
assign n36173 =  ( n263 ) ? ( n36172 ) : ( VREG_12_15 ) ;
assign n36174 =  ( n148 ) ? ( n18946 ) : ( VREG_12_2 ) ;
assign n36175 =  ( n146 ) ? ( n18945 ) : ( n36174 ) ;
assign n36176 =  ( n144 ) ? ( n18944 ) : ( n36175 ) ;
assign n36177 =  ( n142 ) ? ( n18943 ) : ( n36176 ) ;
assign n36178 =  ( n10 ) ? ( n18942 ) : ( n36177 ) ;
assign n36179 =  ( n148 ) ? ( n19980 ) : ( VREG_12_2 ) ;
assign n36180 =  ( n146 ) ? ( n19979 ) : ( n36179 ) ;
assign n36181 =  ( n144 ) ? ( n19978 ) : ( n36180 ) ;
assign n36182 =  ( n142 ) ? ( n19977 ) : ( n36181 ) ;
assign n36183 =  ( n10 ) ? ( n19976 ) : ( n36182 ) ;
assign n36184 =  ( n19987 ) ? ( VREG_12_2 ) : ( n36178 ) ;
assign n36185 =  ( n19987 ) ? ( VREG_12_2 ) : ( n36183 ) ;
assign n36186 =  ( n3034 ) ? ( n36185 ) : ( VREG_12_2 ) ;
assign n36187 =  ( n2965 ) ? ( n36184 ) : ( n36186 ) ;
assign n36188 =  ( n1930 ) ? ( n36183 ) : ( n36187 ) ;
assign n36189 =  ( n879 ) ? ( n36178 ) : ( n36188 ) ;
assign n36190 =  ( n172 ) ? ( n19998 ) : ( VREG_12_2 ) ;
assign n36191 =  ( n170 ) ? ( n19997 ) : ( n36190 ) ;
assign n36192 =  ( n168 ) ? ( n19996 ) : ( n36191 ) ;
assign n36193 =  ( n166 ) ? ( n19995 ) : ( n36192 ) ;
assign n36194 =  ( n162 ) ? ( n19994 ) : ( n36193 ) ;
assign n36195 =  ( n172 ) ? ( n20008 ) : ( VREG_12_2 ) ;
assign n36196 =  ( n170 ) ? ( n20007 ) : ( n36195 ) ;
assign n36197 =  ( n168 ) ? ( n20006 ) : ( n36196 ) ;
assign n36198 =  ( n166 ) ? ( n20005 ) : ( n36197 ) ;
assign n36199 =  ( n162 ) ? ( n20004 ) : ( n36198 ) ;
assign n36200 =  ( n19987 ) ? ( VREG_12_2 ) : ( n36199 ) ;
assign n36201 =  ( n3051 ) ? ( n36200 ) : ( VREG_12_2 ) ;
assign n36202 =  ( n3040 ) ? ( n36194 ) : ( n36201 ) ;
assign n36203 =  ( n192 ) ? ( VREG_12_2 ) : ( VREG_12_2 ) ;
assign n36204 =  ( n157 ) ? ( n36202 ) : ( n36203 ) ;
assign n36205 =  ( n6 ) ? ( n36189 ) : ( n36204 ) ;
assign n36206 =  ( n263 ) ? ( n36205 ) : ( VREG_12_2 ) ;
assign n36207 =  ( n148 ) ? ( n21065 ) : ( VREG_12_3 ) ;
assign n36208 =  ( n146 ) ? ( n21064 ) : ( n36207 ) ;
assign n36209 =  ( n144 ) ? ( n21063 ) : ( n36208 ) ;
assign n36210 =  ( n142 ) ? ( n21062 ) : ( n36209 ) ;
assign n36211 =  ( n10 ) ? ( n21061 ) : ( n36210 ) ;
assign n36212 =  ( n148 ) ? ( n22099 ) : ( VREG_12_3 ) ;
assign n36213 =  ( n146 ) ? ( n22098 ) : ( n36212 ) ;
assign n36214 =  ( n144 ) ? ( n22097 ) : ( n36213 ) ;
assign n36215 =  ( n142 ) ? ( n22096 ) : ( n36214 ) ;
assign n36216 =  ( n10 ) ? ( n22095 ) : ( n36215 ) ;
assign n36217 =  ( n22106 ) ? ( VREG_12_3 ) : ( n36211 ) ;
assign n36218 =  ( n22106 ) ? ( VREG_12_3 ) : ( n36216 ) ;
assign n36219 =  ( n3034 ) ? ( n36218 ) : ( VREG_12_3 ) ;
assign n36220 =  ( n2965 ) ? ( n36217 ) : ( n36219 ) ;
assign n36221 =  ( n1930 ) ? ( n36216 ) : ( n36220 ) ;
assign n36222 =  ( n879 ) ? ( n36211 ) : ( n36221 ) ;
assign n36223 =  ( n172 ) ? ( n22117 ) : ( VREG_12_3 ) ;
assign n36224 =  ( n170 ) ? ( n22116 ) : ( n36223 ) ;
assign n36225 =  ( n168 ) ? ( n22115 ) : ( n36224 ) ;
assign n36226 =  ( n166 ) ? ( n22114 ) : ( n36225 ) ;
assign n36227 =  ( n162 ) ? ( n22113 ) : ( n36226 ) ;
assign n36228 =  ( n172 ) ? ( n22127 ) : ( VREG_12_3 ) ;
assign n36229 =  ( n170 ) ? ( n22126 ) : ( n36228 ) ;
assign n36230 =  ( n168 ) ? ( n22125 ) : ( n36229 ) ;
assign n36231 =  ( n166 ) ? ( n22124 ) : ( n36230 ) ;
assign n36232 =  ( n162 ) ? ( n22123 ) : ( n36231 ) ;
assign n36233 =  ( n22106 ) ? ( VREG_12_3 ) : ( n36232 ) ;
assign n36234 =  ( n3051 ) ? ( n36233 ) : ( VREG_12_3 ) ;
assign n36235 =  ( n3040 ) ? ( n36227 ) : ( n36234 ) ;
assign n36236 =  ( n192 ) ? ( VREG_12_3 ) : ( VREG_12_3 ) ;
assign n36237 =  ( n157 ) ? ( n36235 ) : ( n36236 ) ;
assign n36238 =  ( n6 ) ? ( n36222 ) : ( n36237 ) ;
assign n36239 =  ( n263 ) ? ( n36238 ) : ( VREG_12_3 ) ;
assign n36240 =  ( n148 ) ? ( n23184 ) : ( VREG_12_4 ) ;
assign n36241 =  ( n146 ) ? ( n23183 ) : ( n36240 ) ;
assign n36242 =  ( n144 ) ? ( n23182 ) : ( n36241 ) ;
assign n36243 =  ( n142 ) ? ( n23181 ) : ( n36242 ) ;
assign n36244 =  ( n10 ) ? ( n23180 ) : ( n36243 ) ;
assign n36245 =  ( n148 ) ? ( n24218 ) : ( VREG_12_4 ) ;
assign n36246 =  ( n146 ) ? ( n24217 ) : ( n36245 ) ;
assign n36247 =  ( n144 ) ? ( n24216 ) : ( n36246 ) ;
assign n36248 =  ( n142 ) ? ( n24215 ) : ( n36247 ) ;
assign n36249 =  ( n10 ) ? ( n24214 ) : ( n36248 ) ;
assign n36250 =  ( n24225 ) ? ( VREG_12_4 ) : ( n36244 ) ;
assign n36251 =  ( n24225 ) ? ( VREG_12_4 ) : ( n36249 ) ;
assign n36252 =  ( n3034 ) ? ( n36251 ) : ( VREG_12_4 ) ;
assign n36253 =  ( n2965 ) ? ( n36250 ) : ( n36252 ) ;
assign n36254 =  ( n1930 ) ? ( n36249 ) : ( n36253 ) ;
assign n36255 =  ( n879 ) ? ( n36244 ) : ( n36254 ) ;
assign n36256 =  ( n172 ) ? ( n24236 ) : ( VREG_12_4 ) ;
assign n36257 =  ( n170 ) ? ( n24235 ) : ( n36256 ) ;
assign n36258 =  ( n168 ) ? ( n24234 ) : ( n36257 ) ;
assign n36259 =  ( n166 ) ? ( n24233 ) : ( n36258 ) ;
assign n36260 =  ( n162 ) ? ( n24232 ) : ( n36259 ) ;
assign n36261 =  ( n172 ) ? ( n24246 ) : ( VREG_12_4 ) ;
assign n36262 =  ( n170 ) ? ( n24245 ) : ( n36261 ) ;
assign n36263 =  ( n168 ) ? ( n24244 ) : ( n36262 ) ;
assign n36264 =  ( n166 ) ? ( n24243 ) : ( n36263 ) ;
assign n36265 =  ( n162 ) ? ( n24242 ) : ( n36264 ) ;
assign n36266 =  ( n24225 ) ? ( VREG_12_4 ) : ( n36265 ) ;
assign n36267 =  ( n3051 ) ? ( n36266 ) : ( VREG_12_4 ) ;
assign n36268 =  ( n3040 ) ? ( n36260 ) : ( n36267 ) ;
assign n36269 =  ( n192 ) ? ( VREG_12_4 ) : ( VREG_12_4 ) ;
assign n36270 =  ( n157 ) ? ( n36268 ) : ( n36269 ) ;
assign n36271 =  ( n6 ) ? ( n36255 ) : ( n36270 ) ;
assign n36272 =  ( n263 ) ? ( n36271 ) : ( VREG_12_4 ) ;
assign n36273 =  ( n148 ) ? ( n25303 ) : ( VREG_12_5 ) ;
assign n36274 =  ( n146 ) ? ( n25302 ) : ( n36273 ) ;
assign n36275 =  ( n144 ) ? ( n25301 ) : ( n36274 ) ;
assign n36276 =  ( n142 ) ? ( n25300 ) : ( n36275 ) ;
assign n36277 =  ( n10 ) ? ( n25299 ) : ( n36276 ) ;
assign n36278 =  ( n148 ) ? ( n26337 ) : ( VREG_12_5 ) ;
assign n36279 =  ( n146 ) ? ( n26336 ) : ( n36278 ) ;
assign n36280 =  ( n144 ) ? ( n26335 ) : ( n36279 ) ;
assign n36281 =  ( n142 ) ? ( n26334 ) : ( n36280 ) ;
assign n36282 =  ( n10 ) ? ( n26333 ) : ( n36281 ) ;
assign n36283 =  ( n26344 ) ? ( VREG_12_5 ) : ( n36277 ) ;
assign n36284 =  ( n26344 ) ? ( VREG_12_5 ) : ( n36282 ) ;
assign n36285 =  ( n3034 ) ? ( n36284 ) : ( VREG_12_5 ) ;
assign n36286 =  ( n2965 ) ? ( n36283 ) : ( n36285 ) ;
assign n36287 =  ( n1930 ) ? ( n36282 ) : ( n36286 ) ;
assign n36288 =  ( n879 ) ? ( n36277 ) : ( n36287 ) ;
assign n36289 =  ( n172 ) ? ( n26355 ) : ( VREG_12_5 ) ;
assign n36290 =  ( n170 ) ? ( n26354 ) : ( n36289 ) ;
assign n36291 =  ( n168 ) ? ( n26353 ) : ( n36290 ) ;
assign n36292 =  ( n166 ) ? ( n26352 ) : ( n36291 ) ;
assign n36293 =  ( n162 ) ? ( n26351 ) : ( n36292 ) ;
assign n36294 =  ( n172 ) ? ( n26365 ) : ( VREG_12_5 ) ;
assign n36295 =  ( n170 ) ? ( n26364 ) : ( n36294 ) ;
assign n36296 =  ( n168 ) ? ( n26363 ) : ( n36295 ) ;
assign n36297 =  ( n166 ) ? ( n26362 ) : ( n36296 ) ;
assign n36298 =  ( n162 ) ? ( n26361 ) : ( n36297 ) ;
assign n36299 =  ( n26344 ) ? ( VREG_12_5 ) : ( n36298 ) ;
assign n36300 =  ( n3051 ) ? ( n36299 ) : ( VREG_12_5 ) ;
assign n36301 =  ( n3040 ) ? ( n36293 ) : ( n36300 ) ;
assign n36302 =  ( n192 ) ? ( VREG_12_5 ) : ( VREG_12_5 ) ;
assign n36303 =  ( n157 ) ? ( n36301 ) : ( n36302 ) ;
assign n36304 =  ( n6 ) ? ( n36288 ) : ( n36303 ) ;
assign n36305 =  ( n263 ) ? ( n36304 ) : ( VREG_12_5 ) ;
assign n36306 =  ( n148 ) ? ( n27422 ) : ( VREG_12_6 ) ;
assign n36307 =  ( n146 ) ? ( n27421 ) : ( n36306 ) ;
assign n36308 =  ( n144 ) ? ( n27420 ) : ( n36307 ) ;
assign n36309 =  ( n142 ) ? ( n27419 ) : ( n36308 ) ;
assign n36310 =  ( n10 ) ? ( n27418 ) : ( n36309 ) ;
assign n36311 =  ( n148 ) ? ( n28456 ) : ( VREG_12_6 ) ;
assign n36312 =  ( n146 ) ? ( n28455 ) : ( n36311 ) ;
assign n36313 =  ( n144 ) ? ( n28454 ) : ( n36312 ) ;
assign n36314 =  ( n142 ) ? ( n28453 ) : ( n36313 ) ;
assign n36315 =  ( n10 ) ? ( n28452 ) : ( n36314 ) ;
assign n36316 =  ( n28463 ) ? ( VREG_12_6 ) : ( n36310 ) ;
assign n36317 =  ( n28463 ) ? ( VREG_12_6 ) : ( n36315 ) ;
assign n36318 =  ( n3034 ) ? ( n36317 ) : ( VREG_12_6 ) ;
assign n36319 =  ( n2965 ) ? ( n36316 ) : ( n36318 ) ;
assign n36320 =  ( n1930 ) ? ( n36315 ) : ( n36319 ) ;
assign n36321 =  ( n879 ) ? ( n36310 ) : ( n36320 ) ;
assign n36322 =  ( n172 ) ? ( n28474 ) : ( VREG_12_6 ) ;
assign n36323 =  ( n170 ) ? ( n28473 ) : ( n36322 ) ;
assign n36324 =  ( n168 ) ? ( n28472 ) : ( n36323 ) ;
assign n36325 =  ( n166 ) ? ( n28471 ) : ( n36324 ) ;
assign n36326 =  ( n162 ) ? ( n28470 ) : ( n36325 ) ;
assign n36327 =  ( n172 ) ? ( n28484 ) : ( VREG_12_6 ) ;
assign n36328 =  ( n170 ) ? ( n28483 ) : ( n36327 ) ;
assign n36329 =  ( n168 ) ? ( n28482 ) : ( n36328 ) ;
assign n36330 =  ( n166 ) ? ( n28481 ) : ( n36329 ) ;
assign n36331 =  ( n162 ) ? ( n28480 ) : ( n36330 ) ;
assign n36332 =  ( n28463 ) ? ( VREG_12_6 ) : ( n36331 ) ;
assign n36333 =  ( n3051 ) ? ( n36332 ) : ( VREG_12_6 ) ;
assign n36334 =  ( n3040 ) ? ( n36326 ) : ( n36333 ) ;
assign n36335 =  ( n192 ) ? ( VREG_12_6 ) : ( VREG_12_6 ) ;
assign n36336 =  ( n157 ) ? ( n36334 ) : ( n36335 ) ;
assign n36337 =  ( n6 ) ? ( n36321 ) : ( n36336 ) ;
assign n36338 =  ( n263 ) ? ( n36337 ) : ( VREG_12_6 ) ;
assign n36339 =  ( n148 ) ? ( n29541 ) : ( VREG_12_7 ) ;
assign n36340 =  ( n146 ) ? ( n29540 ) : ( n36339 ) ;
assign n36341 =  ( n144 ) ? ( n29539 ) : ( n36340 ) ;
assign n36342 =  ( n142 ) ? ( n29538 ) : ( n36341 ) ;
assign n36343 =  ( n10 ) ? ( n29537 ) : ( n36342 ) ;
assign n36344 =  ( n148 ) ? ( n30575 ) : ( VREG_12_7 ) ;
assign n36345 =  ( n146 ) ? ( n30574 ) : ( n36344 ) ;
assign n36346 =  ( n144 ) ? ( n30573 ) : ( n36345 ) ;
assign n36347 =  ( n142 ) ? ( n30572 ) : ( n36346 ) ;
assign n36348 =  ( n10 ) ? ( n30571 ) : ( n36347 ) ;
assign n36349 =  ( n30582 ) ? ( VREG_12_7 ) : ( n36343 ) ;
assign n36350 =  ( n30582 ) ? ( VREG_12_7 ) : ( n36348 ) ;
assign n36351 =  ( n3034 ) ? ( n36350 ) : ( VREG_12_7 ) ;
assign n36352 =  ( n2965 ) ? ( n36349 ) : ( n36351 ) ;
assign n36353 =  ( n1930 ) ? ( n36348 ) : ( n36352 ) ;
assign n36354 =  ( n879 ) ? ( n36343 ) : ( n36353 ) ;
assign n36355 =  ( n172 ) ? ( n30593 ) : ( VREG_12_7 ) ;
assign n36356 =  ( n170 ) ? ( n30592 ) : ( n36355 ) ;
assign n36357 =  ( n168 ) ? ( n30591 ) : ( n36356 ) ;
assign n36358 =  ( n166 ) ? ( n30590 ) : ( n36357 ) ;
assign n36359 =  ( n162 ) ? ( n30589 ) : ( n36358 ) ;
assign n36360 =  ( n172 ) ? ( n30603 ) : ( VREG_12_7 ) ;
assign n36361 =  ( n170 ) ? ( n30602 ) : ( n36360 ) ;
assign n36362 =  ( n168 ) ? ( n30601 ) : ( n36361 ) ;
assign n36363 =  ( n166 ) ? ( n30600 ) : ( n36362 ) ;
assign n36364 =  ( n162 ) ? ( n30599 ) : ( n36363 ) ;
assign n36365 =  ( n30582 ) ? ( VREG_12_7 ) : ( n36364 ) ;
assign n36366 =  ( n3051 ) ? ( n36365 ) : ( VREG_12_7 ) ;
assign n36367 =  ( n3040 ) ? ( n36359 ) : ( n36366 ) ;
assign n36368 =  ( n192 ) ? ( VREG_12_7 ) : ( VREG_12_7 ) ;
assign n36369 =  ( n157 ) ? ( n36367 ) : ( n36368 ) ;
assign n36370 =  ( n6 ) ? ( n36354 ) : ( n36369 ) ;
assign n36371 =  ( n263 ) ? ( n36370 ) : ( VREG_12_7 ) ;
assign n36372 =  ( n148 ) ? ( n31660 ) : ( VREG_12_8 ) ;
assign n36373 =  ( n146 ) ? ( n31659 ) : ( n36372 ) ;
assign n36374 =  ( n144 ) ? ( n31658 ) : ( n36373 ) ;
assign n36375 =  ( n142 ) ? ( n31657 ) : ( n36374 ) ;
assign n36376 =  ( n10 ) ? ( n31656 ) : ( n36375 ) ;
assign n36377 =  ( n148 ) ? ( n32694 ) : ( VREG_12_8 ) ;
assign n36378 =  ( n146 ) ? ( n32693 ) : ( n36377 ) ;
assign n36379 =  ( n144 ) ? ( n32692 ) : ( n36378 ) ;
assign n36380 =  ( n142 ) ? ( n32691 ) : ( n36379 ) ;
assign n36381 =  ( n10 ) ? ( n32690 ) : ( n36380 ) ;
assign n36382 =  ( n32701 ) ? ( VREG_12_8 ) : ( n36376 ) ;
assign n36383 =  ( n32701 ) ? ( VREG_12_8 ) : ( n36381 ) ;
assign n36384 =  ( n3034 ) ? ( n36383 ) : ( VREG_12_8 ) ;
assign n36385 =  ( n2965 ) ? ( n36382 ) : ( n36384 ) ;
assign n36386 =  ( n1930 ) ? ( n36381 ) : ( n36385 ) ;
assign n36387 =  ( n879 ) ? ( n36376 ) : ( n36386 ) ;
assign n36388 =  ( n172 ) ? ( n32712 ) : ( VREG_12_8 ) ;
assign n36389 =  ( n170 ) ? ( n32711 ) : ( n36388 ) ;
assign n36390 =  ( n168 ) ? ( n32710 ) : ( n36389 ) ;
assign n36391 =  ( n166 ) ? ( n32709 ) : ( n36390 ) ;
assign n36392 =  ( n162 ) ? ( n32708 ) : ( n36391 ) ;
assign n36393 =  ( n172 ) ? ( n32722 ) : ( VREG_12_8 ) ;
assign n36394 =  ( n170 ) ? ( n32721 ) : ( n36393 ) ;
assign n36395 =  ( n168 ) ? ( n32720 ) : ( n36394 ) ;
assign n36396 =  ( n166 ) ? ( n32719 ) : ( n36395 ) ;
assign n36397 =  ( n162 ) ? ( n32718 ) : ( n36396 ) ;
assign n36398 =  ( n32701 ) ? ( VREG_12_8 ) : ( n36397 ) ;
assign n36399 =  ( n3051 ) ? ( n36398 ) : ( VREG_12_8 ) ;
assign n36400 =  ( n3040 ) ? ( n36392 ) : ( n36399 ) ;
assign n36401 =  ( n192 ) ? ( VREG_12_8 ) : ( VREG_12_8 ) ;
assign n36402 =  ( n157 ) ? ( n36400 ) : ( n36401 ) ;
assign n36403 =  ( n6 ) ? ( n36387 ) : ( n36402 ) ;
assign n36404 =  ( n263 ) ? ( n36403 ) : ( VREG_12_8 ) ;
assign n36405 =  ( n148 ) ? ( n33779 ) : ( VREG_12_9 ) ;
assign n36406 =  ( n146 ) ? ( n33778 ) : ( n36405 ) ;
assign n36407 =  ( n144 ) ? ( n33777 ) : ( n36406 ) ;
assign n36408 =  ( n142 ) ? ( n33776 ) : ( n36407 ) ;
assign n36409 =  ( n10 ) ? ( n33775 ) : ( n36408 ) ;
assign n36410 =  ( n148 ) ? ( n34813 ) : ( VREG_12_9 ) ;
assign n36411 =  ( n146 ) ? ( n34812 ) : ( n36410 ) ;
assign n36412 =  ( n144 ) ? ( n34811 ) : ( n36411 ) ;
assign n36413 =  ( n142 ) ? ( n34810 ) : ( n36412 ) ;
assign n36414 =  ( n10 ) ? ( n34809 ) : ( n36413 ) ;
assign n36415 =  ( n34820 ) ? ( VREG_12_9 ) : ( n36409 ) ;
assign n36416 =  ( n34820 ) ? ( VREG_12_9 ) : ( n36414 ) ;
assign n36417 =  ( n3034 ) ? ( n36416 ) : ( VREG_12_9 ) ;
assign n36418 =  ( n2965 ) ? ( n36415 ) : ( n36417 ) ;
assign n36419 =  ( n1930 ) ? ( n36414 ) : ( n36418 ) ;
assign n36420 =  ( n879 ) ? ( n36409 ) : ( n36419 ) ;
assign n36421 =  ( n172 ) ? ( n34831 ) : ( VREG_12_9 ) ;
assign n36422 =  ( n170 ) ? ( n34830 ) : ( n36421 ) ;
assign n36423 =  ( n168 ) ? ( n34829 ) : ( n36422 ) ;
assign n36424 =  ( n166 ) ? ( n34828 ) : ( n36423 ) ;
assign n36425 =  ( n162 ) ? ( n34827 ) : ( n36424 ) ;
assign n36426 =  ( n172 ) ? ( n34841 ) : ( VREG_12_9 ) ;
assign n36427 =  ( n170 ) ? ( n34840 ) : ( n36426 ) ;
assign n36428 =  ( n168 ) ? ( n34839 ) : ( n36427 ) ;
assign n36429 =  ( n166 ) ? ( n34838 ) : ( n36428 ) ;
assign n36430 =  ( n162 ) ? ( n34837 ) : ( n36429 ) ;
assign n36431 =  ( n34820 ) ? ( VREG_12_9 ) : ( n36430 ) ;
assign n36432 =  ( n3051 ) ? ( n36431 ) : ( VREG_12_9 ) ;
assign n36433 =  ( n3040 ) ? ( n36425 ) : ( n36432 ) ;
assign n36434 =  ( n192 ) ? ( VREG_12_9 ) : ( VREG_12_9 ) ;
assign n36435 =  ( n157 ) ? ( n36433 ) : ( n36434 ) ;
assign n36436 =  ( n6 ) ? ( n36420 ) : ( n36435 ) ;
assign n36437 =  ( n263 ) ? ( n36436 ) : ( VREG_12_9 ) ;
assign n36438 =  ( n148 ) ? ( n1924 ) : ( VREG_13_0 ) ;
assign n36439 =  ( n146 ) ? ( n1923 ) : ( n36438 ) ;
assign n36440 =  ( n144 ) ? ( n1922 ) : ( n36439 ) ;
assign n36441 =  ( n142 ) ? ( n1921 ) : ( n36440 ) ;
assign n36442 =  ( n10 ) ? ( n1920 ) : ( n36441 ) ;
assign n36443 =  ( n148 ) ? ( n2959 ) : ( VREG_13_0 ) ;
assign n36444 =  ( n146 ) ? ( n2958 ) : ( n36443 ) ;
assign n36445 =  ( n144 ) ? ( n2957 ) : ( n36444 ) ;
assign n36446 =  ( n142 ) ? ( n2956 ) : ( n36445 ) ;
assign n36447 =  ( n10 ) ? ( n2955 ) : ( n36446 ) ;
assign n36448 =  ( n3032 ) ? ( VREG_13_0 ) : ( n36442 ) ;
assign n36449 =  ( n3032 ) ? ( VREG_13_0 ) : ( n36447 ) ;
assign n36450 =  ( n3034 ) ? ( n36449 ) : ( VREG_13_0 ) ;
assign n36451 =  ( n2965 ) ? ( n36448 ) : ( n36450 ) ;
assign n36452 =  ( n1930 ) ? ( n36447 ) : ( n36451 ) ;
assign n36453 =  ( n879 ) ? ( n36442 ) : ( n36452 ) ;
assign n36454 =  ( n172 ) ? ( n3045 ) : ( VREG_13_0 ) ;
assign n36455 =  ( n170 ) ? ( n3044 ) : ( n36454 ) ;
assign n36456 =  ( n168 ) ? ( n3043 ) : ( n36455 ) ;
assign n36457 =  ( n166 ) ? ( n3042 ) : ( n36456 ) ;
assign n36458 =  ( n162 ) ? ( n3041 ) : ( n36457 ) ;
assign n36459 =  ( n172 ) ? ( n3056 ) : ( VREG_13_0 ) ;
assign n36460 =  ( n170 ) ? ( n3055 ) : ( n36459 ) ;
assign n36461 =  ( n168 ) ? ( n3054 ) : ( n36460 ) ;
assign n36462 =  ( n166 ) ? ( n3053 ) : ( n36461 ) ;
assign n36463 =  ( n162 ) ? ( n3052 ) : ( n36462 ) ;
assign n36464 =  ( n3032 ) ? ( VREG_13_0 ) : ( n36463 ) ;
assign n36465 =  ( n3051 ) ? ( n36464 ) : ( VREG_13_0 ) ;
assign n36466 =  ( n3040 ) ? ( n36458 ) : ( n36465 ) ;
assign n36467 =  ( n192 ) ? ( VREG_13_0 ) : ( VREG_13_0 ) ;
assign n36468 =  ( n157 ) ? ( n36466 ) : ( n36467 ) ;
assign n36469 =  ( n6 ) ? ( n36453 ) : ( n36468 ) ;
assign n36470 =  ( n285 ) ? ( n36469 ) : ( VREG_13_0 ) ;
assign n36471 =  ( n148 ) ? ( n4113 ) : ( VREG_13_1 ) ;
assign n36472 =  ( n146 ) ? ( n4112 ) : ( n36471 ) ;
assign n36473 =  ( n144 ) ? ( n4111 ) : ( n36472 ) ;
assign n36474 =  ( n142 ) ? ( n4110 ) : ( n36473 ) ;
assign n36475 =  ( n10 ) ? ( n4109 ) : ( n36474 ) ;
assign n36476 =  ( n148 ) ? ( n5147 ) : ( VREG_13_1 ) ;
assign n36477 =  ( n146 ) ? ( n5146 ) : ( n36476 ) ;
assign n36478 =  ( n144 ) ? ( n5145 ) : ( n36477 ) ;
assign n36479 =  ( n142 ) ? ( n5144 ) : ( n36478 ) ;
assign n36480 =  ( n10 ) ? ( n5143 ) : ( n36479 ) ;
assign n36481 =  ( n5154 ) ? ( VREG_13_1 ) : ( n36475 ) ;
assign n36482 =  ( n5154 ) ? ( VREG_13_1 ) : ( n36480 ) ;
assign n36483 =  ( n3034 ) ? ( n36482 ) : ( VREG_13_1 ) ;
assign n36484 =  ( n2965 ) ? ( n36481 ) : ( n36483 ) ;
assign n36485 =  ( n1930 ) ? ( n36480 ) : ( n36484 ) ;
assign n36486 =  ( n879 ) ? ( n36475 ) : ( n36485 ) ;
assign n36487 =  ( n172 ) ? ( n5165 ) : ( VREG_13_1 ) ;
assign n36488 =  ( n170 ) ? ( n5164 ) : ( n36487 ) ;
assign n36489 =  ( n168 ) ? ( n5163 ) : ( n36488 ) ;
assign n36490 =  ( n166 ) ? ( n5162 ) : ( n36489 ) ;
assign n36491 =  ( n162 ) ? ( n5161 ) : ( n36490 ) ;
assign n36492 =  ( n172 ) ? ( n5175 ) : ( VREG_13_1 ) ;
assign n36493 =  ( n170 ) ? ( n5174 ) : ( n36492 ) ;
assign n36494 =  ( n168 ) ? ( n5173 ) : ( n36493 ) ;
assign n36495 =  ( n166 ) ? ( n5172 ) : ( n36494 ) ;
assign n36496 =  ( n162 ) ? ( n5171 ) : ( n36495 ) ;
assign n36497 =  ( n5154 ) ? ( VREG_13_1 ) : ( n36496 ) ;
assign n36498 =  ( n3051 ) ? ( n36497 ) : ( VREG_13_1 ) ;
assign n36499 =  ( n3040 ) ? ( n36491 ) : ( n36498 ) ;
assign n36500 =  ( n192 ) ? ( VREG_13_1 ) : ( VREG_13_1 ) ;
assign n36501 =  ( n157 ) ? ( n36499 ) : ( n36500 ) ;
assign n36502 =  ( n6 ) ? ( n36486 ) : ( n36501 ) ;
assign n36503 =  ( n285 ) ? ( n36502 ) : ( VREG_13_1 ) ;
assign n36504 =  ( n148 ) ? ( n6232 ) : ( VREG_13_10 ) ;
assign n36505 =  ( n146 ) ? ( n6231 ) : ( n36504 ) ;
assign n36506 =  ( n144 ) ? ( n6230 ) : ( n36505 ) ;
assign n36507 =  ( n142 ) ? ( n6229 ) : ( n36506 ) ;
assign n36508 =  ( n10 ) ? ( n6228 ) : ( n36507 ) ;
assign n36509 =  ( n148 ) ? ( n7266 ) : ( VREG_13_10 ) ;
assign n36510 =  ( n146 ) ? ( n7265 ) : ( n36509 ) ;
assign n36511 =  ( n144 ) ? ( n7264 ) : ( n36510 ) ;
assign n36512 =  ( n142 ) ? ( n7263 ) : ( n36511 ) ;
assign n36513 =  ( n10 ) ? ( n7262 ) : ( n36512 ) ;
assign n36514 =  ( n7273 ) ? ( VREG_13_10 ) : ( n36508 ) ;
assign n36515 =  ( n7273 ) ? ( VREG_13_10 ) : ( n36513 ) ;
assign n36516 =  ( n3034 ) ? ( n36515 ) : ( VREG_13_10 ) ;
assign n36517 =  ( n2965 ) ? ( n36514 ) : ( n36516 ) ;
assign n36518 =  ( n1930 ) ? ( n36513 ) : ( n36517 ) ;
assign n36519 =  ( n879 ) ? ( n36508 ) : ( n36518 ) ;
assign n36520 =  ( n172 ) ? ( n7284 ) : ( VREG_13_10 ) ;
assign n36521 =  ( n170 ) ? ( n7283 ) : ( n36520 ) ;
assign n36522 =  ( n168 ) ? ( n7282 ) : ( n36521 ) ;
assign n36523 =  ( n166 ) ? ( n7281 ) : ( n36522 ) ;
assign n36524 =  ( n162 ) ? ( n7280 ) : ( n36523 ) ;
assign n36525 =  ( n172 ) ? ( n7294 ) : ( VREG_13_10 ) ;
assign n36526 =  ( n170 ) ? ( n7293 ) : ( n36525 ) ;
assign n36527 =  ( n168 ) ? ( n7292 ) : ( n36526 ) ;
assign n36528 =  ( n166 ) ? ( n7291 ) : ( n36527 ) ;
assign n36529 =  ( n162 ) ? ( n7290 ) : ( n36528 ) ;
assign n36530 =  ( n7273 ) ? ( VREG_13_10 ) : ( n36529 ) ;
assign n36531 =  ( n3051 ) ? ( n36530 ) : ( VREG_13_10 ) ;
assign n36532 =  ( n3040 ) ? ( n36524 ) : ( n36531 ) ;
assign n36533 =  ( n192 ) ? ( VREG_13_10 ) : ( VREG_13_10 ) ;
assign n36534 =  ( n157 ) ? ( n36532 ) : ( n36533 ) ;
assign n36535 =  ( n6 ) ? ( n36519 ) : ( n36534 ) ;
assign n36536 =  ( n285 ) ? ( n36535 ) : ( VREG_13_10 ) ;
assign n36537 =  ( n148 ) ? ( n8351 ) : ( VREG_13_11 ) ;
assign n36538 =  ( n146 ) ? ( n8350 ) : ( n36537 ) ;
assign n36539 =  ( n144 ) ? ( n8349 ) : ( n36538 ) ;
assign n36540 =  ( n142 ) ? ( n8348 ) : ( n36539 ) ;
assign n36541 =  ( n10 ) ? ( n8347 ) : ( n36540 ) ;
assign n36542 =  ( n148 ) ? ( n9385 ) : ( VREG_13_11 ) ;
assign n36543 =  ( n146 ) ? ( n9384 ) : ( n36542 ) ;
assign n36544 =  ( n144 ) ? ( n9383 ) : ( n36543 ) ;
assign n36545 =  ( n142 ) ? ( n9382 ) : ( n36544 ) ;
assign n36546 =  ( n10 ) ? ( n9381 ) : ( n36545 ) ;
assign n36547 =  ( n9392 ) ? ( VREG_13_11 ) : ( n36541 ) ;
assign n36548 =  ( n9392 ) ? ( VREG_13_11 ) : ( n36546 ) ;
assign n36549 =  ( n3034 ) ? ( n36548 ) : ( VREG_13_11 ) ;
assign n36550 =  ( n2965 ) ? ( n36547 ) : ( n36549 ) ;
assign n36551 =  ( n1930 ) ? ( n36546 ) : ( n36550 ) ;
assign n36552 =  ( n879 ) ? ( n36541 ) : ( n36551 ) ;
assign n36553 =  ( n172 ) ? ( n9403 ) : ( VREG_13_11 ) ;
assign n36554 =  ( n170 ) ? ( n9402 ) : ( n36553 ) ;
assign n36555 =  ( n168 ) ? ( n9401 ) : ( n36554 ) ;
assign n36556 =  ( n166 ) ? ( n9400 ) : ( n36555 ) ;
assign n36557 =  ( n162 ) ? ( n9399 ) : ( n36556 ) ;
assign n36558 =  ( n172 ) ? ( n9413 ) : ( VREG_13_11 ) ;
assign n36559 =  ( n170 ) ? ( n9412 ) : ( n36558 ) ;
assign n36560 =  ( n168 ) ? ( n9411 ) : ( n36559 ) ;
assign n36561 =  ( n166 ) ? ( n9410 ) : ( n36560 ) ;
assign n36562 =  ( n162 ) ? ( n9409 ) : ( n36561 ) ;
assign n36563 =  ( n9392 ) ? ( VREG_13_11 ) : ( n36562 ) ;
assign n36564 =  ( n3051 ) ? ( n36563 ) : ( VREG_13_11 ) ;
assign n36565 =  ( n3040 ) ? ( n36557 ) : ( n36564 ) ;
assign n36566 =  ( n192 ) ? ( VREG_13_11 ) : ( VREG_13_11 ) ;
assign n36567 =  ( n157 ) ? ( n36565 ) : ( n36566 ) ;
assign n36568 =  ( n6 ) ? ( n36552 ) : ( n36567 ) ;
assign n36569 =  ( n285 ) ? ( n36568 ) : ( VREG_13_11 ) ;
assign n36570 =  ( n148 ) ? ( n10470 ) : ( VREG_13_12 ) ;
assign n36571 =  ( n146 ) ? ( n10469 ) : ( n36570 ) ;
assign n36572 =  ( n144 ) ? ( n10468 ) : ( n36571 ) ;
assign n36573 =  ( n142 ) ? ( n10467 ) : ( n36572 ) ;
assign n36574 =  ( n10 ) ? ( n10466 ) : ( n36573 ) ;
assign n36575 =  ( n148 ) ? ( n11504 ) : ( VREG_13_12 ) ;
assign n36576 =  ( n146 ) ? ( n11503 ) : ( n36575 ) ;
assign n36577 =  ( n144 ) ? ( n11502 ) : ( n36576 ) ;
assign n36578 =  ( n142 ) ? ( n11501 ) : ( n36577 ) ;
assign n36579 =  ( n10 ) ? ( n11500 ) : ( n36578 ) ;
assign n36580 =  ( n11511 ) ? ( VREG_13_12 ) : ( n36574 ) ;
assign n36581 =  ( n11511 ) ? ( VREG_13_12 ) : ( n36579 ) ;
assign n36582 =  ( n3034 ) ? ( n36581 ) : ( VREG_13_12 ) ;
assign n36583 =  ( n2965 ) ? ( n36580 ) : ( n36582 ) ;
assign n36584 =  ( n1930 ) ? ( n36579 ) : ( n36583 ) ;
assign n36585 =  ( n879 ) ? ( n36574 ) : ( n36584 ) ;
assign n36586 =  ( n172 ) ? ( n11522 ) : ( VREG_13_12 ) ;
assign n36587 =  ( n170 ) ? ( n11521 ) : ( n36586 ) ;
assign n36588 =  ( n168 ) ? ( n11520 ) : ( n36587 ) ;
assign n36589 =  ( n166 ) ? ( n11519 ) : ( n36588 ) ;
assign n36590 =  ( n162 ) ? ( n11518 ) : ( n36589 ) ;
assign n36591 =  ( n172 ) ? ( n11532 ) : ( VREG_13_12 ) ;
assign n36592 =  ( n170 ) ? ( n11531 ) : ( n36591 ) ;
assign n36593 =  ( n168 ) ? ( n11530 ) : ( n36592 ) ;
assign n36594 =  ( n166 ) ? ( n11529 ) : ( n36593 ) ;
assign n36595 =  ( n162 ) ? ( n11528 ) : ( n36594 ) ;
assign n36596 =  ( n11511 ) ? ( VREG_13_12 ) : ( n36595 ) ;
assign n36597 =  ( n3051 ) ? ( n36596 ) : ( VREG_13_12 ) ;
assign n36598 =  ( n3040 ) ? ( n36590 ) : ( n36597 ) ;
assign n36599 =  ( n192 ) ? ( VREG_13_12 ) : ( VREG_13_12 ) ;
assign n36600 =  ( n157 ) ? ( n36598 ) : ( n36599 ) ;
assign n36601 =  ( n6 ) ? ( n36585 ) : ( n36600 ) ;
assign n36602 =  ( n285 ) ? ( n36601 ) : ( VREG_13_12 ) ;
assign n36603 =  ( n148 ) ? ( n12589 ) : ( VREG_13_13 ) ;
assign n36604 =  ( n146 ) ? ( n12588 ) : ( n36603 ) ;
assign n36605 =  ( n144 ) ? ( n12587 ) : ( n36604 ) ;
assign n36606 =  ( n142 ) ? ( n12586 ) : ( n36605 ) ;
assign n36607 =  ( n10 ) ? ( n12585 ) : ( n36606 ) ;
assign n36608 =  ( n148 ) ? ( n13623 ) : ( VREG_13_13 ) ;
assign n36609 =  ( n146 ) ? ( n13622 ) : ( n36608 ) ;
assign n36610 =  ( n144 ) ? ( n13621 ) : ( n36609 ) ;
assign n36611 =  ( n142 ) ? ( n13620 ) : ( n36610 ) ;
assign n36612 =  ( n10 ) ? ( n13619 ) : ( n36611 ) ;
assign n36613 =  ( n13630 ) ? ( VREG_13_13 ) : ( n36607 ) ;
assign n36614 =  ( n13630 ) ? ( VREG_13_13 ) : ( n36612 ) ;
assign n36615 =  ( n3034 ) ? ( n36614 ) : ( VREG_13_13 ) ;
assign n36616 =  ( n2965 ) ? ( n36613 ) : ( n36615 ) ;
assign n36617 =  ( n1930 ) ? ( n36612 ) : ( n36616 ) ;
assign n36618 =  ( n879 ) ? ( n36607 ) : ( n36617 ) ;
assign n36619 =  ( n172 ) ? ( n13641 ) : ( VREG_13_13 ) ;
assign n36620 =  ( n170 ) ? ( n13640 ) : ( n36619 ) ;
assign n36621 =  ( n168 ) ? ( n13639 ) : ( n36620 ) ;
assign n36622 =  ( n166 ) ? ( n13638 ) : ( n36621 ) ;
assign n36623 =  ( n162 ) ? ( n13637 ) : ( n36622 ) ;
assign n36624 =  ( n172 ) ? ( n13651 ) : ( VREG_13_13 ) ;
assign n36625 =  ( n170 ) ? ( n13650 ) : ( n36624 ) ;
assign n36626 =  ( n168 ) ? ( n13649 ) : ( n36625 ) ;
assign n36627 =  ( n166 ) ? ( n13648 ) : ( n36626 ) ;
assign n36628 =  ( n162 ) ? ( n13647 ) : ( n36627 ) ;
assign n36629 =  ( n13630 ) ? ( VREG_13_13 ) : ( n36628 ) ;
assign n36630 =  ( n3051 ) ? ( n36629 ) : ( VREG_13_13 ) ;
assign n36631 =  ( n3040 ) ? ( n36623 ) : ( n36630 ) ;
assign n36632 =  ( n192 ) ? ( VREG_13_13 ) : ( VREG_13_13 ) ;
assign n36633 =  ( n157 ) ? ( n36631 ) : ( n36632 ) ;
assign n36634 =  ( n6 ) ? ( n36618 ) : ( n36633 ) ;
assign n36635 =  ( n285 ) ? ( n36634 ) : ( VREG_13_13 ) ;
assign n36636 =  ( n148 ) ? ( n14708 ) : ( VREG_13_14 ) ;
assign n36637 =  ( n146 ) ? ( n14707 ) : ( n36636 ) ;
assign n36638 =  ( n144 ) ? ( n14706 ) : ( n36637 ) ;
assign n36639 =  ( n142 ) ? ( n14705 ) : ( n36638 ) ;
assign n36640 =  ( n10 ) ? ( n14704 ) : ( n36639 ) ;
assign n36641 =  ( n148 ) ? ( n15742 ) : ( VREG_13_14 ) ;
assign n36642 =  ( n146 ) ? ( n15741 ) : ( n36641 ) ;
assign n36643 =  ( n144 ) ? ( n15740 ) : ( n36642 ) ;
assign n36644 =  ( n142 ) ? ( n15739 ) : ( n36643 ) ;
assign n36645 =  ( n10 ) ? ( n15738 ) : ( n36644 ) ;
assign n36646 =  ( n15749 ) ? ( VREG_13_14 ) : ( n36640 ) ;
assign n36647 =  ( n15749 ) ? ( VREG_13_14 ) : ( n36645 ) ;
assign n36648 =  ( n3034 ) ? ( n36647 ) : ( VREG_13_14 ) ;
assign n36649 =  ( n2965 ) ? ( n36646 ) : ( n36648 ) ;
assign n36650 =  ( n1930 ) ? ( n36645 ) : ( n36649 ) ;
assign n36651 =  ( n879 ) ? ( n36640 ) : ( n36650 ) ;
assign n36652 =  ( n172 ) ? ( n15760 ) : ( VREG_13_14 ) ;
assign n36653 =  ( n170 ) ? ( n15759 ) : ( n36652 ) ;
assign n36654 =  ( n168 ) ? ( n15758 ) : ( n36653 ) ;
assign n36655 =  ( n166 ) ? ( n15757 ) : ( n36654 ) ;
assign n36656 =  ( n162 ) ? ( n15756 ) : ( n36655 ) ;
assign n36657 =  ( n172 ) ? ( n15770 ) : ( VREG_13_14 ) ;
assign n36658 =  ( n170 ) ? ( n15769 ) : ( n36657 ) ;
assign n36659 =  ( n168 ) ? ( n15768 ) : ( n36658 ) ;
assign n36660 =  ( n166 ) ? ( n15767 ) : ( n36659 ) ;
assign n36661 =  ( n162 ) ? ( n15766 ) : ( n36660 ) ;
assign n36662 =  ( n15749 ) ? ( VREG_13_14 ) : ( n36661 ) ;
assign n36663 =  ( n3051 ) ? ( n36662 ) : ( VREG_13_14 ) ;
assign n36664 =  ( n3040 ) ? ( n36656 ) : ( n36663 ) ;
assign n36665 =  ( n192 ) ? ( VREG_13_14 ) : ( VREG_13_14 ) ;
assign n36666 =  ( n157 ) ? ( n36664 ) : ( n36665 ) ;
assign n36667 =  ( n6 ) ? ( n36651 ) : ( n36666 ) ;
assign n36668 =  ( n285 ) ? ( n36667 ) : ( VREG_13_14 ) ;
assign n36669 =  ( n148 ) ? ( n16827 ) : ( VREG_13_15 ) ;
assign n36670 =  ( n146 ) ? ( n16826 ) : ( n36669 ) ;
assign n36671 =  ( n144 ) ? ( n16825 ) : ( n36670 ) ;
assign n36672 =  ( n142 ) ? ( n16824 ) : ( n36671 ) ;
assign n36673 =  ( n10 ) ? ( n16823 ) : ( n36672 ) ;
assign n36674 =  ( n148 ) ? ( n17861 ) : ( VREG_13_15 ) ;
assign n36675 =  ( n146 ) ? ( n17860 ) : ( n36674 ) ;
assign n36676 =  ( n144 ) ? ( n17859 ) : ( n36675 ) ;
assign n36677 =  ( n142 ) ? ( n17858 ) : ( n36676 ) ;
assign n36678 =  ( n10 ) ? ( n17857 ) : ( n36677 ) ;
assign n36679 =  ( n17868 ) ? ( VREG_13_15 ) : ( n36673 ) ;
assign n36680 =  ( n17868 ) ? ( VREG_13_15 ) : ( n36678 ) ;
assign n36681 =  ( n3034 ) ? ( n36680 ) : ( VREG_13_15 ) ;
assign n36682 =  ( n2965 ) ? ( n36679 ) : ( n36681 ) ;
assign n36683 =  ( n1930 ) ? ( n36678 ) : ( n36682 ) ;
assign n36684 =  ( n879 ) ? ( n36673 ) : ( n36683 ) ;
assign n36685 =  ( n172 ) ? ( n17879 ) : ( VREG_13_15 ) ;
assign n36686 =  ( n170 ) ? ( n17878 ) : ( n36685 ) ;
assign n36687 =  ( n168 ) ? ( n17877 ) : ( n36686 ) ;
assign n36688 =  ( n166 ) ? ( n17876 ) : ( n36687 ) ;
assign n36689 =  ( n162 ) ? ( n17875 ) : ( n36688 ) ;
assign n36690 =  ( n172 ) ? ( n17889 ) : ( VREG_13_15 ) ;
assign n36691 =  ( n170 ) ? ( n17888 ) : ( n36690 ) ;
assign n36692 =  ( n168 ) ? ( n17887 ) : ( n36691 ) ;
assign n36693 =  ( n166 ) ? ( n17886 ) : ( n36692 ) ;
assign n36694 =  ( n162 ) ? ( n17885 ) : ( n36693 ) ;
assign n36695 =  ( n17868 ) ? ( VREG_13_15 ) : ( n36694 ) ;
assign n36696 =  ( n3051 ) ? ( n36695 ) : ( VREG_13_15 ) ;
assign n36697 =  ( n3040 ) ? ( n36689 ) : ( n36696 ) ;
assign n36698 =  ( n192 ) ? ( VREG_13_15 ) : ( VREG_13_15 ) ;
assign n36699 =  ( n157 ) ? ( n36697 ) : ( n36698 ) ;
assign n36700 =  ( n6 ) ? ( n36684 ) : ( n36699 ) ;
assign n36701 =  ( n285 ) ? ( n36700 ) : ( VREG_13_15 ) ;
assign n36702 =  ( n148 ) ? ( n18946 ) : ( VREG_13_2 ) ;
assign n36703 =  ( n146 ) ? ( n18945 ) : ( n36702 ) ;
assign n36704 =  ( n144 ) ? ( n18944 ) : ( n36703 ) ;
assign n36705 =  ( n142 ) ? ( n18943 ) : ( n36704 ) ;
assign n36706 =  ( n10 ) ? ( n18942 ) : ( n36705 ) ;
assign n36707 =  ( n148 ) ? ( n19980 ) : ( VREG_13_2 ) ;
assign n36708 =  ( n146 ) ? ( n19979 ) : ( n36707 ) ;
assign n36709 =  ( n144 ) ? ( n19978 ) : ( n36708 ) ;
assign n36710 =  ( n142 ) ? ( n19977 ) : ( n36709 ) ;
assign n36711 =  ( n10 ) ? ( n19976 ) : ( n36710 ) ;
assign n36712 =  ( n19987 ) ? ( VREG_13_2 ) : ( n36706 ) ;
assign n36713 =  ( n19987 ) ? ( VREG_13_2 ) : ( n36711 ) ;
assign n36714 =  ( n3034 ) ? ( n36713 ) : ( VREG_13_2 ) ;
assign n36715 =  ( n2965 ) ? ( n36712 ) : ( n36714 ) ;
assign n36716 =  ( n1930 ) ? ( n36711 ) : ( n36715 ) ;
assign n36717 =  ( n879 ) ? ( n36706 ) : ( n36716 ) ;
assign n36718 =  ( n172 ) ? ( n19998 ) : ( VREG_13_2 ) ;
assign n36719 =  ( n170 ) ? ( n19997 ) : ( n36718 ) ;
assign n36720 =  ( n168 ) ? ( n19996 ) : ( n36719 ) ;
assign n36721 =  ( n166 ) ? ( n19995 ) : ( n36720 ) ;
assign n36722 =  ( n162 ) ? ( n19994 ) : ( n36721 ) ;
assign n36723 =  ( n172 ) ? ( n20008 ) : ( VREG_13_2 ) ;
assign n36724 =  ( n170 ) ? ( n20007 ) : ( n36723 ) ;
assign n36725 =  ( n168 ) ? ( n20006 ) : ( n36724 ) ;
assign n36726 =  ( n166 ) ? ( n20005 ) : ( n36725 ) ;
assign n36727 =  ( n162 ) ? ( n20004 ) : ( n36726 ) ;
assign n36728 =  ( n19987 ) ? ( VREG_13_2 ) : ( n36727 ) ;
assign n36729 =  ( n3051 ) ? ( n36728 ) : ( VREG_13_2 ) ;
assign n36730 =  ( n3040 ) ? ( n36722 ) : ( n36729 ) ;
assign n36731 =  ( n192 ) ? ( VREG_13_2 ) : ( VREG_13_2 ) ;
assign n36732 =  ( n157 ) ? ( n36730 ) : ( n36731 ) ;
assign n36733 =  ( n6 ) ? ( n36717 ) : ( n36732 ) ;
assign n36734 =  ( n285 ) ? ( n36733 ) : ( VREG_13_2 ) ;
assign n36735 =  ( n148 ) ? ( n21065 ) : ( VREG_13_3 ) ;
assign n36736 =  ( n146 ) ? ( n21064 ) : ( n36735 ) ;
assign n36737 =  ( n144 ) ? ( n21063 ) : ( n36736 ) ;
assign n36738 =  ( n142 ) ? ( n21062 ) : ( n36737 ) ;
assign n36739 =  ( n10 ) ? ( n21061 ) : ( n36738 ) ;
assign n36740 =  ( n148 ) ? ( n22099 ) : ( VREG_13_3 ) ;
assign n36741 =  ( n146 ) ? ( n22098 ) : ( n36740 ) ;
assign n36742 =  ( n144 ) ? ( n22097 ) : ( n36741 ) ;
assign n36743 =  ( n142 ) ? ( n22096 ) : ( n36742 ) ;
assign n36744 =  ( n10 ) ? ( n22095 ) : ( n36743 ) ;
assign n36745 =  ( n22106 ) ? ( VREG_13_3 ) : ( n36739 ) ;
assign n36746 =  ( n22106 ) ? ( VREG_13_3 ) : ( n36744 ) ;
assign n36747 =  ( n3034 ) ? ( n36746 ) : ( VREG_13_3 ) ;
assign n36748 =  ( n2965 ) ? ( n36745 ) : ( n36747 ) ;
assign n36749 =  ( n1930 ) ? ( n36744 ) : ( n36748 ) ;
assign n36750 =  ( n879 ) ? ( n36739 ) : ( n36749 ) ;
assign n36751 =  ( n172 ) ? ( n22117 ) : ( VREG_13_3 ) ;
assign n36752 =  ( n170 ) ? ( n22116 ) : ( n36751 ) ;
assign n36753 =  ( n168 ) ? ( n22115 ) : ( n36752 ) ;
assign n36754 =  ( n166 ) ? ( n22114 ) : ( n36753 ) ;
assign n36755 =  ( n162 ) ? ( n22113 ) : ( n36754 ) ;
assign n36756 =  ( n172 ) ? ( n22127 ) : ( VREG_13_3 ) ;
assign n36757 =  ( n170 ) ? ( n22126 ) : ( n36756 ) ;
assign n36758 =  ( n168 ) ? ( n22125 ) : ( n36757 ) ;
assign n36759 =  ( n166 ) ? ( n22124 ) : ( n36758 ) ;
assign n36760 =  ( n162 ) ? ( n22123 ) : ( n36759 ) ;
assign n36761 =  ( n22106 ) ? ( VREG_13_3 ) : ( n36760 ) ;
assign n36762 =  ( n3051 ) ? ( n36761 ) : ( VREG_13_3 ) ;
assign n36763 =  ( n3040 ) ? ( n36755 ) : ( n36762 ) ;
assign n36764 =  ( n192 ) ? ( VREG_13_3 ) : ( VREG_13_3 ) ;
assign n36765 =  ( n157 ) ? ( n36763 ) : ( n36764 ) ;
assign n36766 =  ( n6 ) ? ( n36750 ) : ( n36765 ) ;
assign n36767 =  ( n285 ) ? ( n36766 ) : ( VREG_13_3 ) ;
assign n36768 =  ( n148 ) ? ( n23184 ) : ( VREG_13_4 ) ;
assign n36769 =  ( n146 ) ? ( n23183 ) : ( n36768 ) ;
assign n36770 =  ( n144 ) ? ( n23182 ) : ( n36769 ) ;
assign n36771 =  ( n142 ) ? ( n23181 ) : ( n36770 ) ;
assign n36772 =  ( n10 ) ? ( n23180 ) : ( n36771 ) ;
assign n36773 =  ( n148 ) ? ( n24218 ) : ( VREG_13_4 ) ;
assign n36774 =  ( n146 ) ? ( n24217 ) : ( n36773 ) ;
assign n36775 =  ( n144 ) ? ( n24216 ) : ( n36774 ) ;
assign n36776 =  ( n142 ) ? ( n24215 ) : ( n36775 ) ;
assign n36777 =  ( n10 ) ? ( n24214 ) : ( n36776 ) ;
assign n36778 =  ( n24225 ) ? ( VREG_13_4 ) : ( n36772 ) ;
assign n36779 =  ( n24225 ) ? ( VREG_13_4 ) : ( n36777 ) ;
assign n36780 =  ( n3034 ) ? ( n36779 ) : ( VREG_13_4 ) ;
assign n36781 =  ( n2965 ) ? ( n36778 ) : ( n36780 ) ;
assign n36782 =  ( n1930 ) ? ( n36777 ) : ( n36781 ) ;
assign n36783 =  ( n879 ) ? ( n36772 ) : ( n36782 ) ;
assign n36784 =  ( n172 ) ? ( n24236 ) : ( VREG_13_4 ) ;
assign n36785 =  ( n170 ) ? ( n24235 ) : ( n36784 ) ;
assign n36786 =  ( n168 ) ? ( n24234 ) : ( n36785 ) ;
assign n36787 =  ( n166 ) ? ( n24233 ) : ( n36786 ) ;
assign n36788 =  ( n162 ) ? ( n24232 ) : ( n36787 ) ;
assign n36789 =  ( n172 ) ? ( n24246 ) : ( VREG_13_4 ) ;
assign n36790 =  ( n170 ) ? ( n24245 ) : ( n36789 ) ;
assign n36791 =  ( n168 ) ? ( n24244 ) : ( n36790 ) ;
assign n36792 =  ( n166 ) ? ( n24243 ) : ( n36791 ) ;
assign n36793 =  ( n162 ) ? ( n24242 ) : ( n36792 ) ;
assign n36794 =  ( n24225 ) ? ( VREG_13_4 ) : ( n36793 ) ;
assign n36795 =  ( n3051 ) ? ( n36794 ) : ( VREG_13_4 ) ;
assign n36796 =  ( n3040 ) ? ( n36788 ) : ( n36795 ) ;
assign n36797 =  ( n192 ) ? ( VREG_13_4 ) : ( VREG_13_4 ) ;
assign n36798 =  ( n157 ) ? ( n36796 ) : ( n36797 ) ;
assign n36799 =  ( n6 ) ? ( n36783 ) : ( n36798 ) ;
assign n36800 =  ( n285 ) ? ( n36799 ) : ( VREG_13_4 ) ;
assign n36801 =  ( n148 ) ? ( n25303 ) : ( VREG_13_5 ) ;
assign n36802 =  ( n146 ) ? ( n25302 ) : ( n36801 ) ;
assign n36803 =  ( n144 ) ? ( n25301 ) : ( n36802 ) ;
assign n36804 =  ( n142 ) ? ( n25300 ) : ( n36803 ) ;
assign n36805 =  ( n10 ) ? ( n25299 ) : ( n36804 ) ;
assign n36806 =  ( n148 ) ? ( n26337 ) : ( VREG_13_5 ) ;
assign n36807 =  ( n146 ) ? ( n26336 ) : ( n36806 ) ;
assign n36808 =  ( n144 ) ? ( n26335 ) : ( n36807 ) ;
assign n36809 =  ( n142 ) ? ( n26334 ) : ( n36808 ) ;
assign n36810 =  ( n10 ) ? ( n26333 ) : ( n36809 ) ;
assign n36811 =  ( n26344 ) ? ( VREG_13_5 ) : ( n36805 ) ;
assign n36812 =  ( n26344 ) ? ( VREG_13_5 ) : ( n36810 ) ;
assign n36813 =  ( n3034 ) ? ( n36812 ) : ( VREG_13_5 ) ;
assign n36814 =  ( n2965 ) ? ( n36811 ) : ( n36813 ) ;
assign n36815 =  ( n1930 ) ? ( n36810 ) : ( n36814 ) ;
assign n36816 =  ( n879 ) ? ( n36805 ) : ( n36815 ) ;
assign n36817 =  ( n172 ) ? ( n26355 ) : ( VREG_13_5 ) ;
assign n36818 =  ( n170 ) ? ( n26354 ) : ( n36817 ) ;
assign n36819 =  ( n168 ) ? ( n26353 ) : ( n36818 ) ;
assign n36820 =  ( n166 ) ? ( n26352 ) : ( n36819 ) ;
assign n36821 =  ( n162 ) ? ( n26351 ) : ( n36820 ) ;
assign n36822 =  ( n172 ) ? ( n26365 ) : ( VREG_13_5 ) ;
assign n36823 =  ( n170 ) ? ( n26364 ) : ( n36822 ) ;
assign n36824 =  ( n168 ) ? ( n26363 ) : ( n36823 ) ;
assign n36825 =  ( n166 ) ? ( n26362 ) : ( n36824 ) ;
assign n36826 =  ( n162 ) ? ( n26361 ) : ( n36825 ) ;
assign n36827 =  ( n26344 ) ? ( VREG_13_5 ) : ( n36826 ) ;
assign n36828 =  ( n3051 ) ? ( n36827 ) : ( VREG_13_5 ) ;
assign n36829 =  ( n3040 ) ? ( n36821 ) : ( n36828 ) ;
assign n36830 =  ( n192 ) ? ( VREG_13_5 ) : ( VREG_13_5 ) ;
assign n36831 =  ( n157 ) ? ( n36829 ) : ( n36830 ) ;
assign n36832 =  ( n6 ) ? ( n36816 ) : ( n36831 ) ;
assign n36833 =  ( n285 ) ? ( n36832 ) : ( VREG_13_5 ) ;
assign n36834 =  ( n148 ) ? ( n27422 ) : ( VREG_13_6 ) ;
assign n36835 =  ( n146 ) ? ( n27421 ) : ( n36834 ) ;
assign n36836 =  ( n144 ) ? ( n27420 ) : ( n36835 ) ;
assign n36837 =  ( n142 ) ? ( n27419 ) : ( n36836 ) ;
assign n36838 =  ( n10 ) ? ( n27418 ) : ( n36837 ) ;
assign n36839 =  ( n148 ) ? ( n28456 ) : ( VREG_13_6 ) ;
assign n36840 =  ( n146 ) ? ( n28455 ) : ( n36839 ) ;
assign n36841 =  ( n144 ) ? ( n28454 ) : ( n36840 ) ;
assign n36842 =  ( n142 ) ? ( n28453 ) : ( n36841 ) ;
assign n36843 =  ( n10 ) ? ( n28452 ) : ( n36842 ) ;
assign n36844 =  ( n28463 ) ? ( VREG_13_6 ) : ( n36838 ) ;
assign n36845 =  ( n28463 ) ? ( VREG_13_6 ) : ( n36843 ) ;
assign n36846 =  ( n3034 ) ? ( n36845 ) : ( VREG_13_6 ) ;
assign n36847 =  ( n2965 ) ? ( n36844 ) : ( n36846 ) ;
assign n36848 =  ( n1930 ) ? ( n36843 ) : ( n36847 ) ;
assign n36849 =  ( n879 ) ? ( n36838 ) : ( n36848 ) ;
assign n36850 =  ( n172 ) ? ( n28474 ) : ( VREG_13_6 ) ;
assign n36851 =  ( n170 ) ? ( n28473 ) : ( n36850 ) ;
assign n36852 =  ( n168 ) ? ( n28472 ) : ( n36851 ) ;
assign n36853 =  ( n166 ) ? ( n28471 ) : ( n36852 ) ;
assign n36854 =  ( n162 ) ? ( n28470 ) : ( n36853 ) ;
assign n36855 =  ( n172 ) ? ( n28484 ) : ( VREG_13_6 ) ;
assign n36856 =  ( n170 ) ? ( n28483 ) : ( n36855 ) ;
assign n36857 =  ( n168 ) ? ( n28482 ) : ( n36856 ) ;
assign n36858 =  ( n166 ) ? ( n28481 ) : ( n36857 ) ;
assign n36859 =  ( n162 ) ? ( n28480 ) : ( n36858 ) ;
assign n36860 =  ( n28463 ) ? ( VREG_13_6 ) : ( n36859 ) ;
assign n36861 =  ( n3051 ) ? ( n36860 ) : ( VREG_13_6 ) ;
assign n36862 =  ( n3040 ) ? ( n36854 ) : ( n36861 ) ;
assign n36863 =  ( n192 ) ? ( VREG_13_6 ) : ( VREG_13_6 ) ;
assign n36864 =  ( n157 ) ? ( n36862 ) : ( n36863 ) ;
assign n36865 =  ( n6 ) ? ( n36849 ) : ( n36864 ) ;
assign n36866 =  ( n285 ) ? ( n36865 ) : ( VREG_13_6 ) ;
assign n36867 =  ( n148 ) ? ( n29541 ) : ( VREG_13_7 ) ;
assign n36868 =  ( n146 ) ? ( n29540 ) : ( n36867 ) ;
assign n36869 =  ( n144 ) ? ( n29539 ) : ( n36868 ) ;
assign n36870 =  ( n142 ) ? ( n29538 ) : ( n36869 ) ;
assign n36871 =  ( n10 ) ? ( n29537 ) : ( n36870 ) ;
assign n36872 =  ( n148 ) ? ( n30575 ) : ( VREG_13_7 ) ;
assign n36873 =  ( n146 ) ? ( n30574 ) : ( n36872 ) ;
assign n36874 =  ( n144 ) ? ( n30573 ) : ( n36873 ) ;
assign n36875 =  ( n142 ) ? ( n30572 ) : ( n36874 ) ;
assign n36876 =  ( n10 ) ? ( n30571 ) : ( n36875 ) ;
assign n36877 =  ( n30582 ) ? ( VREG_13_7 ) : ( n36871 ) ;
assign n36878 =  ( n30582 ) ? ( VREG_13_7 ) : ( n36876 ) ;
assign n36879 =  ( n3034 ) ? ( n36878 ) : ( VREG_13_7 ) ;
assign n36880 =  ( n2965 ) ? ( n36877 ) : ( n36879 ) ;
assign n36881 =  ( n1930 ) ? ( n36876 ) : ( n36880 ) ;
assign n36882 =  ( n879 ) ? ( n36871 ) : ( n36881 ) ;
assign n36883 =  ( n172 ) ? ( n30593 ) : ( VREG_13_7 ) ;
assign n36884 =  ( n170 ) ? ( n30592 ) : ( n36883 ) ;
assign n36885 =  ( n168 ) ? ( n30591 ) : ( n36884 ) ;
assign n36886 =  ( n166 ) ? ( n30590 ) : ( n36885 ) ;
assign n36887 =  ( n162 ) ? ( n30589 ) : ( n36886 ) ;
assign n36888 =  ( n172 ) ? ( n30603 ) : ( VREG_13_7 ) ;
assign n36889 =  ( n170 ) ? ( n30602 ) : ( n36888 ) ;
assign n36890 =  ( n168 ) ? ( n30601 ) : ( n36889 ) ;
assign n36891 =  ( n166 ) ? ( n30600 ) : ( n36890 ) ;
assign n36892 =  ( n162 ) ? ( n30599 ) : ( n36891 ) ;
assign n36893 =  ( n30582 ) ? ( VREG_13_7 ) : ( n36892 ) ;
assign n36894 =  ( n3051 ) ? ( n36893 ) : ( VREG_13_7 ) ;
assign n36895 =  ( n3040 ) ? ( n36887 ) : ( n36894 ) ;
assign n36896 =  ( n192 ) ? ( VREG_13_7 ) : ( VREG_13_7 ) ;
assign n36897 =  ( n157 ) ? ( n36895 ) : ( n36896 ) ;
assign n36898 =  ( n6 ) ? ( n36882 ) : ( n36897 ) ;
assign n36899 =  ( n285 ) ? ( n36898 ) : ( VREG_13_7 ) ;
assign n36900 =  ( n148 ) ? ( n31660 ) : ( VREG_13_8 ) ;
assign n36901 =  ( n146 ) ? ( n31659 ) : ( n36900 ) ;
assign n36902 =  ( n144 ) ? ( n31658 ) : ( n36901 ) ;
assign n36903 =  ( n142 ) ? ( n31657 ) : ( n36902 ) ;
assign n36904 =  ( n10 ) ? ( n31656 ) : ( n36903 ) ;
assign n36905 =  ( n148 ) ? ( n32694 ) : ( VREG_13_8 ) ;
assign n36906 =  ( n146 ) ? ( n32693 ) : ( n36905 ) ;
assign n36907 =  ( n144 ) ? ( n32692 ) : ( n36906 ) ;
assign n36908 =  ( n142 ) ? ( n32691 ) : ( n36907 ) ;
assign n36909 =  ( n10 ) ? ( n32690 ) : ( n36908 ) ;
assign n36910 =  ( n32701 ) ? ( VREG_13_8 ) : ( n36904 ) ;
assign n36911 =  ( n32701 ) ? ( VREG_13_8 ) : ( n36909 ) ;
assign n36912 =  ( n3034 ) ? ( n36911 ) : ( VREG_13_8 ) ;
assign n36913 =  ( n2965 ) ? ( n36910 ) : ( n36912 ) ;
assign n36914 =  ( n1930 ) ? ( n36909 ) : ( n36913 ) ;
assign n36915 =  ( n879 ) ? ( n36904 ) : ( n36914 ) ;
assign n36916 =  ( n172 ) ? ( n32712 ) : ( VREG_13_8 ) ;
assign n36917 =  ( n170 ) ? ( n32711 ) : ( n36916 ) ;
assign n36918 =  ( n168 ) ? ( n32710 ) : ( n36917 ) ;
assign n36919 =  ( n166 ) ? ( n32709 ) : ( n36918 ) ;
assign n36920 =  ( n162 ) ? ( n32708 ) : ( n36919 ) ;
assign n36921 =  ( n172 ) ? ( n32722 ) : ( VREG_13_8 ) ;
assign n36922 =  ( n170 ) ? ( n32721 ) : ( n36921 ) ;
assign n36923 =  ( n168 ) ? ( n32720 ) : ( n36922 ) ;
assign n36924 =  ( n166 ) ? ( n32719 ) : ( n36923 ) ;
assign n36925 =  ( n162 ) ? ( n32718 ) : ( n36924 ) ;
assign n36926 =  ( n32701 ) ? ( VREG_13_8 ) : ( n36925 ) ;
assign n36927 =  ( n3051 ) ? ( n36926 ) : ( VREG_13_8 ) ;
assign n36928 =  ( n3040 ) ? ( n36920 ) : ( n36927 ) ;
assign n36929 =  ( n192 ) ? ( VREG_13_8 ) : ( VREG_13_8 ) ;
assign n36930 =  ( n157 ) ? ( n36928 ) : ( n36929 ) ;
assign n36931 =  ( n6 ) ? ( n36915 ) : ( n36930 ) ;
assign n36932 =  ( n285 ) ? ( n36931 ) : ( VREG_13_8 ) ;
assign n36933 =  ( n148 ) ? ( n33779 ) : ( VREG_13_9 ) ;
assign n36934 =  ( n146 ) ? ( n33778 ) : ( n36933 ) ;
assign n36935 =  ( n144 ) ? ( n33777 ) : ( n36934 ) ;
assign n36936 =  ( n142 ) ? ( n33776 ) : ( n36935 ) ;
assign n36937 =  ( n10 ) ? ( n33775 ) : ( n36936 ) ;
assign n36938 =  ( n148 ) ? ( n34813 ) : ( VREG_13_9 ) ;
assign n36939 =  ( n146 ) ? ( n34812 ) : ( n36938 ) ;
assign n36940 =  ( n144 ) ? ( n34811 ) : ( n36939 ) ;
assign n36941 =  ( n142 ) ? ( n34810 ) : ( n36940 ) ;
assign n36942 =  ( n10 ) ? ( n34809 ) : ( n36941 ) ;
assign n36943 =  ( n34820 ) ? ( VREG_13_9 ) : ( n36937 ) ;
assign n36944 =  ( n34820 ) ? ( VREG_13_9 ) : ( n36942 ) ;
assign n36945 =  ( n3034 ) ? ( n36944 ) : ( VREG_13_9 ) ;
assign n36946 =  ( n2965 ) ? ( n36943 ) : ( n36945 ) ;
assign n36947 =  ( n1930 ) ? ( n36942 ) : ( n36946 ) ;
assign n36948 =  ( n879 ) ? ( n36937 ) : ( n36947 ) ;
assign n36949 =  ( n172 ) ? ( n34831 ) : ( VREG_13_9 ) ;
assign n36950 =  ( n170 ) ? ( n34830 ) : ( n36949 ) ;
assign n36951 =  ( n168 ) ? ( n34829 ) : ( n36950 ) ;
assign n36952 =  ( n166 ) ? ( n34828 ) : ( n36951 ) ;
assign n36953 =  ( n162 ) ? ( n34827 ) : ( n36952 ) ;
assign n36954 =  ( n172 ) ? ( n34841 ) : ( VREG_13_9 ) ;
assign n36955 =  ( n170 ) ? ( n34840 ) : ( n36954 ) ;
assign n36956 =  ( n168 ) ? ( n34839 ) : ( n36955 ) ;
assign n36957 =  ( n166 ) ? ( n34838 ) : ( n36956 ) ;
assign n36958 =  ( n162 ) ? ( n34837 ) : ( n36957 ) ;
assign n36959 =  ( n34820 ) ? ( VREG_13_9 ) : ( n36958 ) ;
assign n36960 =  ( n3051 ) ? ( n36959 ) : ( VREG_13_9 ) ;
assign n36961 =  ( n3040 ) ? ( n36953 ) : ( n36960 ) ;
assign n36962 =  ( n192 ) ? ( VREG_13_9 ) : ( VREG_13_9 ) ;
assign n36963 =  ( n157 ) ? ( n36961 ) : ( n36962 ) ;
assign n36964 =  ( n6 ) ? ( n36948 ) : ( n36963 ) ;
assign n36965 =  ( n285 ) ? ( n36964 ) : ( VREG_13_9 ) ;
assign n36966 =  ( n148 ) ? ( n1924 ) : ( VREG_14_0 ) ;
assign n36967 =  ( n146 ) ? ( n1923 ) : ( n36966 ) ;
assign n36968 =  ( n144 ) ? ( n1922 ) : ( n36967 ) ;
assign n36969 =  ( n142 ) ? ( n1921 ) : ( n36968 ) ;
assign n36970 =  ( n10 ) ? ( n1920 ) : ( n36969 ) ;
assign n36971 =  ( n148 ) ? ( n2959 ) : ( VREG_14_0 ) ;
assign n36972 =  ( n146 ) ? ( n2958 ) : ( n36971 ) ;
assign n36973 =  ( n144 ) ? ( n2957 ) : ( n36972 ) ;
assign n36974 =  ( n142 ) ? ( n2956 ) : ( n36973 ) ;
assign n36975 =  ( n10 ) ? ( n2955 ) : ( n36974 ) ;
assign n36976 =  ( n3032 ) ? ( VREG_14_0 ) : ( n36970 ) ;
assign n36977 =  ( n3032 ) ? ( VREG_14_0 ) : ( n36975 ) ;
assign n36978 =  ( n3034 ) ? ( n36977 ) : ( VREG_14_0 ) ;
assign n36979 =  ( n2965 ) ? ( n36976 ) : ( n36978 ) ;
assign n36980 =  ( n1930 ) ? ( n36975 ) : ( n36979 ) ;
assign n36981 =  ( n879 ) ? ( n36970 ) : ( n36980 ) ;
assign n36982 =  ( n172 ) ? ( n3045 ) : ( VREG_14_0 ) ;
assign n36983 =  ( n170 ) ? ( n3044 ) : ( n36982 ) ;
assign n36984 =  ( n168 ) ? ( n3043 ) : ( n36983 ) ;
assign n36985 =  ( n166 ) ? ( n3042 ) : ( n36984 ) ;
assign n36986 =  ( n162 ) ? ( n3041 ) : ( n36985 ) ;
assign n36987 =  ( n172 ) ? ( n3056 ) : ( VREG_14_0 ) ;
assign n36988 =  ( n170 ) ? ( n3055 ) : ( n36987 ) ;
assign n36989 =  ( n168 ) ? ( n3054 ) : ( n36988 ) ;
assign n36990 =  ( n166 ) ? ( n3053 ) : ( n36989 ) ;
assign n36991 =  ( n162 ) ? ( n3052 ) : ( n36990 ) ;
assign n36992 =  ( n3032 ) ? ( VREG_14_0 ) : ( n36991 ) ;
assign n36993 =  ( n3051 ) ? ( n36992 ) : ( VREG_14_0 ) ;
assign n36994 =  ( n3040 ) ? ( n36986 ) : ( n36993 ) ;
assign n36995 =  ( n192 ) ? ( VREG_14_0 ) : ( VREG_14_0 ) ;
assign n36996 =  ( n157 ) ? ( n36994 ) : ( n36995 ) ;
assign n36997 =  ( n6 ) ? ( n36981 ) : ( n36996 ) ;
assign n36998 =  ( n307 ) ? ( n36997 ) : ( VREG_14_0 ) ;
assign n36999 =  ( n148 ) ? ( n4113 ) : ( VREG_14_1 ) ;
assign n37000 =  ( n146 ) ? ( n4112 ) : ( n36999 ) ;
assign n37001 =  ( n144 ) ? ( n4111 ) : ( n37000 ) ;
assign n37002 =  ( n142 ) ? ( n4110 ) : ( n37001 ) ;
assign n37003 =  ( n10 ) ? ( n4109 ) : ( n37002 ) ;
assign n37004 =  ( n148 ) ? ( n5147 ) : ( VREG_14_1 ) ;
assign n37005 =  ( n146 ) ? ( n5146 ) : ( n37004 ) ;
assign n37006 =  ( n144 ) ? ( n5145 ) : ( n37005 ) ;
assign n37007 =  ( n142 ) ? ( n5144 ) : ( n37006 ) ;
assign n37008 =  ( n10 ) ? ( n5143 ) : ( n37007 ) ;
assign n37009 =  ( n5154 ) ? ( VREG_14_1 ) : ( n37003 ) ;
assign n37010 =  ( n5154 ) ? ( VREG_14_1 ) : ( n37008 ) ;
assign n37011 =  ( n3034 ) ? ( n37010 ) : ( VREG_14_1 ) ;
assign n37012 =  ( n2965 ) ? ( n37009 ) : ( n37011 ) ;
assign n37013 =  ( n1930 ) ? ( n37008 ) : ( n37012 ) ;
assign n37014 =  ( n879 ) ? ( n37003 ) : ( n37013 ) ;
assign n37015 =  ( n172 ) ? ( n5165 ) : ( VREG_14_1 ) ;
assign n37016 =  ( n170 ) ? ( n5164 ) : ( n37015 ) ;
assign n37017 =  ( n168 ) ? ( n5163 ) : ( n37016 ) ;
assign n37018 =  ( n166 ) ? ( n5162 ) : ( n37017 ) ;
assign n37019 =  ( n162 ) ? ( n5161 ) : ( n37018 ) ;
assign n37020 =  ( n172 ) ? ( n5175 ) : ( VREG_14_1 ) ;
assign n37021 =  ( n170 ) ? ( n5174 ) : ( n37020 ) ;
assign n37022 =  ( n168 ) ? ( n5173 ) : ( n37021 ) ;
assign n37023 =  ( n166 ) ? ( n5172 ) : ( n37022 ) ;
assign n37024 =  ( n162 ) ? ( n5171 ) : ( n37023 ) ;
assign n37025 =  ( n5154 ) ? ( VREG_14_1 ) : ( n37024 ) ;
assign n37026 =  ( n3051 ) ? ( n37025 ) : ( VREG_14_1 ) ;
assign n37027 =  ( n3040 ) ? ( n37019 ) : ( n37026 ) ;
assign n37028 =  ( n192 ) ? ( VREG_14_1 ) : ( VREG_14_1 ) ;
assign n37029 =  ( n157 ) ? ( n37027 ) : ( n37028 ) ;
assign n37030 =  ( n6 ) ? ( n37014 ) : ( n37029 ) ;
assign n37031 =  ( n307 ) ? ( n37030 ) : ( VREG_14_1 ) ;
assign n37032 =  ( n148 ) ? ( n6232 ) : ( VREG_14_10 ) ;
assign n37033 =  ( n146 ) ? ( n6231 ) : ( n37032 ) ;
assign n37034 =  ( n144 ) ? ( n6230 ) : ( n37033 ) ;
assign n37035 =  ( n142 ) ? ( n6229 ) : ( n37034 ) ;
assign n37036 =  ( n10 ) ? ( n6228 ) : ( n37035 ) ;
assign n37037 =  ( n148 ) ? ( n7266 ) : ( VREG_14_10 ) ;
assign n37038 =  ( n146 ) ? ( n7265 ) : ( n37037 ) ;
assign n37039 =  ( n144 ) ? ( n7264 ) : ( n37038 ) ;
assign n37040 =  ( n142 ) ? ( n7263 ) : ( n37039 ) ;
assign n37041 =  ( n10 ) ? ( n7262 ) : ( n37040 ) ;
assign n37042 =  ( n7273 ) ? ( VREG_14_10 ) : ( n37036 ) ;
assign n37043 =  ( n7273 ) ? ( VREG_14_10 ) : ( n37041 ) ;
assign n37044 =  ( n3034 ) ? ( n37043 ) : ( VREG_14_10 ) ;
assign n37045 =  ( n2965 ) ? ( n37042 ) : ( n37044 ) ;
assign n37046 =  ( n1930 ) ? ( n37041 ) : ( n37045 ) ;
assign n37047 =  ( n879 ) ? ( n37036 ) : ( n37046 ) ;
assign n37048 =  ( n172 ) ? ( n7284 ) : ( VREG_14_10 ) ;
assign n37049 =  ( n170 ) ? ( n7283 ) : ( n37048 ) ;
assign n37050 =  ( n168 ) ? ( n7282 ) : ( n37049 ) ;
assign n37051 =  ( n166 ) ? ( n7281 ) : ( n37050 ) ;
assign n37052 =  ( n162 ) ? ( n7280 ) : ( n37051 ) ;
assign n37053 =  ( n172 ) ? ( n7294 ) : ( VREG_14_10 ) ;
assign n37054 =  ( n170 ) ? ( n7293 ) : ( n37053 ) ;
assign n37055 =  ( n168 ) ? ( n7292 ) : ( n37054 ) ;
assign n37056 =  ( n166 ) ? ( n7291 ) : ( n37055 ) ;
assign n37057 =  ( n162 ) ? ( n7290 ) : ( n37056 ) ;
assign n37058 =  ( n7273 ) ? ( VREG_14_10 ) : ( n37057 ) ;
assign n37059 =  ( n3051 ) ? ( n37058 ) : ( VREG_14_10 ) ;
assign n37060 =  ( n3040 ) ? ( n37052 ) : ( n37059 ) ;
assign n37061 =  ( n192 ) ? ( VREG_14_10 ) : ( VREG_14_10 ) ;
assign n37062 =  ( n157 ) ? ( n37060 ) : ( n37061 ) ;
assign n37063 =  ( n6 ) ? ( n37047 ) : ( n37062 ) ;
assign n37064 =  ( n307 ) ? ( n37063 ) : ( VREG_14_10 ) ;
assign n37065 =  ( n148 ) ? ( n8351 ) : ( VREG_14_11 ) ;
assign n37066 =  ( n146 ) ? ( n8350 ) : ( n37065 ) ;
assign n37067 =  ( n144 ) ? ( n8349 ) : ( n37066 ) ;
assign n37068 =  ( n142 ) ? ( n8348 ) : ( n37067 ) ;
assign n37069 =  ( n10 ) ? ( n8347 ) : ( n37068 ) ;
assign n37070 =  ( n148 ) ? ( n9385 ) : ( VREG_14_11 ) ;
assign n37071 =  ( n146 ) ? ( n9384 ) : ( n37070 ) ;
assign n37072 =  ( n144 ) ? ( n9383 ) : ( n37071 ) ;
assign n37073 =  ( n142 ) ? ( n9382 ) : ( n37072 ) ;
assign n37074 =  ( n10 ) ? ( n9381 ) : ( n37073 ) ;
assign n37075 =  ( n9392 ) ? ( VREG_14_11 ) : ( n37069 ) ;
assign n37076 =  ( n9392 ) ? ( VREG_14_11 ) : ( n37074 ) ;
assign n37077 =  ( n3034 ) ? ( n37076 ) : ( VREG_14_11 ) ;
assign n37078 =  ( n2965 ) ? ( n37075 ) : ( n37077 ) ;
assign n37079 =  ( n1930 ) ? ( n37074 ) : ( n37078 ) ;
assign n37080 =  ( n879 ) ? ( n37069 ) : ( n37079 ) ;
assign n37081 =  ( n172 ) ? ( n9403 ) : ( VREG_14_11 ) ;
assign n37082 =  ( n170 ) ? ( n9402 ) : ( n37081 ) ;
assign n37083 =  ( n168 ) ? ( n9401 ) : ( n37082 ) ;
assign n37084 =  ( n166 ) ? ( n9400 ) : ( n37083 ) ;
assign n37085 =  ( n162 ) ? ( n9399 ) : ( n37084 ) ;
assign n37086 =  ( n172 ) ? ( n9413 ) : ( VREG_14_11 ) ;
assign n37087 =  ( n170 ) ? ( n9412 ) : ( n37086 ) ;
assign n37088 =  ( n168 ) ? ( n9411 ) : ( n37087 ) ;
assign n37089 =  ( n166 ) ? ( n9410 ) : ( n37088 ) ;
assign n37090 =  ( n162 ) ? ( n9409 ) : ( n37089 ) ;
assign n37091 =  ( n9392 ) ? ( VREG_14_11 ) : ( n37090 ) ;
assign n37092 =  ( n3051 ) ? ( n37091 ) : ( VREG_14_11 ) ;
assign n37093 =  ( n3040 ) ? ( n37085 ) : ( n37092 ) ;
assign n37094 =  ( n192 ) ? ( VREG_14_11 ) : ( VREG_14_11 ) ;
assign n37095 =  ( n157 ) ? ( n37093 ) : ( n37094 ) ;
assign n37096 =  ( n6 ) ? ( n37080 ) : ( n37095 ) ;
assign n37097 =  ( n307 ) ? ( n37096 ) : ( VREG_14_11 ) ;
assign n37098 =  ( n148 ) ? ( n10470 ) : ( VREG_14_12 ) ;
assign n37099 =  ( n146 ) ? ( n10469 ) : ( n37098 ) ;
assign n37100 =  ( n144 ) ? ( n10468 ) : ( n37099 ) ;
assign n37101 =  ( n142 ) ? ( n10467 ) : ( n37100 ) ;
assign n37102 =  ( n10 ) ? ( n10466 ) : ( n37101 ) ;
assign n37103 =  ( n148 ) ? ( n11504 ) : ( VREG_14_12 ) ;
assign n37104 =  ( n146 ) ? ( n11503 ) : ( n37103 ) ;
assign n37105 =  ( n144 ) ? ( n11502 ) : ( n37104 ) ;
assign n37106 =  ( n142 ) ? ( n11501 ) : ( n37105 ) ;
assign n37107 =  ( n10 ) ? ( n11500 ) : ( n37106 ) ;
assign n37108 =  ( n11511 ) ? ( VREG_14_12 ) : ( n37102 ) ;
assign n37109 =  ( n11511 ) ? ( VREG_14_12 ) : ( n37107 ) ;
assign n37110 =  ( n3034 ) ? ( n37109 ) : ( VREG_14_12 ) ;
assign n37111 =  ( n2965 ) ? ( n37108 ) : ( n37110 ) ;
assign n37112 =  ( n1930 ) ? ( n37107 ) : ( n37111 ) ;
assign n37113 =  ( n879 ) ? ( n37102 ) : ( n37112 ) ;
assign n37114 =  ( n172 ) ? ( n11522 ) : ( VREG_14_12 ) ;
assign n37115 =  ( n170 ) ? ( n11521 ) : ( n37114 ) ;
assign n37116 =  ( n168 ) ? ( n11520 ) : ( n37115 ) ;
assign n37117 =  ( n166 ) ? ( n11519 ) : ( n37116 ) ;
assign n37118 =  ( n162 ) ? ( n11518 ) : ( n37117 ) ;
assign n37119 =  ( n172 ) ? ( n11532 ) : ( VREG_14_12 ) ;
assign n37120 =  ( n170 ) ? ( n11531 ) : ( n37119 ) ;
assign n37121 =  ( n168 ) ? ( n11530 ) : ( n37120 ) ;
assign n37122 =  ( n166 ) ? ( n11529 ) : ( n37121 ) ;
assign n37123 =  ( n162 ) ? ( n11528 ) : ( n37122 ) ;
assign n37124 =  ( n11511 ) ? ( VREG_14_12 ) : ( n37123 ) ;
assign n37125 =  ( n3051 ) ? ( n37124 ) : ( VREG_14_12 ) ;
assign n37126 =  ( n3040 ) ? ( n37118 ) : ( n37125 ) ;
assign n37127 =  ( n192 ) ? ( VREG_14_12 ) : ( VREG_14_12 ) ;
assign n37128 =  ( n157 ) ? ( n37126 ) : ( n37127 ) ;
assign n37129 =  ( n6 ) ? ( n37113 ) : ( n37128 ) ;
assign n37130 =  ( n307 ) ? ( n37129 ) : ( VREG_14_12 ) ;
assign n37131 =  ( n148 ) ? ( n12589 ) : ( VREG_14_13 ) ;
assign n37132 =  ( n146 ) ? ( n12588 ) : ( n37131 ) ;
assign n37133 =  ( n144 ) ? ( n12587 ) : ( n37132 ) ;
assign n37134 =  ( n142 ) ? ( n12586 ) : ( n37133 ) ;
assign n37135 =  ( n10 ) ? ( n12585 ) : ( n37134 ) ;
assign n37136 =  ( n148 ) ? ( n13623 ) : ( VREG_14_13 ) ;
assign n37137 =  ( n146 ) ? ( n13622 ) : ( n37136 ) ;
assign n37138 =  ( n144 ) ? ( n13621 ) : ( n37137 ) ;
assign n37139 =  ( n142 ) ? ( n13620 ) : ( n37138 ) ;
assign n37140 =  ( n10 ) ? ( n13619 ) : ( n37139 ) ;
assign n37141 =  ( n13630 ) ? ( VREG_14_13 ) : ( n37135 ) ;
assign n37142 =  ( n13630 ) ? ( VREG_14_13 ) : ( n37140 ) ;
assign n37143 =  ( n3034 ) ? ( n37142 ) : ( VREG_14_13 ) ;
assign n37144 =  ( n2965 ) ? ( n37141 ) : ( n37143 ) ;
assign n37145 =  ( n1930 ) ? ( n37140 ) : ( n37144 ) ;
assign n37146 =  ( n879 ) ? ( n37135 ) : ( n37145 ) ;
assign n37147 =  ( n172 ) ? ( n13641 ) : ( VREG_14_13 ) ;
assign n37148 =  ( n170 ) ? ( n13640 ) : ( n37147 ) ;
assign n37149 =  ( n168 ) ? ( n13639 ) : ( n37148 ) ;
assign n37150 =  ( n166 ) ? ( n13638 ) : ( n37149 ) ;
assign n37151 =  ( n162 ) ? ( n13637 ) : ( n37150 ) ;
assign n37152 =  ( n172 ) ? ( n13651 ) : ( VREG_14_13 ) ;
assign n37153 =  ( n170 ) ? ( n13650 ) : ( n37152 ) ;
assign n37154 =  ( n168 ) ? ( n13649 ) : ( n37153 ) ;
assign n37155 =  ( n166 ) ? ( n13648 ) : ( n37154 ) ;
assign n37156 =  ( n162 ) ? ( n13647 ) : ( n37155 ) ;
assign n37157 =  ( n13630 ) ? ( VREG_14_13 ) : ( n37156 ) ;
assign n37158 =  ( n3051 ) ? ( n37157 ) : ( VREG_14_13 ) ;
assign n37159 =  ( n3040 ) ? ( n37151 ) : ( n37158 ) ;
assign n37160 =  ( n192 ) ? ( VREG_14_13 ) : ( VREG_14_13 ) ;
assign n37161 =  ( n157 ) ? ( n37159 ) : ( n37160 ) ;
assign n37162 =  ( n6 ) ? ( n37146 ) : ( n37161 ) ;
assign n37163 =  ( n307 ) ? ( n37162 ) : ( VREG_14_13 ) ;
assign n37164 =  ( n148 ) ? ( n14708 ) : ( VREG_14_14 ) ;
assign n37165 =  ( n146 ) ? ( n14707 ) : ( n37164 ) ;
assign n37166 =  ( n144 ) ? ( n14706 ) : ( n37165 ) ;
assign n37167 =  ( n142 ) ? ( n14705 ) : ( n37166 ) ;
assign n37168 =  ( n10 ) ? ( n14704 ) : ( n37167 ) ;
assign n37169 =  ( n148 ) ? ( n15742 ) : ( VREG_14_14 ) ;
assign n37170 =  ( n146 ) ? ( n15741 ) : ( n37169 ) ;
assign n37171 =  ( n144 ) ? ( n15740 ) : ( n37170 ) ;
assign n37172 =  ( n142 ) ? ( n15739 ) : ( n37171 ) ;
assign n37173 =  ( n10 ) ? ( n15738 ) : ( n37172 ) ;
assign n37174 =  ( n15749 ) ? ( VREG_14_14 ) : ( n37168 ) ;
assign n37175 =  ( n15749 ) ? ( VREG_14_14 ) : ( n37173 ) ;
assign n37176 =  ( n3034 ) ? ( n37175 ) : ( VREG_14_14 ) ;
assign n37177 =  ( n2965 ) ? ( n37174 ) : ( n37176 ) ;
assign n37178 =  ( n1930 ) ? ( n37173 ) : ( n37177 ) ;
assign n37179 =  ( n879 ) ? ( n37168 ) : ( n37178 ) ;
assign n37180 =  ( n172 ) ? ( n15760 ) : ( VREG_14_14 ) ;
assign n37181 =  ( n170 ) ? ( n15759 ) : ( n37180 ) ;
assign n37182 =  ( n168 ) ? ( n15758 ) : ( n37181 ) ;
assign n37183 =  ( n166 ) ? ( n15757 ) : ( n37182 ) ;
assign n37184 =  ( n162 ) ? ( n15756 ) : ( n37183 ) ;
assign n37185 =  ( n172 ) ? ( n15770 ) : ( VREG_14_14 ) ;
assign n37186 =  ( n170 ) ? ( n15769 ) : ( n37185 ) ;
assign n37187 =  ( n168 ) ? ( n15768 ) : ( n37186 ) ;
assign n37188 =  ( n166 ) ? ( n15767 ) : ( n37187 ) ;
assign n37189 =  ( n162 ) ? ( n15766 ) : ( n37188 ) ;
assign n37190 =  ( n15749 ) ? ( VREG_14_14 ) : ( n37189 ) ;
assign n37191 =  ( n3051 ) ? ( n37190 ) : ( VREG_14_14 ) ;
assign n37192 =  ( n3040 ) ? ( n37184 ) : ( n37191 ) ;
assign n37193 =  ( n192 ) ? ( VREG_14_14 ) : ( VREG_14_14 ) ;
assign n37194 =  ( n157 ) ? ( n37192 ) : ( n37193 ) ;
assign n37195 =  ( n6 ) ? ( n37179 ) : ( n37194 ) ;
assign n37196 =  ( n307 ) ? ( n37195 ) : ( VREG_14_14 ) ;
assign n37197 =  ( n148 ) ? ( n16827 ) : ( VREG_14_15 ) ;
assign n37198 =  ( n146 ) ? ( n16826 ) : ( n37197 ) ;
assign n37199 =  ( n144 ) ? ( n16825 ) : ( n37198 ) ;
assign n37200 =  ( n142 ) ? ( n16824 ) : ( n37199 ) ;
assign n37201 =  ( n10 ) ? ( n16823 ) : ( n37200 ) ;
assign n37202 =  ( n148 ) ? ( n17861 ) : ( VREG_14_15 ) ;
assign n37203 =  ( n146 ) ? ( n17860 ) : ( n37202 ) ;
assign n37204 =  ( n144 ) ? ( n17859 ) : ( n37203 ) ;
assign n37205 =  ( n142 ) ? ( n17858 ) : ( n37204 ) ;
assign n37206 =  ( n10 ) ? ( n17857 ) : ( n37205 ) ;
assign n37207 =  ( n17868 ) ? ( VREG_14_15 ) : ( n37201 ) ;
assign n37208 =  ( n17868 ) ? ( VREG_14_15 ) : ( n37206 ) ;
assign n37209 =  ( n3034 ) ? ( n37208 ) : ( VREG_14_15 ) ;
assign n37210 =  ( n2965 ) ? ( n37207 ) : ( n37209 ) ;
assign n37211 =  ( n1930 ) ? ( n37206 ) : ( n37210 ) ;
assign n37212 =  ( n879 ) ? ( n37201 ) : ( n37211 ) ;
assign n37213 =  ( n172 ) ? ( n17879 ) : ( VREG_14_15 ) ;
assign n37214 =  ( n170 ) ? ( n17878 ) : ( n37213 ) ;
assign n37215 =  ( n168 ) ? ( n17877 ) : ( n37214 ) ;
assign n37216 =  ( n166 ) ? ( n17876 ) : ( n37215 ) ;
assign n37217 =  ( n162 ) ? ( n17875 ) : ( n37216 ) ;
assign n37218 =  ( n172 ) ? ( n17889 ) : ( VREG_14_15 ) ;
assign n37219 =  ( n170 ) ? ( n17888 ) : ( n37218 ) ;
assign n37220 =  ( n168 ) ? ( n17887 ) : ( n37219 ) ;
assign n37221 =  ( n166 ) ? ( n17886 ) : ( n37220 ) ;
assign n37222 =  ( n162 ) ? ( n17885 ) : ( n37221 ) ;
assign n37223 =  ( n17868 ) ? ( VREG_14_15 ) : ( n37222 ) ;
assign n37224 =  ( n3051 ) ? ( n37223 ) : ( VREG_14_15 ) ;
assign n37225 =  ( n3040 ) ? ( n37217 ) : ( n37224 ) ;
assign n37226 =  ( n192 ) ? ( VREG_14_15 ) : ( VREG_14_15 ) ;
assign n37227 =  ( n157 ) ? ( n37225 ) : ( n37226 ) ;
assign n37228 =  ( n6 ) ? ( n37212 ) : ( n37227 ) ;
assign n37229 =  ( n307 ) ? ( n37228 ) : ( VREG_14_15 ) ;
assign n37230 =  ( n148 ) ? ( n18946 ) : ( VREG_14_2 ) ;
assign n37231 =  ( n146 ) ? ( n18945 ) : ( n37230 ) ;
assign n37232 =  ( n144 ) ? ( n18944 ) : ( n37231 ) ;
assign n37233 =  ( n142 ) ? ( n18943 ) : ( n37232 ) ;
assign n37234 =  ( n10 ) ? ( n18942 ) : ( n37233 ) ;
assign n37235 =  ( n148 ) ? ( n19980 ) : ( VREG_14_2 ) ;
assign n37236 =  ( n146 ) ? ( n19979 ) : ( n37235 ) ;
assign n37237 =  ( n144 ) ? ( n19978 ) : ( n37236 ) ;
assign n37238 =  ( n142 ) ? ( n19977 ) : ( n37237 ) ;
assign n37239 =  ( n10 ) ? ( n19976 ) : ( n37238 ) ;
assign n37240 =  ( n19987 ) ? ( VREG_14_2 ) : ( n37234 ) ;
assign n37241 =  ( n19987 ) ? ( VREG_14_2 ) : ( n37239 ) ;
assign n37242 =  ( n3034 ) ? ( n37241 ) : ( VREG_14_2 ) ;
assign n37243 =  ( n2965 ) ? ( n37240 ) : ( n37242 ) ;
assign n37244 =  ( n1930 ) ? ( n37239 ) : ( n37243 ) ;
assign n37245 =  ( n879 ) ? ( n37234 ) : ( n37244 ) ;
assign n37246 =  ( n172 ) ? ( n19998 ) : ( VREG_14_2 ) ;
assign n37247 =  ( n170 ) ? ( n19997 ) : ( n37246 ) ;
assign n37248 =  ( n168 ) ? ( n19996 ) : ( n37247 ) ;
assign n37249 =  ( n166 ) ? ( n19995 ) : ( n37248 ) ;
assign n37250 =  ( n162 ) ? ( n19994 ) : ( n37249 ) ;
assign n37251 =  ( n172 ) ? ( n20008 ) : ( VREG_14_2 ) ;
assign n37252 =  ( n170 ) ? ( n20007 ) : ( n37251 ) ;
assign n37253 =  ( n168 ) ? ( n20006 ) : ( n37252 ) ;
assign n37254 =  ( n166 ) ? ( n20005 ) : ( n37253 ) ;
assign n37255 =  ( n162 ) ? ( n20004 ) : ( n37254 ) ;
assign n37256 =  ( n19987 ) ? ( VREG_14_2 ) : ( n37255 ) ;
assign n37257 =  ( n3051 ) ? ( n37256 ) : ( VREG_14_2 ) ;
assign n37258 =  ( n3040 ) ? ( n37250 ) : ( n37257 ) ;
assign n37259 =  ( n192 ) ? ( VREG_14_2 ) : ( VREG_14_2 ) ;
assign n37260 =  ( n157 ) ? ( n37258 ) : ( n37259 ) ;
assign n37261 =  ( n6 ) ? ( n37245 ) : ( n37260 ) ;
assign n37262 =  ( n307 ) ? ( n37261 ) : ( VREG_14_2 ) ;
assign n37263 =  ( n148 ) ? ( n21065 ) : ( VREG_14_3 ) ;
assign n37264 =  ( n146 ) ? ( n21064 ) : ( n37263 ) ;
assign n37265 =  ( n144 ) ? ( n21063 ) : ( n37264 ) ;
assign n37266 =  ( n142 ) ? ( n21062 ) : ( n37265 ) ;
assign n37267 =  ( n10 ) ? ( n21061 ) : ( n37266 ) ;
assign n37268 =  ( n148 ) ? ( n22099 ) : ( VREG_14_3 ) ;
assign n37269 =  ( n146 ) ? ( n22098 ) : ( n37268 ) ;
assign n37270 =  ( n144 ) ? ( n22097 ) : ( n37269 ) ;
assign n37271 =  ( n142 ) ? ( n22096 ) : ( n37270 ) ;
assign n37272 =  ( n10 ) ? ( n22095 ) : ( n37271 ) ;
assign n37273 =  ( n22106 ) ? ( VREG_14_3 ) : ( n37267 ) ;
assign n37274 =  ( n22106 ) ? ( VREG_14_3 ) : ( n37272 ) ;
assign n37275 =  ( n3034 ) ? ( n37274 ) : ( VREG_14_3 ) ;
assign n37276 =  ( n2965 ) ? ( n37273 ) : ( n37275 ) ;
assign n37277 =  ( n1930 ) ? ( n37272 ) : ( n37276 ) ;
assign n37278 =  ( n879 ) ? ( n37267 ) : ( n37277 ) ;
assign n37279 =  ( n172 ) ? ( n22117 ) : ( VREG_14_3 ) ;
assign n37280 =  ( n170 ) ? ( n22116 ) : ( n37279 ) ;
assign n37281 =  ( n168 ) ? ( n22115 ) : ( n37280 ) ;
assign n37282 =  ( n166 ) ? ( n22114 ) : ( n37281 ) ;
assign n37283 =  ( n162 ) ? ( n22113 ) : ( n37282 ) ;
assign n37284 =  ( n172 ) ? ( n22127 ) : ( VREG_14_3 ) ;
assign n37285 =  ( n170 ) ? ( n22126 ) : ( n37284 ) ;
assign n37286 =  ( n168 ) ? ( n22125 ) : ( n37285 ) ;
assign n37287 =  ( n166 ) ? ( n22124 ) : ( n37286 ) ;
assign n37288 =  ( n162 ) ? ( n22123 ) : ( n37287 ) ;
assign n37289 =  ( n22106 ) ? ( VREG_14_3 ) : ( n37288 ) ;
assign n37290 =  ( n3051 ) ? ( n37289 ) : ( VREG_14_3 ) ;
assign n37291 =  ( n3040 ) ? ( n37283 ) : ( n37290 ) ;
assign n37292 =  ( n192 ) ? ( VREG_14_3 ) : ( VREG_14_3 ) ;
assign n37293 =  ( n157 ) ? ( n37291 ) : ( n37292 ) ;
assign n37294 =  ( n6 ) ? ( n37278 ) : ( n37293 ) ;
assign n37295 =  ( n307 ) ? ( n37294 ) : ( VREG_14_3 ) ;
assign n37296 =  ( n148 ) ? ( n23184 ) : ( VREG_14_4 ) ;
assign n37297 =  ( n146 ) ? ( n23183 ) : ( n37296 ) ;
assign n37298 =  ( n144 ) ? ( n23182 ) : ( n37297 ) ;
assign n37299 =  ( n142 ) ? ( n23181 ) : ( n37298 ) ;
assign n37300 =  ( n10 ) ? ( n23180 ) : ( n37299 ) ;
assign n37301 =  ( n148 ) ? ( n24218 ) : ( VREG_14_4 ) ;
assign n37302 =  ( n146 ) ? ( n24217 ) : ( n37301 ) ;
assign n37303 =  ( n144 ) ? ( n24216 ) : ( n37302 ) ;
assign n37304 =  ( n142 ) ? ( n24215 ) : ( n37303 ) ;
assign n37305 =  ( n10 ) ? ( n24214 ) : ( n37304 ) ;
assign n37306 =  ( n24225 ) ? ( VREG_14_4 ) : ( n37300 ) ;
assign n37307 =  ( n24225 ) ? ( VREG_14_4 ) : ( n37305 ) ;
assign n37308 =  ( n3034 ) ? ( n37307 ) : ( VREG_14_4 ) ;
assign n37309 =  ( n2965 ) ? ( n37306 ) : ( n37308 ) ;
assign n37310 =  ( n1930 ) ? ( n37305 ) : ( n37309 ) ;
assign n37311 =  ( n879 ) ? ( n37300 ) : ( n37310 ) ;
assign n37312 =  ( n172 ) ? ( n24236 ) : ( VREG_14_4 ) ;
assign n37313 =  ( n170 ) ? ( n24235 ) : ( n37312 ) ;
assign n37314 =  ( n168 ) ? ( n24234 ) : ( n37313 ) ;
assign n37315 =  ( n166 ) ? ( n24233 ) : ( n37314 ) ;
assign n37316 =  ( n162 ) ? ( n24232 ) : ( n37315 ) ;
assign n37317 =  ( n172 ) ? ( n24246 ) : ( VREG_14_4 ) ;
assign n37318 =  ( n170 ) ? ( n24245 ) : ( n37317 ) ;
assign n37319 =  ( n168 ) ? ( n24244 ) : ( n37318 ) ;
assign n37320 =  ( n166 ) ? ( n24243 ) : ( n37319 ) ;
assign n37321 =  ( n162 ) ? ( n24242 ) : ( n37320 ) ;
assign n37322 =  ( n24225 ) ? ( VREG_14_4 ) : ( n37321 ) ;
assign n37323 =  ( n3051 ) ? ( n37322 ) : ( VREG_14_4 ) ;
assign n37324 =  ( n3040 ) ? ( n37316 ) : ( n37323 ) ;
assign n37325 =  ( n192 ) ? ( VREG_14_4 ) : ( VREG_14_4 ) ;
assign n37326 =  ( n157 ) ? ( n37324 ) : ( n37325 ) ;
assign n37327 =  ( n6 ) ? ( n37311 ) : ( n37326 ) ;
assign n37328 =  ( n307 ) ? ( n37327 ) : ( VREG_14_4 ) ;
assign n37329 =  ( n148 ) ? ( n25303 ) : ( VREG_14_5 ) ;
assign n37330 =  ( n146 ) ? ( n25302 ) : ( n37329 ) ;
assign n37331 =  ( n144 ) ? ( n25301 ) : ( n37330 ) ;
assign n37332 =  ( n142 ) ? ( n25300 ) : ( n37331 ) ;
assign n37333 =  ( n10 ) ? ( n25299 ) : ( n37332 ) ;
assign n37334 =  ( n148 ) ? ( n26337 ) : ( VREG_14_5 ) ;
assign n37335 =  ( n146 ) ? ( n26336 ) : ( n37334 ) ;
assign n37336 =  ( n144 ) ? ( n26335 ) : ( n37335 ) ;
assign n37337 =  ( n142 ) ? ( n26334 ) : ( n37336 ) ;
assign n37338 =  ( n10 ) ? ( n26333 ) : ( n37337 ) ;
assign n37339 =  ( n26344 ) ? ( VREG_14_5 ) : ( n37333 ) ;
assign n37340 =  ( n26344 ) ? ( VREG_14_5 ) : ( n37338 ) ;
assign n37341 =  ( n3034 ) ? ( n37340 ) : ( VREG_14_5 ) ;
assign n37342 =  ( n2965 ) ? ( n37339 ) : ( n37341 ) ;
assign n37343 =  ( n1930 ) ? ( n37338 ) : ( n37342 ) ;
assign n37344 =  ( n879 ) ? ( n37333 ) : ( n37343 ) ;
assign n37345 =  ( n172 ) ? ( n26355 ) : ( VREG_14_5 ) ;
assign n37346 =  ( n170 ) ? ( n26354 ) : ( n37345 ) ;
assign n37347 =  ( n168 ) ? ( n26353 ) : ( n37346 ) ;
assign n37348 =  ( n166 ) ? ( n26352 ) : ( n37347 ) ;
assign n37349 =  ( n162 ) ? ( n26351 ) : ( n37348 ) ;
assign n37350 =  ( n172 ) ? ( n26365 ) : ( VREG_14_5 ) ;
assign n37351 =  ( n170 ) ? ( n26364 ) : ( n37350 ) ;
assign n37352 =  ( n168 ) ? ( n26363 ) : ( n37351 ) ;
assign n37353 =  ( n166 ) ? ( n26362 ) : ( n37352 ) ;
assign n37354 =  ( n162 ) ? ( n26361 ) : ( n37353 ) ;
assign n37355 =  ( n26344 ) ? ( VREG_14_5 ) : ( n37354 ) ;
assign n37356 =  ( n3051 ) ? ( n37355 ) : ( VREG_14_5 ) ;
assign n37357 =  ( n3040 ) ? ( n37349 ) : ( n37356 ) ;
assign n37358 =  ( n192 ) ? ( VREG_14_5 ) : ( VREG_14_5 ) ;
assign n37359 =  ( n157 ) ? ( n37357 ) : ( n37358 ) ;
assign n37360 =  ( n6 ) ? ( n37344 ) : ( n37359 ) ;
assign n37361 =  ( n307 ) ? ( n37360 ) : ( VREG_14_5 ) ;
assign n37362 =  ( n148 ) ? ( n27422 ) : ( VREG_14_6 ) ;
assign n37363 =  ( n146 ) ? ( n27421 ) : ( n37362 ) ;
assign n37364 =  ( n144 ) ? ( n27420 ) : ( n37363 ) ;
assign n37365 =  ( n142 ) ? ( n27419 ) : ( n37364 ) ;
assign n37366 =  ( n10 ) ? ( n27418 ) : ( n37365 ) ;
assign n37367 =  ( n148 ) ? ( n28456 ) : ( VREG_14_6 ) ;
assign n37368 =  ( n146 ) ? ( n28455 ) : ( n37367 ) ;
assign n37369 =  ( n144 ) ? ( n28454 ) : ( n37368 ) ;
assign n37370 =  ( n142 ) ? ( n28453 ) : ( n37369 ) ;
assign n37371 =  ( n10 ) ? ( n28452 ) : ( n37370 ) ;
assign n37372 =  ( n28463 ) ? ( VREG_14_6 ) : ( n37366 ) ;
assign n37373 =  ( n28463 ) ? ( VREG_14_6 ) : ( n37371 ) ;
assign n37374 =  ( n3034 ) ? ( n37373 ) : ( VREG_14_6 ) ;
assign n37375 =  ( n2965 ) ? ( n37372 ) : ( n37374 ) ;
assign n37376 =  ( n1930 ) ? ( n37371 ) : ( n37375 ) ;
assign n37377 =  ( n879 ) ? ( n37366 ) : ( n37376 ) ;
assign n37378 =  ( n172 ) ? ( n28474 ) : ( VREG_14_6 ) ;
assign n37379 =  ( n170 ) ? ( n28473 ) : ( n37378 ) ;
assign n37380 =  ( n168 ) ? ( n28472 ) : ( n37379 ) ;
assign n37381 =  ( n166 ) ? ( n28471 ) : ( n37380 ) ;
assign n37382 =  ( n162 ) ? ( n28470 ) : ( n37381 ) ;
assign n37383 =  ( n172 ) ? ( n28484 ) : ( VREG_14_6 ) ;
assign n37384 =  ( n170 ) ? ( n28483 ) : ( n37383 ) ;
assign n37385 =  ( n168 ) ? ( n28482 ) : ( n37384 ) ;
assign n37386 =  ( n166 ) ? ( n28481 ) : ( n37385 ) ;
assign n37387 =  ( n162 ) ? ( n28480 ) : ( n37386 ) ;
assign n37388 =  ( n28463 ) ? ( VREG_14_6 ) : ( n37387 ) ;
assign n37389 =  ( n3051 ) ? ( n37388 ) : ( VREG_14_6 ) ;
assign n37390 =  ( n3040 ) ? ( n37382 ) : ( n37389 ) ;
assign n37391 =  ( n192 ) ? ( VREG_14_6 ) : ( VREG_14_6 ) ;
assign n37392 =  ( n157 ) ? ( n37390 ) : ( n37391 ) ;
assign n37393 =  ( n6 ) ? ( n37377 ) : ( n37392 ) ;
assign n37394 =  ( n307 ) ? ( n37393 ) : ( VREG_14_6 ) ;
assign n37395 =  ( n148 ) ? ( n29541 ) : ( VREG_14_7 ) ;
assign n37396 =  ( n146 ) ? ( n29540 ) : ( n37395 ) ;
assign n37397 =  ( n144 ) ? ( n29539 ) : ( n37396 ) ;
assign n37398 =  ( n142 ) ? ( n29538 ) : ( n37397 ) ;
assign n37399 =  ( n10 ) ? ( n29537 ) : ( n37398 ) ;
assign n37400 =  ( n148 ) ? ( n30575 ) : ( VREG_14_7 ) ;
assign n37401 =  ( n146 ) ? ( n30574 ) : ( n37400 ) ;
assign n37402 =  ( n144 ) ? ( n30573 ) : ( n37401 ) ;
assign n37403 =  ( n142 ) ? ( n30572 ) : ( n37402 ) ;
assign n37404 =  ( n10 ) ? ( n30571 ) : ( n37403 ) ;
assign n37405 =  ( n30582 ) ? ( VREG_14_7 ) : ( n37399 ) ;
assign n37406 =  ( n30582 ) ? ( VREG_14_7 ) : ( n37404 ) ;
assign n37407 =  ( n3034 ) ? ( n37406 ) : ( VREG_14_7 ) ;
assign n37408 =  ( n2965 ) ? ( n37405 ) : ( n37407 ) ;
assign n37409 =  ( n1930 ) ? ( n37404 ) : ( n37408 ) ;
assign n37410 =  ( n879 ) ? ( n37399 ) : ( n37409 ) ;
assign n37411 =  ( n172 ) ? ( n30593 ) : ( VREG_14_7 ) ;
assign n37412 =  ( n170 ) ? ( n30592 ) : ( n37411 ) ;
assign n37413 =  ( n168 ) ? ( n30591 ) : ( n37412 ) ;
assign n37414 =  ( n166 ) ? ( n30590 ) : ( n37413 ) ;
assign n37415 =  ( n162 ) ? ( n30589 ) : ( n37414 ) ;
assign n37416 =  ( n172 ) ? ( n30603 ) : ( VREG_14_7 ) ;
assign n37417 =  ( n170 ) ? ( n30602 ) : ( n37416 ) ;
assign n37418 =  ( n168 ) ? ( n30601 ) : ( n37417 ) ;
assign n37419 =  ( n166 ) ? ( n30600 ) : ( n37418 ) ;
assign n37420 =  ( n162 ) ? ( n30599 ) : ( n37419 ) ;
assign n37421 =  ( n30582 ) ? ( VREG_14_7 ) : ( n37420 ) ;
assign n37422 =  ( n3051 ) ? ( n37421 ) : ( VREG_14_7 ) ;
assign n37423 =  ( n3040 ) ? ( n37415 ) : ( n37422 ) ;
assign n37424 =  ( n192 ) ? ( VREG_14_7 ) : ( VREG_14_7 ) ;
assign n37425 =  ( n157 ) ? ( n37423 ) : ( n37424 ) ;
assign n37426 =  ( n6 ) ? ( n37410 ) : ( n37425 ) ;
assign n37427 =  ( n307 ) ? ( n37426 ) : ( VREG_14_7 ) ;
assign n37428 =  ( n148 ) ? ( n31660 ) : ( VREG_14_8 ) ;
assign n37429 =  ( n146 ) ? ( n31659 ) : ( n37428 ) ;
assign n37430 =  ( n144 ) ? ( n31658 ) : ( n37429 ) ;
assign n37431 =  ( n142 ) ? ( n31657 ) : ( n37430 ) ;
assign n37432 =  ( n10 ) ? ( n31656 ) : ( n37431 ) ;
assign n37433 =  ( n148 ) ? ( n32694 ) : ( VREG_14_8 ) ;
assign n37434 =  ( n146 ) ? ( n32693 ) : ( n37433 ) ;
assign n37435 =  ( n144 ) ? ( n32692 ) : ( n37434 ) ;
assign n37436 =  ( n142 ) ? ( n32691 ) : ( n37435 ) ;
assign n37437 =  ( n10 ) ? ( n32690 ) : ( n37436 ) ;
assign n37438 =  ( n32701 ) ? ( VREG_14_8 ) : ( n37432 ) ;
assign n37439 =  ( n32701 ) ? ( VREG_14_8 ) : ( n37437 ) ;
assign n37440 =  ( n3034 ) ? ( n37439 ) : ( VREG_14_8 ) ;
assign n37441 =  ( n2965 ) ? ( n37438 ) : ( n37440 ) ;
assign n37442 =  ( n1930 ) ? ( n37437 ) : ( n37441 ) ;
assign n37443 =  ( n879 ) ? ( n37432 ) : ( n37442 ) ;
assign n37444 =  ( n172 ) ? ( n32712 ) : ( VREG_14_8 ) ;
assign n37445 =  ( n170 ) ? ( n32711 ) : ( n37444 ) ;
assign n37446 =  ( n168 ) ? ( n32710 ) : ( n37445 ) ;
assign n37447 =  ( n166 ) ? ( n32709 ) : ( n37446 ) ;
assign n37448 =  ( n162 ) ? ( n32708 ) : ( n37447 ) ;
assign n37449 =  ( n172 ) ? ( n32722 ) : ( VREG_14_8 ) ;
assign n37450 =  ( n170 ) ? ( n32721 ) : ( n37449 ) ;
assign n37451 =  ( n168 ) ? ( n32720 ) : ( n37450 ) ;
assign n37452 =  ( n166 ) ? ( n32719 ) : ( n37451 ) ;
assign n37453 =  ( n162 ) ? ( n32718 ) : ( n37452 ) ;
assign n37454 =  ( n32701 ) ? ( VREG_14_8 ) : ( n37453 ) ;
assign n37455 =  ( n3051 ) ? ( n37454 ) : ( VREG_14_8 ) ;
assign n37456 =  ( n3040 ) ? ( n37448 ) : ( n37455 ) ;
assign n37457 =  ( n192 ) ? ( VREG_14_8 ) : ( VREG_14_8 ) ;
assign n37458 =  ( n157 ) ? ( n37456 ) : ( n37457 ) ;
assign n37459 =  ( n6 ) ? ( n37443 ) : ( n37458 ) ;
assign n37460 =  ( n307 ) ? ( n37459 ) : ( VREG_14_8 ) ;
assign n37461 =  ( n148 ) ? ( n33779 ) : ( VREG_14_9 ) ;
assign n37462 =  ( n146 ) ? ( n33778 ) : ( n37461 ) ;
assign n37463 =  ( n144 ) ? ( n33777 ) : ( n37462 ) ;
assign n37464 =  ( n142 ) ? ( n33776 ) : ( n37463 ) ;
assign n37465 =  ( n10 ) ? ( n33775 ) : ( n37464 ) ;
assign n37466 =  ( n148 ) ? ( n34813 ) : ( VREG_14_9 ) ;
assign n37467 =  ( n146 ) ? ( n34812 ) : ( n37466 ) ;
assign n37468 =  ( n144 ) ? ( n34811 ) : ( n37467 ) ;
assign n37469 =  ( n142 ) ? ( n34810 ) : ( n37468 ) ;
assign n37470 =  ( n10 ) ? ( n34809 ) : ( n37469 ) ;
assign n37471 =  ( n34820 ) ? ( VREG_14_9 ) : ( n37465 ) ;
assign n37472 =  ( n34820 ) ? ( VREG_14_9 ) : ( n37470 ) ;
assign n37473 =  ( n3034 ) ? ( n37472 ) : ( VREG_14_9 ) ;
assign n37474 =  ( n2965 ) ? ( n37471 ) : ( n37473 ) ;
assign n37475 =  ( n1930 ) ? ( n37470 ) : ( n37474 ) ;
assign n37476 =  ( n879 ) ? ( n37465 ) : ( n37475 ) ;
assign n37477 =  ( n172 ) ? ( n34831 ) : ( VREG_14_9 ) ;
assign n37478 =  ( n170 ) ? ( n34830 ) : ( n37477 ) ;
assign n37479 =  ( n168 ) ? ( n34829 ) : ( n37478 ) ;
assign n37480 =  ( n166 ) ? ( n34828 ) : ( n37479 ) ;
assign n37481 =  ( n162 ) ? ( n34827 ) : ( n37480 ) ;
assign n37482 =  ( n172 ) ? ( n34841 ) : ( VREG_14_9 ) ;
assign n37483 =  ( n170 ) ? ( n34840 ) : ( n37482 ) ;
assign n37484 =  ( n168 ) ? ( n34839 ) : ( n37483 ) ;
assign n37485 =  ( n166 ) ? ( n34838 ) : ( n37484 ) ;
assign n37486 =  ( n162 ) ? ( n34837 ) : ( n37485 ) ;
assign n37487 =  ( n34820 ) ? ( VREG_14_9 ) : ( n37486 ) ;
assign n37488 =  ( n3051 ) ? ( n37487 ) : ( VREG_14_9 ) ;
assign n37489 =  ( n3040 ) ? ( n37481 ) : ( n37488 ) ;
assign n37490 =  ( n192 ) ? ( VREG_14_9 ) : ( VREG_14_9 ) ;
assign n37491 =  ( n157 ) ? ( n37489 ) : ( n37490 ) ;
assign n37492 =  ( n6 ) ? ( n37476 ) : ( n37491 ) ;
assign n37493 =  ( n307 ) ? ( n37492 ) : ( VREG_14_9 ) ;
assign n37494 =  ( n148 ) ? ( n1924 ) : ( VREG_15_0 ) ;
assign n37495 =  ( n146 ) ? ( n1923 ) : ( n37494 ) ;
assign n37496 =  ( n144 ) ? ( n1922 ) : ( n37495 ) ;
assign n37497 =  ( n142 ) ? ( n1921 ) : ( n37496 ) ;
assign n37498 =  ( n10 ) ? ( n1920 ) : ( n37497 ) ;
assign n37499 =  ( n148 ) ? ( n2959 ) : ( VREG_15_0 ) ;
assign n37500 =  ( n146 ) ? ( n2958 ) : ( n37499 ) ;
assign n37501 =  ( n144 ) ? ( n2957 ) : ( n37500 ) ;
assign n37502 =  ( n142 ) ? ( n2956 ) : ( n37501 ) ;
assign n37503 =  ( n10 ) ? ( n2955 ) : ( n37502 ) ;
assign n37504 =  ( n3032 ) ? ( VREG_15_0 ) : ( n37498 ) ;
assign n37505 =  ( n3032 ) ? ( VREG_15_0 ) : ( n37503 ) ;
assign n37506 =  ( n3034 ) ? ( n37505 ) : ( VREG_15_0 ) ;
assign n37507 =  ( n2965 ) ? ( n37504 ) : ( n37506 ) ;
assign n37508 =  ( n1930 ) ? ( n37503 ) : ( n37507 ) ;
assign n37509 =  ( n879 ) ? ( n37498 ) : ( n37508 ) ;
assign n37510 =  ( n172 ) ? ( n3045 ) : ( VREG_15_0 ) ;
assign n37511 =  ( n170 ) ? ( n3044 ) : ( n37510 ) ;
assign n37512 =  ( n168 ) ? ( n3043 ) : ( n37511 ) ;
assign n37513 =  ( n166 ) ? ( n3042 ) : ( n37512 ) ;
assign n37514 =  ( n162 ) ? ( n3041 ) : ( n37513 ) ;
assign n37515 =  ( n172 ) ? ( n3056 ) : ( VREG_15_0 ) ;
assign n37516 =  ( n170 ) ? ( n3055 ) : ( n37515 ) ;
assign n37517 =  ( n168 ) ? ( n3054 ) : ( n37516 ) ;
assign n37518 =  ( n166 ) ? ( n3053 ) : ( n37517 ) ;
assign n37519 =  ( n162 ) ? ( n3052 ) : ( n37518 ) ;
assign n37520 =  ( n3032 ) ? ( VREG_15_0 ) : ( n37519 ) ;
assign n37521 =  ( n3051 ) ? ( n37520 ) : ( VREG_15_0 ) ;
assign n37522 =  ( n3040 ) ? ( n37514 ) : ( n37521 ) ;
assign n37523 =  ( n192 ) ? ( VREG_15_0 ) : ( VREG_15_0 ) ;
assign n37524 =  ( n157 ) ? ( n37522 ) : ( n37523 ) ;
assign n37525 =  ( n6 ) ? ( n37509 ) : ( n37524 ) ;
assign n37526 =  ( n329 ) ? ( n37525 ) : ( VREG_15_0 ) ;
assign n37527 =  ( n148 ) ? ( n4113 ) : ( VREG_15_1 ) ;
assign n37528 =  ( n146 ) ? ( n4112 ) : ( n37527 ) ;
assign n37529 =  ( n144 ) ? ( n4111 ) : ( n37528 ) ;
assign n37530 =  ( n142 ) ? ( n4110 ) : ( n37529 ) ;
assign n37531 =  ( n10 ) ? ( n4109 ) : ( n37530 ) ;
assign n37532 =  ( n148 ) ? ( n5147 ) : ( VREG_15_1 ) ;
assign n37533 =  ( n146 ) ? ( n5146 ) : ( n37532 ) ;
assign n37534 =  ( n144 ) ? ( n5145 ) : ( n37533 ) ;
assign n37535 =  ( n142 ) ? ( n5144 ) : ( n37534 ) ;
assign n37536 =  ( n10 ) ? ( n5143 ) : ( n37535 ) ;
assign n37537 =  ( n5154 ) ? ( VREG_15_1 ) : ( n37531 ) ;
assign n37538 =  ( n5154 ) ? ( VREG_15_1 ) : ( n37536 ) ;
assign n37539 =  ( n3034 ) ? ( n37538 ) : ( VREG_15_1 ) ;
assign n37540 =  ( n2965 ) ? ( n37537 ) : ( n37539 ) ;
assign n37541 =  ( n1930 ) ? ( n37536 ) : ( n37540 ) ;
assign n37542 =  ( n879 ) ? ( n37531 ) : ( n37541 ) ;
assign n37543 =  ( n172 ) ? ( n5165 ) : ( VREG_15_1 ) ;
assign n37544 =  ( n170 ) ? ( n5164 ) : ( n37543 ) ;
assign n37545 =  ( n168 ) ? ( n5163 ) : ( n37544 ) ;
assign n37546 =  ( n166 ) ? ( n5162 ) : ( n37545 ) ;
assign n37547 =  ( n162 ) ? ( n5161 ) : ( n37546 ) ;
assign n37548 =  ( n172 ) ? ( n5175 ) : ( VREG_15_1 ) ;
assign n37549 =  ( n170 ) ? ( n5174 ) : ( n37548 ) ;
assign n37550 =  ( n168 ) ? ( n5173 ) : ( n37549 ) ;
assign n37551 =  ( n166 ) ? ( n5172 ) : ( n37550 ) ;
assign n37552 =  ( n162 ) ? ( n5171 ) : ( n37551 ) ;
assign n37553 =  ( n5154 ) ? ( VREG_15_1 ) : ( n37552 ) ;
assign n37554 =  ( n3051 ) ? ( n37553 ) : ( VREG_15_1 ) ;
assign n37555 =  ( n3040 ) ? ( n37547 ) : ( n37554 ) ;
assign n37556 =  ( n192 ) ? ( VREG_15_1 ) : ( VREG_15_1 ) ;
assign n37557 =  ( n157 ) ? ( n37555 ) : ( n37556 ) ;
assign n37558 =  ( n6 ) ? ( n37542 ) : ( n37557 ) ;
assign n37559 =  ( n329 ) ? ( n37558 ) : ( VREG_15_1 ) ;
assign n37560 =  ( n148 ) ? ( n6232 ) : ( VREG_15_10 ) ;
assign n37561 =  ( n146 ) ? ( n6231 ) : ( n37560 ) ;
assign n37562 =  ( n144 ) ? ( n6230 ) : ( n37561 ) ;
assign n37563 =  ( n142 ) ? ( n6229 ) : ( n37562 ) ;
assign n37564 =  ( n10 ) ? ( n6228 ) : ( n37563 ) ;
assign n37565 =  ( n148 ) ? ( n7266 ) : ( VREG_15_10 ) ;
assign n37566 =  ( n146 ) ? ( n7265 ) : ( n37565 ) ;
assign n37567 =  ( n144 ) ? ( n7264 ) : ( n37566 ) ;
assign n37568 =  ( n142 ) ? ( n7263 ) : ( n37567 ) ;
assign n37569 =  ( n10 ) ? ( n7262 ) : ( n37568 ) ;
assign n37570 =  ( n7273 ) ? ( VREG_15_10 ) : ( n37564 ) ;
assign n37571 =  ( n7273 ) ? ( VREG_15_10 ) : ( n37569 ) ;
assign n37572 =  ( n3034 ) ? ( n37571 ) : ( VREG_15_10 ) ;
assign n37573 =  ( n2965 ) ? ( n37570 ) : ( n37572 ) ;
assign n37574 =  ( n1930 ) ? ( n37569 ) : ( n37573 ) ;
assign n37575 =  ( n879 ) ? ( n37564 ) : ( n37574 ) ;
assign n37576 =  ( n172 ) ? ( n7284 ) : ( VREG_15_10 ) ;
assign n37577 =  ( n170 ) ? ( n7283 ) : ( n37576 ) ;
assign n37578 =  ( n168 ) ? ( n7282 ) : ( n37577 ) ;
assign n37579 =  ( n166 ) ? ( n7281 ) : ( n37578 ) ;
assign n37580 =  ( n162 ) ? ( n7280 ) : ( n37579 ) ;
assign n37581 =  ( n172 ) ? ( n7294 ) : ( VREG_15_10 ) ;
assign n37582 =  ( n170 ) ? ( n7293 ) : ( n37581 ) ;
assign n37583 =  ( n168 ) ? ( n7292 ) : ( n37582 ) ;
assign n37584 =  ( n166 ) ? ( n7291 ) : ( n37583 ) ;
assign n37585 =  ( n162 ) ? ( n7290 ) : ( n37584 ) ;
assign n37586 =  ( n7273 ) ? ( VREG_15_10 ) : ( n37585 ) ;
assign n37587 =  ( n3051 ) ? ( n37586 ) : ( VREG_15_10 ) ;
assign n37588 =  ( n3040 ) ? ( n37580 ) : ( n37587 ) ;
assign n37589 =  ( n192 ) ? ( VREG_15_10 ) : ( VREG_15_10 ) ;
assign n37590 =  ( n157 ) ? ( n37588 ) : ( n37589 ) ;
assign n37591 =  ( n6 ) ? ( n37575 ) : ( n37590 ) ;
assign n37592 =  ( n329 ) ? ( n37591 ) : ( VREG_15_10 ) ;
assign n37593 =  ( n148 ) ? ( n8351 ) : ( VREG_15_11 ) ;
assign n37594 =  ( n146 ) ? ( n8350 ) : ( n37593 ) ;
assign n37595 =  ( n144 ) ? ( n8349 ) : ( n37594 ) ;
assign n37596 =  ( n142 ) ? ( n8348 ) : ( n37595 ) ;
assign n37597 =  ( n10 ) ? ( n8347 ) : ( n37596 ) ;
assign n37598 =  ( n148 ) ? ( n9385 ) : ( VREG_15_11 ) ;
assign n37599 =  ( n146 ) ? ( n9384 ) : ( n37598 ) ;
assign n37600 =  ( n144 ) ? ( n9383 ) : ( n37599 ) ;
assign n37601 =  ( n142 ) ? ( n9382 ) : ( n37600 ) ;
assign n37602 =  ( n10 ) ? ( n9381 ) : ( n37601 ) ;
assign n37603 =  ( n9392 ) ? ( VREG_15_11 ) : ( n37597 ) ;
assign n37604 =  ( n9392 ) ? ( VREG_15_11 ) : ( n37602 ) ;
assign n37605 =  ( n3034 ) ? ( n37604 ) : ( VREG_15_11 ) ;
assign n37606 =  ( n2965 ) ? ( n37603 ) : ( n37605 ) ;
assign n37607 =  ( n1930 ) ? ( n37602 ) : ( n37606 ) ;
assign n37608 =  ( n879 ) ? ( n37597 ) : ( n37607 ) ;
assign n37609 =  ( n172 ) ? ( n9403 ) : ( VREG_15_11 ) ;
assign n37610 =  ( n170 ) ? ( n9402 ) : ( n37609 ) ;
assign n37611 =  ( n168 ) ? ( n9401 ) : ( n37610 ) ;
assign n37612 =  ( n166 ) ? ( n9400 ) : ( n37611 ) ;
assign n37613 =  ( n162 ) ? ( n9399 ) : ( n37612 ) ;
assign n37614 =  ( n172 ) ? ( n9413 ) : ( VREG_15_11 ) ;
assign n37615 =  ( n170 ) ? ( n9412 ) : ( n37614 ) ;
assign n37616 =  ( n168 ) ? ( n9411 ) : ( n37615 ) ;
assign n37617 =  ( n166 ) ? ( n9410 ) : ( n37616 ) ;
assign n37618 =  ( n162 ) ? ( n9409 ) : ( n37617 ) ;
assign n37619 =  ( n9392 ) ? ( VREG_15_11 ) : ( n37618 ) ;
assign n37620 =  ( n3051 ) ? ( n37619 ) : ( VREG_15_11 ) ;
assign n37621 =  ( n3040 ) ? ( n37613 ) : ( n37620 ) ;
assign n37622 =  ( n192 ) ? ( VREG_15_11 ) : ( VREG_15_11 ) ;
assign n37623 =  ( n157 ) ? ( n37621 ) : ( n37622 ) ;
assign n37624 =  ( n6 ) ? ( n37608 ) : ( n37623 ) ;
assign n37625 =  ( n329 ) ? ( n37624 ) : ( VREG_15_11 ) ;
assign n37626 =  ( n148 ) ? ( n10470 ) : ( VREG_15_12 ) ;
assign n37627 =  ( n146 ) ? ( n10469 ) : ( n37626 ) ;
assign n37628 =  ( n144 ) ? ( n10468 ) : ( n37627 ) ;
assign n37629 =  ( n142 ) ? ( n10467 ) : ( n37628 ) ;
assign n37630 =  ( n10 ) ? ( n10466 ) : ( n37629 ) ;
assign n37631 =  ( n148 ) ? ( n11504 ) : ( VREG_15_12 ) ;
assign n37632 =  ( n146 ) ? ( n11503 ) : ( n37631 ) ;
assign n37633 =  ( n144 ) ? ( n11502 ) : ( n37632 ) ;
assign n37634 =  ( n142 ) ? ( n11501 ) : ( n37633 ) ;
assign n37635 =  ( n10 ) ? ( n11500 ) : ( n37634 ) ;
assign n37636 =  ( n11511 ) ? ( VREG_15_12 ) : ( n37630 ) ;
assign n37637 =  ( n11511 ) ? ( VREG_15_12 ) : ( n37635 ) ;
assign n37638 =  ( n3034 ) ? ( n37637 ) : ( VREG_15_12 ) ;
assign n37639 =  ( n2965 ) ? ( n37636 ) : ( n37638 ) ;
assign n37640 =  ( n1930 ) ? ( n37635 ) : ( n37639 ) ;
assign n37641 =  ( n879 ) ? ( n37630 ) : ( n37640 ) ;
assign n37642 =  ( n172 ) ? ( n11522 ) : ( VREG_15_12 ) ;
assign n37643 =  ( n170 ) ? ( n11521 ) : ( n37642 ) ;
assign n37644 =  ( n168 ) ? ( n11520 ) : ( n37643 ) ;
assign n37645 =  ( n166 ) ? ( n11519 ) : ( n37644 ) ;
assign n37646 =  ( n162 ) ? ( n11518 ) : ( n37645 ) ;
assign n37647 =  ( n172 ) ? ( n11532 ) : ( VREG_15_12 ) ;
assign n37648 =  ( n170 ) ? ( n11531 ) : ( n37647 ) ;
assign n37649 =  ( n168 ) ? ( n11530 ) : ( n37648 ) ;
assign n37650 =  ( n166 ) ? ( n11529 ) : ( n37649 ) ;
assign n37651 =  ( n162 ) ? ( n11528 ) : ( n37650 ) ;
assign n37652 =  ( n11511 ) ? ( VREG_15_12 ) : ( n37651 ) ;
assign n37653 =  ( n3051 ) ? ( n37652 ) : ( VREG_15_12 ) ;
assign n37654 =  ( n3040 ) ? ( n37646 ) : ( n37653 ) ;
assign n37655 =  ( n192 ) ? ( VREG_15_12 ) : ( VREG_15_12 ) ;
assign n37656 =  ( n157 ) ? ( n37654 ) : ( n37655 ) ;
assign n37657 =  ( n6 ) ? ( n37641 ) : ( n37656 ) ;
assign n37658 =  ( n329 ) ? ( n37657 ) : ( VREG_15_12 ) ;
assign n37659 =  ( n148 ) ? ( n12589 ) : ( VREG_15_13 ) ;
assign n37660 =  ( n146 ) ? ( n12588 ) : ( n37659 ) ;
assign n37661 =  ( n144 ) ? ( n12587 ) : ( n37660 ) ;
assign n37662 =  ( n142 ) ? ( n12586 ) : ( n37661 ) ;
assign n37663 =  ( n10 ) ? ( n12585 ) : ( n37662 ) ;
assign n37664 =  ( n148 ) ? ( n13623 ) : ( VREG_15_13 ) ;
assign n37665 =  ( n146 ) ? ( n13622 ) : ( n37664 ) ;
assign n37666 =  ( n144 ) ? ( n13621 ) : ( n37665 ) ;
assign n37667 =  ( n142 ) ? ( n13620 ) : ( n37666 ) ;
assign n37668 =  ( n10 ) ? ( n13619 ) : ( n37667 ) ;
assign n37669 =  ( n13630 ) ? ( VREG_15_13 ) : ( n37663 ) ;
assign n37670 =  ( n13630 ) ? ( VREG_15_13 ) : ( n37668 ) ;
assign n37671 =  ( n3034 ) ? ( n37670 ) : ( VREG_15_13 ) ;
assign n37672 =  ( n2965 ) ? ( n37669 ) : ( n37671 ) ;
assign n37673 =  ( n1930 ) ? ( n37668 ) : ( n37672 ) ;
assign n37674 =  ( n879 ) ? ( n37663 ) : ( n37673 ) ;
assign n37675 =  ( n172 ) ? ( n13641 ) : ( VREG_15_13 ) ;
assign n37676 =  ( n170 ) ? ( n13640 ) : ( n37675 ) ;
assign n37677 =  ( n168 ) ? ( n13639 ) : ( n37676 ) ;
assign n37678 =  ( n166 ) ? ( n13638 ) : ( n37677 ) ;
assign n37679 =  ( n162 ) ? ( n13637 ) : ( n37678 ) ;
assign n37680 =  ( n172 ) ? ( n13651 ) : ( VREG_15_13 ) ;
assign n37681 =  ( n170 ) ? ( n13650 ) : ( n37680 ) ;
assign n37682 =  ( n168 ) ? ( n13649 ) : ( n37681 ) ;
assign n37683 =  ( n166 ) ? ( n13648 ) : ( n37682 ) ;
assign n37684 =  ( n162 ) ? ( n13647 ) : ( n37683 ) ;
assign n37685 =  ( n13630 ) ? ( VREG_15_13 ) : ( n37684 ) ;
assign n37686 =  ( n3051 ) ? ( n37685 ) : ( VREG_15_13 ) ;
assign n37687 =  ( n3040 ) ? ( n37679 ) : ( n37686 ) ;
assign n37688 =  ( n192 ) ? ( VREG_15_13 ) : ( VREG_15_13 ) ;
assign n37689 =  ( n157 ) ? ( n37687 ) : ( n37688 ) ;
assign n37690 =  ( n6 ) ? ( n37674 ) : ( n37689 ) ;
assign n37691 =  ( n329 ) ? ( n37690 ) : ( VREG_15_13 ) ;
assign n37692 =  ( n148 ) ? ( n14708 ) : ( VREG_15_14 ) ;
assign n37693 =  ( n146 ) ? ( n14707 ) : ( n37692 ) ;
assign n37694 =  ( n144 ) ? ( n14706 ) : ( n37693 ) ;
assign n37695 =  ( n142 ) ? ( n14705 ) : ( n37694 ) ;
assign n37696 =  ( n10 ) ? ( n14704 ) : ( n37695 ) ;
assign n37697 =  ( n148 ) ? ( n15742 ) : ( VREG_15_14 ) ;
assign n37698 =  ( n146 ) ? ( n15741 ) : ( n37697 ) ;
assign n37699 =  ( n144 ) ? ( n15740 ) : ( n37698 ) ;
assign n37700 =  ( n142 ) ? ( n15739 ) : ( n37699 ) ;
assign n37701 =  ( n10 ) ? ( n15738 ) : ( n37700 ) ;
assign n37702 =  ( n15749 ) ? ( VREG_15_14 ) : ( n37696 ) ;
assign n37703 =  ( n15749 ) ? ( VREG_15_14 ) : ( n37701 ) ;
assign n37704 =  ( n3034 ) ? ( n37703 ) : ( VREG_15_14 ) ;
assign n37705 =  ( n2965 ) ? ( n37702 ) : ( n37704 ) ;
assign n37706 =  ( n1930 ) ? ( n37701 ) : ( n37705 ) ;
assign n37707 =  ( n879 ) ? ( n37696 ) : ( n37706 ) ;
assign n37708 =  ( n172 ) ? ( n15760 ) : ( VREG_15_14 ) ;
assign n37709 =  ( n170 ) ? ( n15759 ) : ( n37708 ) ;
assign n37710 =  ( n168 ) ? ( n15758 ) : ( n37709 ) ;
assign n37711 =  ( n166 ) ? ( n15757 ) : ( n37710 ) ;
assign n37712 =  ( n162 ) ? ( n15756 ) : ( n37711 ) ;
assign n37713 =  ( n172 ) ? ( n15770 ) : ( VREG_15_14 ) ;
assign n37714 =  ( n170 ) ? ( n15769 ) : ( n37713 ) ;
assign n37715 =  ( n168 ) ? ( n15768 ) : ( n37714 ) ;
assign n37716 =  ( n166 ) ? ( n15767 ) : ( n37715 ) ;
assign n37717 =  ( n162 ) ? ( n15766 ) : ( n37716 ) ;
assign n37718 =  ( n15749 ) ? ( VREG_15_14 ) : ( n37717 ) ;
assign n37719 =  ( n3051 ) ? ( n37718 ) : ( VREG_15_14 ) ;
assign n37720 =  ( n3040 ) ? ( n37712 ) : ( n37719 ) ;
assign n37721 =  ( n192 ) ? ( VREG_15_14 ) : ( VREG_15_14 ) ;
assign n37722 =  ( n157 ) ? ( n37720 ) : ( n37721 ) ;
assign n37723 =  ( n6 ) ? ( n37707 ) : ( n37722 ) ;
assign n37724 =  ( n329 ) ? ( n37723 ) : ( VREG_15_14 ) ;
assign n37725 =  ( n148 ) ? ( n16827 ) : ( VREG_15_15 ) ;
assign n37726 =  ( n146 ) ? ( n16826 ) : ( n37725 ) ;
assign n37727 =  ( n144 ) ? ( n16825 ) : ( n37726 ) ;
assign n37728 =  ( n142 ) ? ( n16824 ) : ( n37727 ) ;
assign n37729 =  ( n10 ) ? ( n16823 ) : ( n37728 ) ;
assign n37730 =  ( n148 ) ? ( n17861 ) : ( VREG_15_15 ) ;
assign n37731 =  ( n146 ) ? ( n17860 ) : ( n37730 ) ;
assign n37732 =  ( n144 ) ? ( n17859 ) : ( n37731 ) ;
assign n37733 =  ( n142 ) ? ( n17858 ) : ( n37732 ) ;
assign n37734 =  ( n10 ) ? ( n17857 ) : ( n37733 ) ;
assign n37735 =  ( n17868 ) ? ( VREG_15_15 ) : ( n37729 ) ;
assign n37736 =  ( n17868 ) ? ( VREG_15_15 ) : ( n37734 ) ;
assign n37737 =  ( n3034 ) ? ( n37736 ) : ( VREG_15_15 ) ;
assign n37738 =  ( n2965 ) ? ( n37735 ) : ( n37737 ) ;
assign n37739 =  ( n1930 ) ? ( n37734 ) : ( n37738 ) ;
assign n37740 =  ( n879 ) ? ( n37729 ) : ( n37739 ) ;
assign n37741 =  ( n172 ) ? ( n17879 ) : ( VREG_15_15 ) ;
assign n37742 =  ( n170 ) ? ( n17878 ) : ( n37741 ) ;
assign n37743 =  ( n168 ) ? ( n17877 ) : ( n37742 ) ;
assign n37744 =  ( n166 ) ? ( n17876 ) : ( n37743 ) ;
assign n37745 =  ( n162 ) ? ( n17875 ) : ( n37744 ) ;
assign n37746 =  ( n172 ) ? ( n17889 ) : ( VREG_15_15 ) ;
assign n37747 =  ( n170 ) ? ( n17888 ) : ( n37746 ) ;
assign n37748 =  ( n168 ) ? ( n17887 ) : ( n37747 ) ;
assign n37749 =  ( n166 ) ? ( n17886 ) : ( n37748 ) ;
assign n37750 =  ( n162 ) ? ( n17885 ) : ( n37749 ) ;
assign n37751 =  ( n17868 ) ? ( VREG_15_15 ) : ( n37750 ) ;
assign n37752 =  ( n3051 ) ? ( n37751 ) : ( VREG_15_15 ) ;
assign n37753 =  ( n3040 ) ? ( n37745 ) : ( n37752 ) ;
assign n37754 =  ( n192 ) ? ( VREG_15_15 ) : ( VREG_15_15 ) ;
assign n37755 =  ( n157 ) ? ( n37753 ) : ( n37754 ) ;
assign n37756 =  ( n6 ) ? ( n37740 ) : ( n37755 ) ;
assign n37757 =  ( n329 ) ? ( n37756 ) : ( VREG_15_15 ) ;
assign n37758 =  ( n148 ) ? ( n18946 ) : ( VREG_15_2 ) ;
assign n37759 =  ( n146 ) ? ( n18945 ) : ( n37758 ) ;
assign n37760 =  ( n144 ) ? ( n18944 ) : ( n37759 ) ;
assign n37761 =  ( n142 ) ? ( n18943 ) : ( n37760 ) ;
assign n37762 =  ( n10 ) ? ( n18942 ) : ( n37761 ) ;
assign n37763 =  ( n148 ) ? ( n19980 ) : ( VREG_15_2 ) ;
assign n37764 =  ( n146 ) ? ( n19979 ) : ( n37763 ) ;
assign n37765 =  ( n144 ) ? ( n19978 ) : ( n37764 ) ;
assign n37766 =  ( n142 ) ? ( n19977 ) : ( n37765 ) ;
assign n37767 =  ( n10 ) ? ( n19976 ) : ( n37766 ) ;
assign n37768 =  ( n19987 ) ? ( VREG_15_2 ) : ( n37762 ) ;
assign n37769 =  ( n19987 ) ? ( VREG_15_2 ) : ( n37767 ) ;
assign n37770 =  ( n3034 ) ? ( n37769 ) : ( VREG_15_2 ) ;
assign n37771 =  ( n2965 ) ? ( n37768 ) : ( n37770 ) ;
assign n37772 =  ( n1930 ) ? ( n37767 ) : ( n37771 ) ;
assign n37773 =  ( n879 ) ? ( n37762 ) : ( n37772 ) ;
assign n37774 =  ( n172 ) ? ( n19998 ) : ( VREG_15_2 ) ;
assign n37775 =  ( n170 ) ? ( n19997 ) : ( n37774 ) ;
assign n37776 =  ( n168 ) ? ( n19996 ) : ( n37775 ) ;
assign n37777 =  ( n166 ) ? ( n19995 ) : ( n37776 ) ;
assign n37778 =  ( n162 ) ? ( n19994 ) : ( n37777 ) ;
assign n37779 =  ( n172 ) ? ( n20008 ) : ( VREG_15_2 ) ;
assign n37780 =  ( n170 ) ? ( n20007 ) : ( n37779 ) ;
assign n37781 =  ( n168 ) ? ( n20006 ) : ( n37780 ) ;
assign n37782 =  ( n166 ) ? ( n20005 ) : ( n37781 ) ;
assign n37783 =  ( n162 ) ? ( n20004 ) : ( n37782 ) ;
assign n37784 =  ( n19987 ) ? ( VREG_15_2 ) : ( n37783 ) ;
assign n37785 =  ( n3051 ) ? ( n37784 ) : ( VREG_15_2 ) ;
assign n37786 =  ( n3040 ) ? ( n37778 ) : ( n37785 ) ;
assign n37787 =  ( n192 ) ? ( VREG_15_2 ) : ( VREG_15_2 ) ;
assign n37788 =  ( n157 ) ? ( n37786 ) : ( n37787 ) ;
assign n37789 =  ( n6 ) ? ( n37773 ) : ( n37788 ) ;
assign n37790 =  ( n329 ) ? ( n37789 ) : ( VREG_15_2 ) ;
assign n37791 =  ( n148 ) ? ( n21065 ) : ( VREG_15_3 ) ;
assign n37792 =  ( n146 ) ? ( n21064 ) : ( n37791 ) ;
assign n37793 =  ( n144 ) ? ( n21063 ) : ( n37792 ) ;
assign n37794 =  ( n142 ) ? ( n21062 ) : ( n37793 ) ;
assign n37795 =  ( n10 ) ? ( n21061 ) : ( n37794 ) ;
assign n37796 =  ( n148 ) ? ( n22099 ) : ( VREG_15_3 ) ;
assign n37797 =  ( n146 ) ? ( n22098 ) : ( n37796 ) ;
assign n37798 =  ( n144 ) ? ( n22097 ) : ( n37797 ) ;
assign n37799 =  ( n142 ) ? ( n22096 ) : ( n37798 ) ;
assign n37800 =  ( n10 ) ? ( n22095 ) : ( n37799 ) ;
assign n37801 =  ( n22106 ) ? ( VREG_15_3 ) : ( n37795 ) ;
assign n37802 =  ( n22106 ) ? ( VREG_15_3 ) : ( n37800 ) ;
assign n37803 =  ( n3034 ) ? ( n37802 ) : ( VREG_15_3 ) ;
assign n37804 =  ( n2965 ) ? ( n37801 ) : ( n37803 ) ;
assign n37805 =  ( n1930 ) ? ( n37800 ) : ( n37804 ) ;
assign n37806 =  ( n879 ) ? ( n37795 ) : ( n37805 ) ;
assign n37807 =  ( n172 ) ? ( n22117 ) : ( VREG_15_3 ) ;
assign n37808 =  ( n170 ) ? ( n22116 ) : ( n37807 ) ;
assign n37809 =  ( n168 ) ? ( n22115 ) : ( n37808 ) ;
assign n37810 =  ( n166 ) ? ( n22114 ) : ( n37809 ) ;
assign n37811 =  ( n162 ) ? ( n22113 ) : ( n37810 ) ;
assign n37812 =  ( n172 ) ? ( n22127 ) : ( VREG_15_3 ) ;
assign n37813 =  ( n170 ) ? ( n22126 ) : ( n37812 ) ;
assign n37814 =  ( n168 ) ? ( n22125 ) : ( n37813 ) ;
assign n37815 =  ( n166 ) ? ( n22124 ) : ( n37814 ) ;
assign n37816 =  ( n162 ) ? ( n22123 ) : ( n37815 ) ;
assign n37817 =  ( n22106 ) ? ( VREG_15_3 ) : ( n37816 ) ;
assign n37818 =  ( n3051 ) ? ( n37817 ) : ( VREG_15_3 ) ;
assign n37819 =  ( n3040 ) ? ( n37811 ) : ( n37818 ) ;
assign n37820 =  ( n192 ) ? ( VREG_15_3 ) : ( VREG_15_3 ) ;
assign n37821 =  ( n157 ) ? ( n37819 ) : ( n37820 ) ;
assign n37822 =  ( n6 ) ? ( n37806 ) : ( n37821 ) ;
assign n37823 =  ( n329 ) ? ( n37822 ) : ( VREG_15_3 ) ;
assign n37824 =  ( n148 ) ? ( n23184 ) : ( VREG_15_4 ) ;
assign n37825 =  ( n146 ) ? ( n23183 ) : ( n37824 ) ;
assign n37826 =  ( n144 ) ? ( n23182 ) : ( n37825 ) ;
assign n37827 =  ( n142 ) ? ( n23181 ) : ( n37826 ) ;
assign n37828 =  ( n10 ) ? ( n23180 ) : ( n37827 ) ;
assign n37829 =  ( n148 ) ? ( n24218 ) : ( VREG_15_4 ) ;
assign n37830 =  ( n146 ) ? ( n24217 ) : ( n37829 ) ;
assign n37831 =  ( n144 ) ? ( n24216 ) : ( n37830 ) ;
assign n37832 =  ( n142 ) ? ( n24215 ) : ( n37831 ) ;
assign n37833 =  ( n10 ) ? ( n24214 ) : ( n37832 ) ;
assign n37834 =  ( n24225 ) ? ( VREG_15_4 ) : ( n37828 ) ;
assign n37835 =  ( n24225 ) ? ( VREG_15_4 ) : ( n37833 ) ;
assign n37836 =  ( n3034 ) ? ( n37835 ) : ( VREG_15_4 ) ;
assign n37837 =  ( n2965 ) ? ( n37834 ) : ( n37836 ) ;
assign n37838 =  ( n1930 ) ? ( n37833 ) : ( n37837 ) ;
assign n37839 =  ( n879 ) ? ( n37828 ) : ( n37838 ) ;
assign n37840 =  ( n172 ) ? ( n24236 ) : ( VREG_15_4 ) ;
assign n37841 =  ( n170 ) ? ( n24235 ) : ( n37840 ) ;
assign n37842 =  ( n168 ) ? ( n24234 ) : ( n37841 ) ;
assign n37843 =  ( n166 ) ? ( n24233 ) : ( n37842 ) ;
assign n37844 =  ( n162 ) ? ( n24232 ) : ( n37843 ) ;
assign n37845 =  ( n172 ) ? ( n24246 ) : ( VREG_15_4 ) ;
assign n37846 =  ( n170 ) ? ( n24245 ) : ( n37845 ) ;
assign n37847 =  ( n168 ) ? ( n24244 ) : ( n37846 ) ;
assign n37848 =  ( n166 ) ? ( n24243 ) : ( n37847 ) ;
assign n37849 =  ( n162 ) ? ( n24242 ) : ( n37848 ) ;
assign n37850 =  ( n24225 ) ? ( VREG_15_4 ) : ( n37849 ) ;
assign n37851 =  ( n3051 ) ? ( n37850 ) : ( VREG_15_4 ) ;
assign n37852 =  ( n3040 ) ? ( n37844 ) : ( n37851 ) ;
assign n37853 =  ( n192 ) ? ( VREG_15_4 ) : ( VREG_15_4 ) ;
assign n37854 =  ( n157 ) ? ( n37852 ) : ( n37853 ) ;
assign n37855 =  ( n6 ) ? ( n37839 ) : ( n37854 ) ;
assign n37856 =  ( n329 ) ? ( n37855 ) : ( VREG_15_4 ) ;
assign n37857 =  ( n148 ) ? ( n25303 ) : ( VREG_15_5 ) ;
assign n37858 =  ( n146 ) ? ( n25302 ) : ( n37857 ) ;
assign n37859 =  ( n144 ) ? ( n25301 ) : ( n37858 ) ;
assign n37860 =  ( n142 ) ? ( n25300 ) : ( n37859 ) ;
assign n37861 =  ( n10 ) ? ( n25299 ) : ( n37860 ) ;
assign n37862 =  ( n148 ) ? ( n26337 ) : ( VREG_15_5 ) ;
assign n37863 =  ( n146 ) ? ( n26336 ) : ( n37862 ) ;
assign n37864 =  ( n144 ) ? ( n26335 ) : ( n37863 ) ;
assign n37865 =  ( n142 ) ? ( n26334 ) : ( n37864 ) ;
assign n37866 =  ( n10 ) ? ( n26333 ) : ( n37865 ) ;
assign n37867 =  ( n26344 ) ? ( VREG_15_5 ) : ( n37861 ) ;
assign n37868 =  ( n26344 ) ? ( VREG_15_5 ) : ( n37866 ) ;
assign n37869 =  ( n3034 ) ? ( n37868 ) : ( VREG_15_5 ) ;
assign n37870 =  ( n2965 ) ? ( n37867 ) : ( n37869 ) ;
assign n37871 =  ( n1930 ) ? ( n37866 ) : ( n37870 ) ;
assign n37872 =  ( n879 ) ? ( n37861 ) : ( n37871 ) ;
assign n37873 =  ( n172 ) ? ( n26355 ) : ( VREG_15_5 ) ;
assign n37874 =  ( n170 ) ? ( n26354 ) : ( n37873 ) ;
assign n37875 =  ( n168 ) ? ( n26353 ) : ( n37874 ) ;
assign n37876 =  ( n166 ) ? ( n26352 ) : ( n37875 ) ;
assign n37877 =  ( n162 ) ? ( n26351 ) : ( n37876 ) ;
assign n37878 =  ( n172 ) ? ( n26365 ) : ( VREG_15_5 ) ;
assign n37879 =  ( n170 ) ? ( n26364 ) : ( n37878 ) ;
assign n37880 =  ( n168 ) ? ( n26363 ) : ( n37879 ) ;
assign n37881 =  ( n166 ) ? ( n26362 ) : ( n37880 ) ;
assign n37882 =  ( n162 ) ? ( n26361 ) : ( n37881 ) ;
assign n37883 =  ( n26344 ) ? ( VREG_15_5 ) : ( n37882 ) ;
assign n37884 =  ( n3051 ) ? ( n37883 ) : ( VREG_15_5 ) ;
assign n37885 =  ( n3040 ) ? ( n37877 ) : ( n37884 ) ;
assign n37886 =  ( n192 ) ? ( VREG_15_5 ) : ( VREG_15_5 ) ;
assign n37887 =  ( n157 ) ? ( n37885 ) : ( n37886 ) ;
assign n37888 =  ( n6 ) ? ( n37872 ) : ( n37887 ) ;
assign n37889 =  ( n329 ) ? ( n37888 ) : ( VREG_15_5 ) ;
assign n37890 =  ( n148 ) ? ( n27422 ) : ( VREG_15_6 ) ;
assign n37891 =  ( n146 ) ? ( n27421 ) : ( n37890 ) ;
assign n37892 =  ( n144 ) ? ( n27420 ) : ( n37891 ) ;
assign n37893 =  ( n142 ) ? ( n27419 ) : ( n37892 ) ;
assign n37894 =  ( n10 ) ? ( n27418 ) : ( n37893 ) ;
assign n37895 =  ( n148 ) ? ( n28456 ) : ( VREG_15_6 ) ;
assign n37896 =  ( n146 ) ? ( n28455 ) : ( n37895 ) ;
assign n37897 =  ( n144 ) ? ( n28454 ) : ( n37896 ) ;
assign n37898 =  ( n142 ) ? ( n28453 ) : ( n37897 ) ;
assign n37899 =  ( n10 ) ? ( n28452 ) : ( n37898 ) ;
assign n37900 =  ( n28463 ) ? ( VREG_15_6 ) : ( n37894 ) ;
assign n37901 =  ( n28463 ) ? ( VREG_15_6 ) : ( n37899 ) ;
assign n37902 =  ( n3034 ) ? ( n37901 ) : ( VREG_15_6 ) ;
assign n37903 =  ( n2965 ) ? ( n37900 ) : ( n37902 ) ;
assign n37904 =  ( n1930 ) ? ( n37899 ) : ( n37903 ) ;
assign n37905 =  ( n879 ) ? ( n37894 ) : ( n37904 ) ;
assign n37906 =  ( n172 ) ? ( n28474 ) : ( VREG_15_6 ) ;
assign n37907 =  ( n170 ) ? ( n28473 ) : ( n37906 ) ;
assign n37908 =  ( n168 ) ? ( n28472 ) : ( n37907 ) ;
assign n37909 =  ( n166 ) ? ( n28471 ) : ( n37908 ) ;
assign n37910 =  ( n162 ) ? ( n28470 ) : ( n37909 ) ;
assign n37911 =  ( n172 ) ? ( n28484 ) : ( VREG_15_6 ) ;
assign n37912 =  ( n170 ) ? ( n28483 ) : ( n37911 ) ;
assign n37913 =  ( n168 ) ? ( n28482 ) : ( n37912 ) ;
assign n37914 =  ( n166 ) ? ( n28481 ) : ( n37913 ) ;
assign n37915 =  ( n162 ) ? ( n28480 ) : ( n37914 ) ;
assign n37916 =  ( n28463 ) ? ( VREG_15_6 ) : ( n37915 ) ;
assign n37917 =  ( n3051 ) ? ( n37916 ) : ( VREG_15_6 ) ;
assign n37918 =  ( n3040 ) ? ( n37910 ) : ( n37917 ) ;
assign n37919 =  ( n192 ) ? ( VREG_15_6 ) : ( VREG_15_6 ) ;
assign n37920 =  ( n157 ) ? ( n37918 ) : ( n37919 ) ;
assign n37921 =  ( n6 ) ? ( n37905 ) : ( n37920 ) ;
assign n37922 =  ( n329 ) ? ( n37921 ) : ( VREG_15_6 ) ;
assign n37923 =  ( n148 ) ? ( n29541 ) : ( VREG_15_7 ) ;
assign n37924 =  ( n146 ) ? ( n29540 ) : ( n37923 ) ;
assign n37925 =  ( n144 ) ? ( n29539 ) : ( n37924 ) ;
assign n37926 =  ( n142 ) ? ( n29538 ) : ( n37925 ) ;
assign n37927 =  ( n10 ) ? ( n29537 ) : ( n37926 ) ;
assign n37928 =  ( n148 ) ? ( n30575 ) : ( VREG_15_7 ) ;
assign n37929 =  ( n146 ) ? ( n30574 ) : ( n37928 ) ;
assign n37930 =  ( n144 ) ? ( n30573 ) : ( n37929 ) ;
assign n37931 =  ( n142 ) ? ( n30572 ) : ( n37930 ) ;
assign n37932 =  ( n10 ) ? ( n30571 ) : ( n37931 ) ;
assign n37933 =  ( n30582 ) ? ( VREG_15_7 ) : ( n37927 ) ;
assign n37934 =  ( n30582 ) ? ( VREG_15_7 ) : ( n37932 ) ;
assign n37935 =  ( n3034 ) ? ( n37934 ) : ( VREG_15_7 ) ;
assign n37936 =  ( n2965 ) ? ( n37933 ) : ( n37935 ) ;
assign n37937 =  ( n1930 ) ? ( n37932 ) : ( n37936 ) ;
assign n37938 =  ( n879 ) ? ( n37927 ) : ( n37937 ) ;
assign n37939 =  ( n172 ) ? ( n30593 ) : ( VREG_15_7 ) ;
assign n37940 =  ( n170 ) ? ( n30592 ) : ( n37939 ) ;
assign n37941 =  ( n168 ) ? ( n30591 ) : ( n37940 ) ;
assign n37942 =  ( n166 ) ? ( n30590 ) : ( n37941 ) ;
assign n37943 =  ( n162 ) ? ( n30589 ) : ( n37942 ) ;
assign n37944 =  ( n172 ) ? ( n30603 ) : ( VREG_15_7 ) ;
assign n37945 =  ( n170 ) ? ( n30602 ) : ( n37944 ) ;
assign n37946 =  ( n168 ) ? ( n30601 ) : ( n37945 ) ;
assign n37947 =  ( n166 ) ? ( n30600 ) : ( n37946 ) ;
assign n37948 =  ( n162 ) ? ( n30599 ) : ( n37947 ) ;
assign n37949 =  ( n30582 ) ? ( VREG_15_7 ) : ( n37948 ) ;
assign n37950 =  ( n3051 ) ? ( n37949 ) : ( VREG_15_7 ) ;
assign n37951 =  ( n3040 ) ? ( n37943 ) : ( n37950 ) ;
assign n37952 =  ( n192 ) ? ( VREG_15_7 ) : ( VREG_15_7 ) ;
assign n37953 =  ( n157 ) ? ( n37951 ) : ( n37952 ) ;
assign n37954 =  ( n6 ) ? ( n37938 ) : ( n37953 ) ;
assign n37955 =  ( n329 ) ? ( n37954 ) : ( VREG_15_7 ) ;
assign n37956 =  ( n148 ) ? ( n31660 ) : ( VREG_15_8 ) ;
assign n37957 =  ( n146 ) ? ( n31659 ) : ( n37956 ) ;
assign n37958 =  ( n144 ) ? ( n31658 ) : ( n37957 ) ;
assign n37959 =  ( n142 ) ? ( n31657 ) : ( n37958 ) ;
assign n37960 =  ( n10 ) ? ( n31656 ) : ( n37959 ) ;
assign n37961 =  ( n148 ) ? ( n32694 ) : ( VREG_15_8 ) ;
assign n37962 =  ( n146 ) ? ( n32693 ) : ( n37961 ) ;
assign n37963 =  ( n144 ) ? ( n32692 ) : ( n37962 ) ;
assign n37964 =  ( n142 ) ? ( n32691 ) : ( n37963 ) ;
assign n37965 =  ( n10 ) ? ( n32690 ) : ( n37964 ) ;
assign n37966 =  ( n32701 ) ? ( VREG_15_8 ) : ( n37960 ) ;
assign n37967 =  ( n32701 ) ? ( VREG_15_8 ) : ( n37965 ) ;
assign n37968 =  ( n3034 ) ? ( n37967 ) : ( VREG_15_8 ) ;
assign n37969 =  ( n2965 ) ? ( n37966 ) : ( n37968 ) ;
assign n37970 =  ( n1930 ) ? ( n37965 ) : ( n37969 ) ;
assign n37971 =  ( n879 ) ? ( n37960 ) : ( n37970 ) ;
assign n37972 =  ( n172 ) ? ( n32712 ) : ( VREG_15_8 ) ;
assign n37973 =  ( n170 ) ? ( n32711 ) : ( n37972 ) ;
assign n37974 =  ( n168 ) ? ( n32710 ) : ( n37973 ) ;
assign n37975 =  ( n166 ) ? ( n32709 ) : ( n37974 ) ;
assign n37976 =  ( n162 ) ? ( n32708 ) : ( n37975 ) ;
assign n37977 =  ( n172 ) ? ( n32722 ) : ( VREG_15_8 ) ;
assign n37978 =  ( n170 ) ? ( n32721 ) : ( n37977 ) ;
assign n37979 =  ( n168 ) ? ( n32720 ) : ( n37978 ) ;
assign n37980 =  ( n166 ) ? ( n32719 ) : ( n37979 ) ;
assign n37981 =  ( n162 ) ? ( n32718 ) : ( n37980 ) ;
assign n37982 =  ( n32701 ) ? ( VREG_15_8 ) : ( n37981 ) ;
assign n37983 =  ( n3051 ) ? ( n37982 ) : ( VREG_15_8 ) ;
assign n37984 =  ( n3040 ) ? ( n37976 ) : ( n37983 ) ;
assign n37985 =  ( n192 ) ? ( VREG_15_8 ) : ( VREG_15_8 ) ;
assign n37986 =  ( n157 ) ? ( n37984 ) : ( n37985 ) ;
assign n37987 =  ( n6 ) ? ( n37971 ) : ( n37986 ) ;
assign n37988 =  ( n329 ) ? ( n37987 ) : ( VREG_15_8 ) ;
assign n37989 =  ( n148 ) ? ( n33779 ) : ( VREG_15_9 ) ;
assign n37990 =  ( n146 ) ? ( n33778 ) : ( n37989 ) ;
assign n37991 =  ( n144 ) ? ( n33777 ) : ( n37990 ) ;
assign n37992 =  ( n142 ) ? ( n33776 ) : ( n37991 ) ;
assign n37993 =  ( n10 ) ? ( n33775 ) : ( n37992 ) ;
assign n37994 =  ( n148 ) ? ( n34813 ) : ( VREG_15_9 ) ;
assign n37995 =  ( n146 ) ? ( n34812 ) : ( n37994 ) ;
assign n37996 =  ( n144 ) ? ( n34811 ) : ( n37995 ) ;
assign n37997 =  ( n142 ) ? ( n34810 ) : ( n37996 ) ;
assign n37998 =  ( n10 ) ? ( n34809 ) : ( n37997 ) ;
assign n37999 =  ( n34820 ) ? ( VREG_15_9 ) : ( n37993 ) ;
assign n38000 =  ( n34820 ) ? ( VREG_15_9 ) : ( n37998 ) ;
assign n38001 =  ( n3034 ) ? ( n38000 ) : ( VREG_15_9 ) ;
assign n38002 =  ( n2965 ) ? ( n37999 ) : ( n38001 ) ;
assign n38003 =  ( n1930 ) ? ( n37998 ) : ( n38002 ) ;
assign n38004 =  ( n879 ) ? ( n37993 ) : ( n38003 ) ;
assign n38005 =  ( n172 ) ? ( n34831 ) : ( VREG_15_9 ) ;
assign n38006 =  ( n170 ) ? ( n34830 ) : ( n38005 ) ;
assign n38007 =  ( n168 ) ? ( n34829 ) : ( n38006 ) ;
assign n38008 =  ( n166 ) ? ( n34828 ) : ( n38007 ) ;
assign n38009 =  ( n162 ) ? ( n34827 ) : ( n38008 ) ;
assign n38010 =  ( n172 ) ? ( n34841 ) : ( VREG_15_9 ) ;
assign n38011 =  ( n170 ) ? ( n34840 ) : ( n38010 ) ;
assign n38012 =  ( n168 ) ? ( n34839 ) : ( n38011 ) ;
assign n38013 =  ( n166 ) ? ( n34838 ) : ( n38012 ) ;
assign n38014 =  ( n162 ) ? ( n34837 ) : ( n38013 ) ;
assign n38015 =  ( n34820 ) ? ( VREG_15_9 ) : ( n38014 ) ;
assign n38016 =  ( n3051 ) ? ( n38015 ) : ( VREG_15_9 ) ;
assign n38017 =  ( n3040 ) ? ( n38009 ) : ( n38016 ) ;
assign n38018 =  ( n192 ) ? ( VREG_15_9 ) : ( VREG_15_9 ) ;
assign n38019 =  ( n157 ) ? ( n38017 ) : ( n38018 ) ;
assign n38020 =  ( n6 ) ? ( n38004 ) : ( n38019 ) ;
assign n38021 =  ( n329 ) ? ( n38020 ) : ( VREG_15_9 ) ;
assign n38022 =  ( n148 ) ? ( n1924 ) : ( VREG_16_0 ) ;
assign n38023 =  ( n146 ) ? ( n1923 ) : ( n38022 ) ;
assign n38024 =  ( n144 ) ? ( n1922 ) : ( n38023 ) ;
assign n38025 =  ( n142 ) ? ( n1921 ) : ( n38024 ) ;
assign n38026 =  ( n10 ) ? ( n1920 ) : ( n38025 ) ;
assign n38027 =  ( n148 ) ? ( n2959 ) : ( VREG_16_0 ) ;
assign n38028 =  ( n146 ) ? ( n2958 ) : ( n38027 ) ;
assign n38029 =  ( n144 ) ? ( n2957 ) : ( n38028 ) ;
assign n38030 =  ( n142 ) ? ( n2956 ) : ( n38029 ) ;
assign n38031 =  ( n10 ) ? ( n2955 ) : ( n38030 ) ;
assign n38032 =  ( n3032 ) ? ( VREG_16_0 ) : ( n38026 ) ;
assign n38033 =  ( n3032 ) ? ( VREG_16_0 ) : ( n38031 ) ;
assign n38034 =  ( n3034 ) ? ( n38033 ) : ( VREG_16_0 ) ;
assign n38035 =  ( n2965 ) ? ( n38032 ) : ( n38034 ) ;
assign n38036 =  ( n1930 ) ? ( n38031 ) : ( n38035 ) ;
assign n38037 =  ( n879 ) ? ( n38026 ) : ( n38036 ) ;
assign n38038 =  ( n172 ) ? ( n3045 ) : ( VREG_16_0 ) ;
assign n38039 =  ( n170 ) ? ( n3044 ) : ( n38038 ) ;
assign n38040 =  ( n168 ) ? ( n3043 ) : ( n38039 ) ;
assign n38041 =  ( n166 ) ? ( n3042 ) : ( n38040 ) ;
assign n38042 =  ( n162 ) ? ( n3041 ) : ( n38041 ) ;
assign n38043 =  ( n172 ) ? ( n3056 ) : ( VREG_16_0 ) ;
assign n38044 =  ( n170 ) ? ( n3055 ) : ( n38043 ) ;
assign n38045 =  ( n168 ) ? ( n3054 ) : ( n38044 ) ;
assign n38046 =  ( n166 ) ? ( n3053 ) : ( n38045 ) ;
assign n38047 =  ( n162 ) ? ( n3052 ) : ( n38046 ) ;
assign n38048 =  ( n3032 ) ? ( VREG_16_0 ) : ( n38047 ) ;
assign n38049 =  ( n3051 ) ? ( n38048 ) : ( VREG_16_0 ) ;
assign n38050 =  ( n3040 ) ? ( n38042 ) : ( n38049 ) ;
assign n38051 =  ( n192 ) ? ( VREG_16_0 ) : ( VREG_16_0 ) ;
assign n38052 =  ( n157 ) ? ( n38050 ) : ( n38051 ) ;
assign n38053 =  ( n6 ) ? ( n38037 ) : ( n38052 ) ;
assign n38054 =  ( n351 ) ? ( n38053 ) : ( VREG_16_0 ) ;
assign n38055 =  ( n148 ) ? ( n4113 ) : ( VREG_16_1 ) ;
assign n38056 =  ( n146 ) ? ( n4112 ) : ( n38055 ) ;
assign n38057 =  ( n144 ) ? ( n4111 ) : ( n38056 ) ;
assign n38058 =  ( n142 ) ? ( n4110 ) : ( n38057 ) ;
assign n38059 =  ( n10 ) ? ( n4109 ) : ( n38058 ) ;
assign n38060 =  ( n148 ) ? ( n5147 ) : ( VREG_16_1 ) ;
assign n38061 =  ( n146 ) ? ( n5146 ) : ( n38060 ) ;
assign n38062 =  ( n144 ) ? ( n5145 ) : ( n38061 ) ;
assign n38063 =  ( n142 ) ? ( n5144 ) : ( n38062 ) ;
assign n38064 =  ( n10 ) ? ( n5143 ) : ( n38063 ) ;
assign n38065 =  ( n5154 ) ? ( VREG_16_1 ) : ( n38059 ) ;
assign n38066 =  ( n5154 ) ? ( VREG_16_1 ) : ( n38064 ) ;
assign n38067 =  ( n3034 ) ? ( n38066 ) : ( VREG_16_1 ) ;
assign n38068 =  ( n2965 ) ? ( n38065 ) : ( n38067 ) ;
assign n38069 =  ( n1930 ) ? ( n38064 ) : ( n38068 ) ;
assign n38070 =  ( n879 ) ? ( n38059 ) : ( n38069 ) ;
assign n38071 =  ( n172 ) ? ( n5165 ) : ( VREG_16_1 ) ;
assign n38072 =  ( n170 ) ? ( n5164 ) : ( n38071 ) ;
assign n38073 =  ( n168 ) ? ( n5163 ) : ( n38072 ) ;
assign n38074 =  ( n166 ) ? ( n5162 ) : ( n38073 ) ;
assign n38075 =  ( n162 ) ? ( n5161 ) : ( n38074 ) ;
assign n38076 =  ( n172 ) ? ( n5175 ) : ( VREG_16_1 ) ;
assign n38077 =  ( n170 ) ? ( n5174 ) : ( n38076 ) ;
assign n38078 =  ( n168 ) ? ( n5173 ) : ( n38077 ) ;
assign n38079 =  ( n166 ) ? ( n5172 ) : ( n38078 ) ;
assign n38080 =  ( n162 ) ? ( n5171 ) : ( n38079 ) ;
assign n38081 =  ( n5154 ) ? ( VREG_16_1 ) : ( n38080 ) ;
assign n38082 =  ( n3051 ) ? ( n38081 ) : ( VREG_16_1 ) ;
assign n38083 =  ( n3040 ) ? ( n38075 ) : ( n38082 ) ;
assign n38084 =  ( n192 ) ? ( VREG_16_1 ) : ( VREG_16_1 ) ;
assign n38085 =  ( n157 ) ? ( n38083 ) : ( n38084 ) ;
assign n38086 =  ( n6 ) ? ( n38070 ) : ( n38085 ) ;
assign n38087 =  ( n351 ) ? ( n38086 ) : ( VREG_16_1 ) ;
assign n38088 =  ( n148 ) ? ( n6232 ) : ( VREG_16_10 ) ;
assign n38089 =  ( n146 ) ? ( n6231 ) : ( n38088 ) ;
assign n38090 =  ( n144 ) ? ( n6230 ) : ( n38089 ) ;
assign n38091 =  ( n142 ) ? ( n6229 ) : ( n38090 ) ;
assign n38092 =  ( n10 ) ? ( n6228 ) : ( n38091 ) ;
assign n38093 =  ( n148 ) ? ( n7266 ) : ( VREG_16_10 ) ;
assign n38094 =  ( n146 ) ? ( n7265 ) : ( n38093 ) ;
assign n38095 =  ( n144 ) ? ( n7264 ) : ( n38094 ) ;
assign n38096 =  ( n142 ) ? ( n7263 ) : ( n38095 ) ;
assign n38097 =  ( n10 ) ? ( n7262 ) : ( n38096 ) ;
assign n38098 =  ( n7273 ) ? ( VREG_16_10 ) : ( n38092 ) ;
assign n38099 =  ( n7273 ) ? ( VREG_16_10 ) : ( n38097 ) ;
assign n38100 =  ( n3034 ) ? ( n38099 ) : ( VREG_16_10 ) ;
assign n38101 =  ( n2965 ) ? ( n38098 ) : ( n38100 ) ;
assign n38102 =  ( n1930 ) ? ( n38097 ) : ( n38101 ) ;
assign n38103 =  ( n879 ) ? ( n38092 ) : ( n38102 ) ;
assign n38104 =  ( n172 ) ? ( n7284 ) : ( VREG_16_10 ) ;
assign n38105 =  ( n170 ) ? ( n7283 ) : ( n38104 ) ;
assign n38106 =  ( n168 ) ? ( n7282 ) : ( n38105 ) ;
assign n38107 =  ( n166 ) ? ( n7281 ) : ( n38106 ) ;
assign n38108 =  ( n162 ) ? ( n7280 ) : ( n38107 ) ;
assign n38109 =  ( n172 ) ? ( n7294 ) : ( VREG_16_10 ) ;
assign n38110 =  ( n170 ) ? ( n7293 ) : ( n38109 ) ;
assign n38111 =  ( n168 ) ? ( n7292 ) : ( n38110 ) ;
assign n38112 =  ( n166 ) ? ( n7291 ) : ( n38111 ) ;
assign n38113 =  ( n162 ) ? ( n7290 ) : ( n38112 ) ;
assign n38114 =  ( n7273 ) ? ( VREG_16_10 ) : ( n38113 ) ;
assign n38115 =  ( n3051 ) ? ( n38114 ) : ( VREG_16_10 ) ;
assign n38116 =  ( n3040 ) ? ( n38108 ) : ( n38115 ) ;
assign n38117 =  ( n192 ) ? ( VREG_16_10 ) : ( VREG_16_10 ) ;
assign n38118 =  ( n157 ) ? ( n38116 ) : ( n38117 ) ;
assign n38119 =  ( n6 ) ? ( n38103 ) : ( n38118 ) ;
assign n38120 =  ( n351 ) ? ( n38119 ) : ( VREG_16_10 ) ;
assign n38121 =  ( n148 ) ? ( n8351 ) : ( VREG_16_11 ) ;
assign n38122 =  ( n146 ) ? ( n8350 ) : ( n38121 ) ;
assign n38123 =  ( n144 ) ? ( n8349 ) : ( n38122 ) ;
assign n38124 =  ( n142 ) ? ( n8348 ) : ( n38123 ) ;
assign n38125 =  ( n10 ) ? ( n8347 ) : ( n38124 ) ;
assign n38126 =  ( n148 ) ? ( n9385 ) : ( VREG_16_11 ) ;
assign n38127 =  ( n146 ) ? ( n9384 ) : ( n38126 ) ;
assign n38128 =  ( n144 ) ? ( n9383 ) : ( n38127 ) ;
assign n38129 =  ( n142 ) ? ( n9382 ) : ( n38128 ) ;
assign n38130 =  ( n10 ) ? ( n9381 ) : ( n38129 ) ;
assign n38131 =  ( n9392 ) ? ( VREG_16_11 ) : ( n38125 ) ;
assign n38132 =  ( n9392 ) ? ( VREG_16_11 ) : ( n38130 ) ;
assign n38133 =  ( n3034 ) ? ( n38132 ) : ( VREG_16_11 ) ;
assign n38134 =  ( n2965 ) ? ( n38131 ) : ( n38133 ) ;
assign n38135 =  ( n1930 ) ? ( n38130 ) : ( n38134 ) ;
assign n38136 =  ( n879 ) ? ( n38125 ) : ( n38135 ) ;
assign n38137 =  ( n172 ) ? ( n9403 ) : ( VREG_16_11 ) ;
assign n38138 =  ( n170 ) ? ( n9402 ) : ( n38137 ) ;
assign n38139 =  ( n168 ) ? ( n9401 ) : ( n38138 ) ;
assign n38140 =  ( n166 ) ? ( n9400 ) : ( n38139 ) ;
assign n38141 =  ( n162 ) ? ( n9399 ) : ( n38140 ) ;
assign n38142 =  ( n172 ) ? ( n9413 ) : ( VREG_16_11 ) ;
assign n38143 =  ( n170 ) ? ( n9412 ) : ( n38142 ) ;
assign n38144 =  ( n168 ) ? ( n9411 ) : ( n38143 ) ;
assign n38145 =  ( n166 ) ? ( n9410 ) : ( n38144 ) ;
assign n38146 =  ( n162 ) ? ( n9409 ) : ( n38145 ) ;
assign n38147 =  ( n9392 ) ? ( VREG_16_11 ) : ( n38146 ) ;
assign n38148 =  ( n3051 ) ? ( n38147 ) : ( VREG_16_11 ) ;
assign n38149 =  ( n3040 ) ? ( n38141 ) : ( n38148 ) ;
assign n38150 =  ( n192 ) ? ( VREG_16_11 ) : ( VREG_16_11 ) ;
assign n38151 =  ( n157 ) ? ( n38149 ) : ( n38150 ) ;
assign n38152 =  ( n6 ) ? ( n38136 ) : ( n38151 ) ;
assign n38153 =  ( n351 ) ? ( n38152 ) : ( VREG_16_11 ) ;
assign n38154 =  ( n148 ) ? ( n10470 ) : ( VREG_16_12 ) ;
assign n38155 =  ( n146 ) ? ( n10469 ) : ( n38154 ) ;
assign n38156 =  ( n144 ) ? ( n10468 ) : ( n38155 ) ;
assign n38157 =  ( n142 ) ? ( n10467 ) : ( n38156 ) ;
assign n38158 =  ( n10 ) ? ( n10466 ) : ( n38157 ) ;
assign n38159 =  ( n148 ) ? ( n11504 ) : ( VREG_16_12 ) ;
assign n38160 =  ( n146 ) ? ( n11503 ) : ( n38159 ) ;
assign n38161 =  ( n144 ) ? ( n11502 ) : ( n38160 ) ;
assign n38162 =  ( n142 ) ? ( n11501 ) : ( n38161 ) ;
assign n38163 =  ( n10 ) ? ( n11500 ) : ( n38162 ) ;
assign n38164 =  ( n11511 ) ? ( VREG_16_12 ) : ( n38158 ) ;
assign n38165 =  ( n11511 ) ? ( VREG_16_12 ) : ( n38163 ) ;
assign n38166 =  ( n3034 ) ? ( n38165 ) : ( VREG_16_12 ) ;
assign n38167 =  ( n2965 ) ? ( n38164 ) : ( n38166 ) ;
assign n38168 =  ( n1930 ) ? ( n38163 ) : ( n38167 ) ;
assign n38169 =  ( n879 ) ? ( n38158 ) : ( n38168 ) ;
assign n38170 =  ( n172 ) ? ( n11522 ) : ( VREG_16_12 ) ;
assign n38171 =  ( n170 ) ? ( n11521 ) : ( n38170 ) ;
assign n38172 =  ( n168 ) ? ( n11520 ) : ( n38171 ) ;
assign n38173 =  ( n166 ) ? ( n11519 ) : ( n38172 ) ;
assign n38174 =  ( n162 ) ? ( n11518 ) : ( n38173 ) ;
assign n38175 =  ( n172 ) ? ( n11532 ) : ( VREG_16_12 ) ;
assign n38176 =  ( n170 ) ? ( n11531 ) : ( n38175 ) ;
assign n38177 =  ( n168 ) ? ( n11530 ) : ( n38176 ) ;
assign n38178 =  ( n166 ) ? ( n11529 ) : ( n38177 ) ;
assign n38179 =  ( n162 ) ? ( n11528 ) : ( n38178 ) ;
assign n38180 =  ( n11511 ) ? ( VREG_16_12 ) : ( n38179 ) ;
assign n38181 =  ( n3051 ) ? ( n38180 ) : ( VREG_16_12 ) ;
assign n38182 =  ( n3040 ) ? ( n38174 ) : ( n38181 ) ;
assign n38183 =  ( n192 ) ? ( VREG_16_12 ) : ( VREG_16_12 ) ;
assign n38184 =  ( n157 ) ? ( n38182 ) : ( n38183 ) ;
assign n38185 =  ( n6 ) ? ( n38169 ) : ( n38184 ) ;
assign n38186 =  ( n351 ) ? ( n38185 ) : ( VREG_16_12 ) ;
assign n38187 =  ( n148 ) ? ( n12589 ) : ( VREG_16_13 ) ;
assign n38188 =  ( n146 ) ? ( n12588 ) : ( n38187 ) ;
assign n38189 =  ( n144 ) ? ( n12587 ) : ( n38188 ) ;
assign n38190 =  ( n142 ) ? ( n12586 ) : ( n38189 ) ;
assign n38191 =  ( n10 ) ? ( n12585 ) : ( n38190 ) ;
assign n38192 =  ( n148 ) ? ( n13623 ) : ( VREG_16_13 ) ;
assign n38193 =  ( n146 ) ? ( n13622 ) : ( n38192 ) ;
assign n38194 =  ( n144 ) ? ( n13621 ) : ( n38193 ) ;
assign n38195 =  ( n142 ) ? ( n13620 ) : ( n38194 ) ;
assign n38196 =  ( n10 ) ? ( n13619 ) : ( n38195 ) ;
assign n38197 =  ( n13630 ) ? ( VREG_16_13 ) : ( n38191 ) ;
assign n38198 =  ( n13630 ) ? ( VREG_16_13 ) : ( n38196 ) ;
assign n38199 =  ( n3034 ) ? ( n38198 ) : ( VREG_16_13 ) ;
assign n38200 =  ( n2965 ) ? ( n38197 ) : ( n38199 ) ;
assign n38201 =  ( n1930 ) ? ( n38196 ) : ( n38200 ) ;
assign n38202 =  ( n879 ) ? ( n38191 ) : ( n38201 ) ;
assign n38203 =  ( n172 ) ? ( n13641 ) : ( VREG_16_13 ) ;
assign n38204 =  ( n170 ) ? ( n13640 ) : ( n38203 ) ;
assign n38205 =  ( n168 ) ? ( n13639 ) : ( n38204 ) ;
assign n38206 =  ( n166 ) ? ( n13638 ) : ( n38205 ) ;
assign n38207 =  ( n162 ) ? ( n13637 ) : ( n38206 ) ;
assign n38208 =  ( n172 ) ? ( n13651 ) : ( VREG_16_13 ) ;
assign n38209 =  ( n170 ) ? ( n13650 ) : ( n38208 ) ;
assign n38210 =  ( n168 ) ? ( n13649 ) : ( n38209 ) ;
assign n38211 =  ( n166 ) ? ( n13648 ) : ( n38210 ) ;
assign n38212 =  ( n162 ) ? ( n13647 ) : ( n38211 ) ;
assign n38213 =  ( n13630 ) ? ( VREG_16_13 ) : ( n38212 ) ;
assign n38214 =  ( n3051 ) ? ( n38213 ) : ( VREG_16_13 ) ;
assign n38215 =  ( n3040 ) ? ( n38207 ) : ( n38214 ) ;
assign n38216 =  ( n192 ) ? ( VREG_16_13 ) : ( VREG_16_13 ) ;
assign n38217 =  ( n157 ) ? ( n38215 ) : ( n38216 ) ;
assign n38218 =  ( n6 ) ? ( n38202 ) : ( n38217 ) ;
assign n38219 =  ( n351 ) ? ( n38218 ) : ( VREG_16_13 ) ;
assign n38220 =  ( n148 ) ? ( n14708 ) : ( VREG_16_14 ) ;
assign n38221 =  ( n146 ) ? ( n14707 ) : ( n38220 ) ;
assign n38222 =  ( n144 ) ? ( n14706 ) : ( n38221 ) ;
assign n38223 =  ( n142 ) ? ( n14705 ) : ( n38222 ) ;
assign n38224 =  ( n10 ) ? ( n14704 ) : ( n38223 ) ;
assign n38225 =  ( n148 ) ? ( n15742 ) : ( VREG_16_14 ) ;
assign n38226 =  ( n146 ) ? ( n15741 ) : ( n38225 ) ;
assign n38227 =  ( n144 ) ? ( n15740 ) : ( n38226 ) ;
assign n38228 =  ( n142 ) ? ( n15739 ) : ( n38227 ) ;
assign n38229 =  ( n10 ) ? ( n15738 ) : ( n38228 ) ;
assign n38230 =  ( n15749 ) ? ( VREG_16_14 ) : ( n38224 ) ;
assign n38231 =  ( n15749 ) ? ( VREG_16_14 ) : ( n38229 ) ;
assign n38232 =  ( n3034 ) ? ( n38231 ) : ( VREG_16_14 ) ;
assign n38233 =  ( n2965 ) ? ( n38230 ) : ( n38232 ) ;
assign n38234 =  ( n1930 ) ? ( n38229 ) : ( n38233 ) ;
assign n38235 =  ( n879 ) ? ( n38224 ) : ( n38234 ) ;
assign n38236 =  ( n172 ) ? ( n15760 ) : ( VREG_16_14 ) ;
assign n38237 =  ( n170 ) ? ( n15759 ) : ( n38236 ) ;
assign n38238 =  ( n168 ) ? ( n15758 ) : ( n38237 ) ;
assign n38239 =  ( n166 ) ? ( n15757 ) : ( n38238 ) ;
assign n38240 =  ( n162 ) ? ( n15756 ) : ( n38239 ) ;
assign n38241 =  ( n172 ) ? ( n15770 ) : ( VREG_16_14 ) ;
assign n38242 =  ( n170 ) ? ( n15769 ) : ( n38241 ) ;
assign n38243 =  ( n168 ) ? ( n15768 ) : ( n38242 ) ;
assign n38244 =  ( n166 ) ? ( n15767 ) : ( n38243 ) ;
assign n38245 =  ( n162 ) ? ( n15766 ) : ( n38244 ) ;
assign n38246 =  ( n15749 ) ? ( VREG_16_14 ) : ( n38245 ) ;
assign n38247 =  ( n3051 ) ? ( n38246 ) : ( VREG_16_14 ) ;
assign n38248 =  ( n3040 ) ? ( n38240 ) : ( n38247 ) ;
assign n38249 =  ( n192 ) ? ( VREG_16_14 ) : ( VREG_16_14 ) ;
assign n38250 =  ( n157 ) ? ( n38248 ) : ( n38249 ) ;
assign n38251 =  ( n6 ) ? ( n38235 ) : ( n38250 ) ;
assign n38252 =  ( n351 ) ? ( n38251 ) : ( VREG_16_14 ) ;
assign n38253 =  ( n148 ) ? ( n16827 ) : ( VREG_16_15 ) ;
assign n38254 =  ( n146 ) ? ( n16826 ) : ( n38253 ) ;
assign n38255 =  ( n144 ) ? ( n16825 ) : ( n38254 ) ;
assign n38256 =  ( n142 ) ? ( n16824 ) : ( n38255 ) ;
assign n38257 =  ( n10 ) ? ( n16823 ) : ( n38256 ) ;
assign n38258 =  ( n148 ) ? ( n17861 ) : ( VREG_16_15 ) ;
assign n38259 =  ( n146 ) ? ( n17860 ) : ( n38258 ) ;
assign n38260 =  ( n144 ) ? ( n17859 ) : ( n38259 ) ;
assign n38261 =  ( n142 ) ? ( n17858 ) : ( n38260 ) ;
assign n38262 =  ( n10 ) ? ( n17857 ) : ( n38261 ) ;
assign n38263 =  ( n17868 ) ? ( VREG_16_15 ) : ( n38257 ) ;
assign n38264 =  ( n17868 ) ? ( VREG_16_15 ) : ( n38262 ) ;
assign n38265 =  ( n3034 ) ? ( n38264 ) : ( VREG_16_15 ) ;
assign n38266 =  ( n2965 ) ? ( n38263 ) : ( n38265 ) ;
assign n38267 =  ( n1930 ) ? ( n38262 ) : ( n38266 ) ;
assign n38268 =  ( n879 ) ? ( n38257 ) : ( n38267 ) ;
assign n38269 =  ( n172 ) ? ( n17879 ) : ( VREG_16_15 ) ;
assign n38270 =  ( n170 ) ? ( n17878 ) : ( n38269 ) ;
assign n38271 =  ( n168 ) ? ( n17877 ) : ( n38270 ) ;
assign n38272 =  ( n166 ) ? ( n17876 ) : ( n38271 ) ;
assign n38273 =  ( n162 ) ? ( n17875 ) : ( n38272 ) ;
assign n38274 =  ( n172 ) ? ( n17889 ) : ( VREG_16_15 ) ;
assign n38275 =  ( n170 ) ? ( n17888 ) : ( n38274 ) ;
assign n38276 =  ( n168 ) ? ( n17887 ) : ( n38275 ) ;
assign n38277 =  ( n166 ) ? ( n17886 ) : ( n38276 ) ;
assign n38278 =  ( n162 ) ? ( n17885 ) : ( n38277 ) ;
assign n38279 =  ( n17868 ) ? ( VREG_16_15 ) : ( n38278 ) ;
assign n38280 =  ( n3051 ) ? ( n38279 ) : ( VREG_16_15 ) ;
assign n38281 =  ( n3040 ) ? ( n38273 ) : ( n38280 ) ;
assign n38282 =  ( n192 ) ? ( VREG_16_15 ) : ( VREG_16_15 ) ;
assign n38283 =  ( n157 ) ? ( n38281 ) : ( n38282 ) ;
assign n38284 =  ( n6 ) ? ( n38268 ) : ( n38283 ) ;
assign n38285 =  ( n351 ) ? ( n38284 ) : ( VREG_16_15 ) ;
assign n38286 =  ( n148 ) ? ( n18946 ) : ( VREG_16_2 ) ;
assign n38287 =  ( n146 ) ? ( n18945 ) : ( n38286 ) ;
assign n38288 =  ( n144 ) ? ( n18944 ) : ( n38287 ) ;
assign n38289 =  ( n142 ) ? ( n18943 ) : ( n38288 ) ;
assign n38290 =  ( n10 ) ? ( n18942 ) : ( n38289 ) ;
assign n38291 =  ( n148 ) ? ( n19980 ) : ( VREG_16_2 ) ;
assign n38292 =  ( n146 ) ? ( n19979 ) : ( n38291 ) ;
assign n38293 =  ( n144 ) ? ( n19978 ) : ( n38292 ) ;
assign n38294 =  ( n142 ) ? ( n19977 ) : ( n38293 ) ;
assign n38295 =  ( n10 ) ? ( n19976 ) : ( n38294 ) ;
assign n38296 =  ( n19987 ) ? ( VREG_16_2 ) : ( n38290 ) ;
assign n38297 =  ( n19987 ) ? ( VREG_16_2 ) : ( n38295 ) ;
assign n38298 =  ( n3034 ) ? ( n38297 ) : ( VREG_16_2 ) ;
assign n38299 =  ( n2965 ) ? ( n38296 ) : ( n38298 ) ;
assign n38300 =  ( n1930 ) ? ( n38295 ) : ( n38299 ) ;
assign n38301 =  ( n879 ) ? ( n38290 ) : ( n38300 ) ;
assign n38302 =  ( n172 ) ? ( n19998 ) : ( VREG_16_2 ) ;
assign n38303 =  ( n170 ) ? ( n19997 ) : ( n38302 ) ;
assign n38304 =  ( n168 ) ? ( n19996 ) : ( n38303 ) ;
assign n38305 =  ( n166 ) ? ( n19995 ) : ( n38304 ) ;
assign n38306 =  ( n162 ) ? ( n19994 ) : ( n38305 ) ;
assign n38307 =  ( n172 ) ? ( n20008 ) : ( VREG_16_2 ) ;
assign n38308 =  ( n170 ) ? ( n20007 ) : ( n38307 ) ;
assign n38309 =  ( n168 ) ? ( n20006 ) : ( n38308 ) ;
assign n38310 =  ( n166 ) ? ( n20005 ) : ( n38309 ) ;
assign n38311 =  ( n162 ) ? ( n20004 ) : ( n38310 ) ;
assign n38312 =  ( n19987 ) ? ( VREG_16_2 ) : ( n38311 ) ;
assign n38313 =  ( n3051 ) ? ( n38312 ) : ( VREG_16_2 ) ;
assign n38314 =  ( n3040 ) ? ( n38306 ) : ( n38313 ) ;
assign n38315 =  ( n192 ) ? ( VREG_16_2 ) : ( VREG_16_2 ) ;
assign n38316 =  ( n157 ) ? ( n38314 ) : ( n38315 ) ;
assign n38317 =  ( n6 ) ? ( n38301 ) : ( n38316 ) ;
assign n38318 =  ( n351 ) ? ( n38317 ) : ( VREG_16_2 ) ;
assign n38319 =  ( n148 ) ? ( n21065 ) : ( VREG_16_3 ) ;
assign n38320 =  ( n146 ) ? ( n21064 ) : ( n38319 ) ;
assign n38321 =  ( n144 ) ? ( n21063 ) : ( n38320 ) ;
assign n38322 =  ( n142 ) ? ( n21062 ) : ( n38321 ) ;
assign n38323 =  ( n10 ) ? ( n21061 ) : ( n38322 ) ;
assign n38324 =  ( n148 ) ? ( n22099 ) : ( VREG_16_3 ) ;
assign n38325 =  ( n146 ) ? ( n22098 ) : ( n38324 ) ;
assign n38326 =  ( n144 ) ? ( n22097 ) : ( n38325 ) ;
assign n38327 =  ( n142 ) ? ( n22096 ) : ( n38326 ) ;
assign n38328 =  ( n10 ) ? ( n22095 ) : ( n38327 ) ;
assign n38329 =  ( n22106 ) ? ( VREG_16_3 ) : ( n38323 ) ;
assign n38330 =  ( n22106 ) ? ( VREG_16_3 ) : ( n38328 ) ;
assign n38331 =  ( n3034 ) ? ( n38330 ) : ( VREG_16_3 ) ;
assign n38332 =  ( n2965 ) ? ( n38329 ) : ( n38331 ) ;
assign n38333 =  ( n1930 ) ? ( n38328 ) : ( n38332 ) ;
assign n38334 =  ( n879 ) ? ( n38323 ) : ( n38333 ) ;
assign n38335 =  ( n172 ) ? ( n22117 ) : ( VREG_16_3 ) ;
assign n38336 =  ( n170 ) ? ( n22116 ) : ( n38335 ) ;
assign n38337 =  ( n168 ) ? ( n22115 ) : ( n38336 ) ;
assign n38338 =  ( n166 ) ? ( n22114 ) : ( n38337 ) ;
assign n38339 =  ( n162 ) ? ( n22113 ) : ( n38338 ) ;
assign n38340 =  ( n172 ) ? ( n22127 ) : ( VREG_16_3 ) ;
assign n38341 =  ( n170 ) ? ( n22126 ) : ( n38340 ) ;
assign n38342 =  ( n168 ) ? ( n22125 ) : ( n38341 ) ;
assign n38343 =  ( n166 ) ? ( n22124 ) : ( n38342 ) ;
assign n38344 =  ( n162 ) ? ( n22123 ) : ( n38343 ) ;
assign n38345 =  ( n22106 ) ? ( VREG_16_3 ) : ( n38344 ) ;
assign n38346 =  ( n3051 ) ? ( n38345 ) : ( VREG_16_3 ) ;
assign n38347 =  ( n3040 ) ? ( n38339 ) : ( n38346 ) ;
assign n38348 =  ( n192 ) ? ( VREG_16_3 ) : ( VREG_16_3 ) ;
assign n38349 =  ( n157 ) ? ( n38347 ) : ( n38348 ) ;
assign n38350 =  ( n6 ) ? ( n38334 ) : ( n38349 ) ;
assign n38351 =  ( n351 ) ? ( n38350 ) : ( VREG_16_3 ) ;
assign n38352 =  ( n148 ) ? ( n23184 ) : ( VREG_16_4 ) ;
assign n38353 =  ( n146 ) ? ( n23183 ) : ( n38352 ) ;
assign n38354 =  ( n144 ) ? ( n23182 ) : ( n38353 ) ;
assign n38355 =  ( n142 ) ? ( n23181 ) : ( n38354 ) ;
assign n38356 =  ( n10 ) ? ( n23180 ) : ( n38355 ) ;
assign n38357 =  ( n148 ) ? ( n24218 ) : ( VREG_16_4 ) ;
assign n38358 =  ( n146 ) ? ( n24217 ) : ( n38357 ) ;
assign n38359 =  ( n144 ) ? ( n24216 ) : ( n38358 ) ;
assign n38360 =  ( n142 ) ? ( n24215 ) : ( n38359 ) ;
assign n38361 =  ( n10 ) ? ( n24214 ) : ( n38360 ) ;
assign n38362 =  ( n24225 ) ? ( VREG_16_4 ) : ( n38356 ) ;
assign n38363 =  ( n24225 ) ? ( VREG_16_4 ) : ( n38361 ) ;
assign n38364 =  ( n3034 ) ? ( n38363 ) : ( VREG_16_4 ) ;
assign n38365 =  ( n2965 ) ? ( n38362 ) : ( n38364 ) ;
assign n38366 =  ( n1930 ) ? ( n38361 ) : ( n38365 ) ;
assign n38367 =  ( n879 ) ? ( n38356 ) : ( n38366 ) ;
assign n38368 =  ( n172 ) ? ( n24236 ) : ( VREG_16_4 ) ;
assign n38369 =  ( n170 ) ? ( n24235 ) : ( n38368 ) ;
assign n38370 =  ( n168 ) ? ( n24234 ) : ( n38369 ) ;
assign n38371 =  ( n166 ) ? ( n24233 ) : ( n38370 ) ;
assign n38372 =  ( n162 ) ? ( n24232 ) : ( n38371 ) ;
assign n38373 =  ( n172 ) ? ( n24246 ) : ( VREG_16_4 ) ;
assign n38374 =  ( n170 ) ? ( n24245 ) : ( n38373 ) ;
assign n38375 =  ( n168 ) ? ( n24244 ) : ( n38374 ) ;
assign n38376 =  ( n166 ) ? ( n24243 ) : ( n38375 ) ;
assign n38377 =  ( n162 ) ? ( n24242 ) : ( n38376 ) ;
assign n38378 =  ( n24225 ) ? ( VREG_16_4 ) : ( n38377 ) ;
assign n38379 =  ( n3051 ) ? ( n38378 ) : ( VREG_16_4 ) ;
assign n38380 =  ( n3040 ) ? ( n38372 ) : ( n38379 ) ;
assign n38381 =  ( n192 ) ? ( VREG_16_4 ) : ( VREG_16_4 ) ;
assign n38382 =  ( n157 ) ? ( n38380 ) : ( n38381 ) ;
assign n38383 =  ( n6 ) ? ( n38367 ) : ( n38382 ) ;
assign n38384 =  ( n351 ) ? ( n38383 ) : ( VREG_16_4 ) ;
assign n38385 =  ( n148 ) ? ( n25303 ) : ( VREG_16_5 ) ;
assign n38386 =  ( n146 ) ? ( n25302 ) : ( n38385 ) ;
assign n38387 =  ( n144 ) ? ( n25301 ) : ( n38386 ) ;
assign n38388 =  ( n142 ) ? ( n25300 ) : ( n38387 ) ;
assign n38389 =  ( n10 ) ? ( n25299 ) : ( n38388 ) ;
assign n38390 =  ( n148 ) ? ( n26337 ) : ( VREG_16_5 ) ;
assign n38391 =  ( n146 ) ? ( n26336 ) : ( n38390 ) ;
assign n38392 =  ( n144 ) ? ( n26335 ) : ( n38391 ) ;
assign n38393 =  ( n142 ) ? ( n26334 ) : ( n38392 ) ;
assign n38394 =  ( n10 ) ? ( n26333 ) : ( n38393 ) ;
assign n38395 =  ( n26344 ) ? ( VREG_16_5 ) : ( n38389 ) ;
assign n38396 =  ( n26344 ) ? ( VREG_16_5 ) : ( n38394 ) ;
assign n38397 =  ( n3034 ) ? ( n38396 ) : ( VREG_16_5 ) ;
assign n38398 =  ( n2965 ) ? ( n38395 ) : ( n38397 ) ;
assign n38399 =  ( n1930 ) ? ( n38394 ) : ( n38398 ) ;
assign n38400 =  ( n879 ) ? ( n38389 ) : ( n38399 ) ;
assign n38401 =  ( n172 ) ? ( n26355 ) : ( VREG_16_5 ) ;
assign n38402 =  ( n170 ) ? ( n26354 ) : ( n38401 ) ;
assign n38403 =  ( n168 ) ? ( n26353 ) : ( n38402 ) ;
assign n38404 =  ( n166 ) ? ( n26352 ) : ( n38403 ) ;
assign n38405 =  ( n162 ) ? ( n26351 ) : ( n38404 ) ;
assign n38406 =  ( n172 ) ? ( n26365 ) : ( VREG_16_5 ) ;
assign n38407 =  ( n170 ) ? ( n26364 ) : ( n38406 ) ;
assign n38408 =  ( n168 ) ? ( n26363 ) : ( n38407 ) ;
assign n38409 =  ( n166 ) ? ( n26362 ) : ( n38408 ) ;
assign n38410 =  ( n162 ) ? ( n26361 ) : ( n38409 ) ;
assign n38411 =  ( n26344 ) ? ( VREG_16_5 ) : ( n38410 ) ;
assign n38412 =  ( n3051 ) ? ( n38411 ) : ( VREG_16_5 ) ;
assign n38413 =  ( n3040 ) ? ( n38405 ) : ( n38412 ) ;
assign n38414 =  ( n192 ) ? ( VREG_16_5 ) : ( VREG_16_5 ) ;
assign n38415 =  ( n157 ) ? ( n38413 ) : ( n38414 ) ;
assign n38416 =  ( n6 ) ? ( n38400 ) : ( n38415 ) ;
assign n38417 =  ( n351 ) ? ( n38416 ) : ( VREG_16_5 ) ;
assign n38418 =  ( n148 ) ? ( n27422 ) : ( VREG_16_6 ) ;
assign n38419 =  ( n146 ) ? ( n27421 ) : ( n38418 ) ;
assign n38420 =  ( n144 ) ? ( n27420 ) : ( n38419 ) ;
assign n38421 =  ( n142 ) ? ( n27419 ) : ( n38420 ) ;
assign n38422 =  ( n10 ) ? ( n27418 ) : ( n38421 ) ;
assign n38423 =  ( n148 ) ? ( n28456 ) : ( VREG_16_6 ) ;
assign n38424 =  ( n146 ) ? ( n28455 ) : ( n38423 ) ;
assign n38425 =  ( n144 ) ? ( n28454 ) : ( n38424 ) ;
assign n38426 =  ( n142 ) ? ( n28453 ) : ( n38425 ) ;
assign n38427 =  ( n10 ) ? ( n28452 ) : ( n38426 ) ;
assign n38428 =  ( n28463 ) ? ( VREG_16_6 ) : ( n38422 ) ;
assign n38429 =  ( n28463 ) ? ( VREG_16_6 ) : ( n38427 ) ;
assign n38430 =  ( n3034 ) ? ( n38429 ) : ( VREG_16_6 ) ;
assign n38431 =  ( n2965 ) ? ( n38428 ) : ( n38430 ) ;
assign n38432 =  ( n1930 ) ? ( n38427 ) : ( n38431 ) ;
assign n38433 =  ( n879 ) ? ( n38422 ) : ( n38432 ) ;
assign n38434 =  ( n172 ) ? ( n28474 ) : ( VREG_16_6 ) ;
assign n38435 =  ( n170 ) ? ( n28473 ) : ( n38434 ) ;
assign n38436 =  ( n168 ) ? ( n28472 ) : ( n38435 ) ;
assign n38437 =  ( n166 ) ? ( n28471 ) : ( n38436 ) ;
assign n38438 =  ( n162 ) ? ( n28470 ) : ( n38437 ) ;
assign n38439 =  ( n172 ) ? ( n28484 ) : ( VREG_16_6 ) ;
assign n38440 =  ( n170 ) ? ( n28483 ) : ( n38439 ) ;
assign n38441 =  ( n168 ) ? ( n28482 ) : ( n38440 ) ;
assign n38442 =  ( n166 ) ? ( n28481 ) : ( n38441 ) ;
assign n38443 =  ( n162 ) ? ( n28480 ) : ( n38442 ) ;
assign n38444 =  ( n28463 ) ? ( VREG_16_6 ) : ( n38443 ) ;
assign n38445 =  ( n3051 ) ? ( n38444 ) : ( VREG_16_6 ) ;
assign n38446 =  ( n3040 ) ? ( n38438 ) : ( n38445 ) ;
assign n38447 =  ( n192 ) ? ( VREG_16_6 ) : ( VREG_16_6 ) ;
assign n38448 =  ( n157 ) ? ( n38446 ) : ( n38447 ) ;
assign n38449 =  ( n6 ) ? ( n38433 ) : ( n38448 ) ;
assign n38450 =  ( n351 ) ? ( n38449 ) : ( VREG_16_6 ) ;
assign n38451 =  ( n148 ) ? ( n29541 ) : ( VREG_16_7 ) ;
assign n38452 =  ( n146 ) ? ( n29540 ) : ( n38451 ) ;
assign n38453 =  ( n144 ) ? ( n29539 ) : ( n38452 ) ;
assign n38454 =  ( n142 ) ? ( n29538 ) : ( n38453 ) ;
assign n38455 =  ( n10 ) ? ( n29537 ) : ( n38454 ) ;
assign n38456 =  ( n148 ) ? ( n30575 ) : ( VREG_16_7 ) ;
assign n38457 =  ( n146 ) ? ( n30574 ) : ( n38456 ) ;
assign n38458 =  ( n144 ) ? ( n30573 ) : ( n38457 ) ;
assign n38459 =  ( n142 ) ? ( n30572 ) : ( n38458 ) ;
assign n38460 =  ( n10 ) ? ( n30571 ) : ( n38459 ) ;
assign n38461 =  ( n30582 ) ? ( VREG_16_7 ) : ( n38455 ) ;
assign n38462 =  ( n30582 ) ? ( VREG_16_7 ) : ( n38460 ) ;
assign n38463 =  ( n3034 ) ? ( n38462 ) : ( VREG_16_7 ) ;
assign n38464 =  ( n2965 ) ? ( n38461 ) : ( n38463 ) ;
assign n38465 =  ( n1930 ) ? ( n38460 ) : ( n38464 ) ;
assign n38466 =  ( n879 ) ? ( n38455 ) : ( n38465 ) ;
assign n38467 =  ( n172 ) ? ( n30593 ) : ( VREG_16_7 ) ;
assign n38468 =  ( n170 ) ? ( n30592 ) : ( n38467 ) ;
assign n38469 =  ( n168 ) ? ( n30591 ) : ( n38468 ) ;
assign n38470 =  ( n166 ) ? ( n30590 ) : ( n38469 ) ;
assign n38471 =  ( n162 ) ? ( n30589 ) : ( n38470 ) ;
assign n38472 =  ( n172 ) ? ( n30603 ) : ( VREG_16_7 ) ;
assign n38473 =  ( n170 ) ? ( n30602 ) : ( n38472 ) ;
assign n38474 =  ( n168 ) ? ( n30601 ) : ( n38473 ) ;
assign n38475 =  ( n166 ) ? ( n30600 ) : ( n38474 ) ;
assign n38476 =  ( n162 ) ? ( n30599 ) : ( n38475 ) ;
assign n38477 =  ( n30582 ) ? ( VREG_16_7 ) : ( n38476 ) ;
assign n38478 =  ( n3051 ) ? ( n38477 ) : ( VREG_16_7 ) ;
assign n38479 =  ( n3040 ) ? ( n38471 ) : ( n38478 ) ;
assign n38480 =  ( n192 ) ? ( VREG_16_7 ) : ( VREG_16_7 ) ;
assign n38481 =  ( n157 ) ? ( n38479 ) : ( n38480 ) ;
assign n38482 =  ( n6 ) ? ( n38466 ) : ( n38481 ) ;
assign n38483 =  ( n351 ) ? ( n38482 ) : ( VREG_16_7 ) ;
assign n38484 =  ( n148 ) ? ( n31660 ) : ( VREG_16_8 ) ;
assign n38485 =  ( n146 ) ? ( n31659 ) : ( n38484 ) ;
assign n38486 =  ( n144 ) ? ( n31658 ) : ( n38485 ) ;
assign n38487 =  ( n142 ) ? ( n31657 ) : ( n38486 ) ;
assign n38488 =  ( n10 ) ? ( n31656 ) : ( n38487 ) ;
assign n38489 =  ( n148 ) ? ( n32694 ) : ( VREG_16_8 ) ;
assign n38490 =  ( n146 ) ? ( n32693 ) : ( n38489 ) ;
assign n38491 =  ( n144 ) ? ( n32692 ) : ( n38490 ) ;
assign n38492 =  ( n142 ) ? ( n32691 ) : ( n38491 ) ;
assign n38493 =  ( n10 ) ? ( n32690 ) : ( n38492 ) ;
assign n38494 =  ( n32701 ) ? ( VREG_16_8 ) : ( n38488 ) ;
assign n38495 =  ( n32701 ) ? ( VREG_16_8 ) : ( n38493 ) ;
assign n38496 =  ( n3034 ) ? ( n38495 ) : ( VREG_16_8 ) ;
assign n38497 =  ( n2965 ) ? ( n38494 ) : ( n38496 ) ;
assign n38498 =  ( n1930 ) ? ( n38493 ) : ( n38497 ) ;
assign n38499 =  ( n879 ) ? ( n38488 ) : ( n38498 ) ;
assign n38500 =  ( n172 ) ? ( n32712 ) : ( VREG_16_8 ) ;
assign n38501 =  ( n170 ) ? ( n32711 ) : ( n38500 ) ;
assign n38502 =  ( n168 ) ? ( n32710 ) : ( n38501 ) ;
assign n38503 =  ( n166 ) ? ( n32709 ) : ( n38502 ) ;
assign n38504 =  ( n162 ) ? ( n32708 ) : ( n38503 ) ;
assign n38505 =  ( n172 ) ? ( n32722 ) : ( VREG_16_8 ) ;
assign n38506 =  ( n170 ) ? ( n32721 ) : ( n38505 ) ;
assign n38507 =  ( n168 ) ? ( n32720 ) : ( n38506 ) ;
assign n38508 =  ( n166 ) ? ( n32719 ) : ( n38507 ) ;
assign n38509 =  ( n162 ) ? ( n32718 ) : ( n38508 ) ;
assign n38510 =  ( n32701 ) ? ( VREG_16_8 ) : ( n38509 ) ;
assign n38511 =  ( n3051 ) ? ( n38510 ) : ( VREG_16_8 ) ;
assign n38512 =  ( n3040 ) ? ( n38504 ) : ( n38511 ) ;
assign n38513 =  ( n192 ) ? ( VREG_16_8 ) : ( VREG_16_8 ) ;
assign n38514 =  ( n157 ) ? ( n38512 ) : ( n38513 ) ;
assign n38515 =  ( n6 ) ? ( n38499 ) : ( n38514 ) ;
assign n38516 =  ( n351 ) ? ( n38515 ) : ( VREG_16_8 ) ;
assign n38517 =  ( n148 ) ? ( n33779 ) : ( VREG_16_9 ) ;
assign n38518 =  ( n146 ) ? ( n33778 ) : ( n38517 ) ;
assign n38519 =  ( n144 ) ? ( n33777 ) : ( n38518 ) ;
assign n38520 =  ( n142 ) ? ( n33776 ) : ( n38519 ) ;
assign n38521 =  ( n10 ) ? ( n33775 ) : ( n38520 ) ;
assign n38522 =  ( n148 ) ? ( n34813 ) : ( VREG_16_9 ) ;
assign n38523 =  ( n146 ) ? ( n34812 ) : ( n38522 ) ;
assign n38524 =  ( n144 ) ? ( n34811 ) : ( n38523 ) ;
assign n38525 =  ( n142 ) ? ( n34810 ) : ( n38524 ) ;
assign n38526 =  ( n10 ) ? ( n34809 ) : ( n38525 ) ;
assign n38527 =  ( n34820 ) ? ( VREG_16_9 ) : ( n38521 ) ;
assign n38528 =  ( n34820 ) ? ( VREG_16_9 ) : ( n38526 ) ;
assign n38529 =  ( n3034 ) ? ( n38528 ) : ( VREG_16_9 ) ;
assign n38530 =  ( n2965 ) ? ( n38527 ) : ( n38529 ) ;
assign n38531 =  ( n1930 ) ? ( n38526 ) : ( n38530 ) ;
assign n38532 =  ( n879 ) ? ( n38521 ) : ( n38531 ) ;
assign n38533 =  ( n172 ) ? ( n34831 ) : ( VREG_16_9 ) ;
assign n38534 =  ( n170 ) ? ( n34830 ) : ( n38533 ) ;
assign n38535 =  ( n168 ) ? ( n34829 ) : ( n38534 ) ;
assign n38536 =  ( n166 ) ? ( n34828 ) : ( n38535 ) ;
assign n38537 =  ( n162 ) ? ( n34827 ) : ( n38536 ) ;
assign n38538 =  ( n172 ) ? ( n34841 ) : ( VREG_16_9 ) ;
assign n38539 =  ( n170 ) ? ( n34840 ) : ( n38538 ) ;
assign n38540 =  ( n168 ) ? ( n34839 ) : ( n38539 ) ;
assign n38541 =  ( n166 ) ? ( n34838 ) : ( n38540 ) ;
assign n38542 =  ( n162 ) ? ( n34837 ) : ( n38541 ) ;
assign n38543 =  ( n34820 ) ? ( VREG_16_9 ) : ( n38542 ) ;
assign n38544 =  ( n3051 ) ? ( n38543 ) : ( VREG_16_9 ) ;
assign n38545 =  ( n3040 ) ? ( n38537 ) : ( n38544 ) ;
assign n38546 =  ( n192 ) ? ( VREG_16_9 ) : ( VREG_16_9 ) ;
assign n38547 =  ( n157 ) ? ( n38545 ) : ( n38546 ) ;
assign n38548 =  ( n6 ) ? ( n38532 ) : ( n38547 ) ;
assign n38549 =  ( n351 ) ? ( n38548 ) : ( VREG_16_9 ) ;
assign n38550 =  ( n148 ) ? ( n1924 ) : ( VREG_17_0 ) ;
assign n38551 =  ( n146 ) ? ( n1923 ) : ( n38550 ) ;
assign n38552 =  ( n144 ) ? ( n1922 ) : ( n38551 ) ;
assign n38553 =  ( n142 ) ? ( n1921 ) : ( n38552 ) ;
assign n38554 =  ( n10 ) ? ( n1920 ) : ( n38553 ) ;
assign n38555 =  ( n148 ) ? ( n2959 ) : ( VREG_17_0 ) ;
assign n38556 =  ( n146 ) ? ( n2958 ) : ( n38555 ) ;
assign n38557 =  ( n144 ) ? ( n2957 ) : ( n38556 ) ;
assign n38558 =  ( n142 ) ? ( n2956 ) : ( n38557 ) ;
assign n38559 =  ( n10 ) ? ( n2955 ) : ( n38558 ) ;
assign n38560 =  ( n3032 ) ? ( VREG_17_0 ) : ( n38554 ) ;
assign n38561 =  ( n3032 ) ? ( VREG_17_0 ) : ( n38559 ) ;
assign n38562 =  ( n3034 ) ? ( n38561 ) : ( VREG_17_0 ) ;
assign n38563 =  ( n2965 ) ? ( n38560 ) : ( n38562 ) ;
assign n38564 =  ( n1930 ) ? ( n38559 ) : ( n38563 ) ;
assign n38565 =  ( n879 ) ? ( n38554 ) : ( n38564 ) ;
assign n38566 =  ( n172 ) ? ( n3045 ) : ( VREG_17_0 ) ;
assign n38567 =  ( n170 ) ? ( n3044 ) : ( n38566 ) ;
assign n38568 =  ( n168 ) ? ( n3043 ) : ( n38567 ) ;
assign n38569 =  ( n166 ) ? ( n3042 ) : ( n38568 ) ;
assign n38570 =  ( n162 ) ? ( n3041 ) : ( n38569 ) ;
assign n38571 =  ( n172 ) ? ( n3056 ) : ( VREG_17_0 ) ;
assign n38572 =  ( n170 ) ? ( n3055 ) : ( n38571 ) ;
assign n38573 =  ( n168 ) ? ( n3054 ) : ( n38572 ) ;
assign n38574 =  ( n166 ) ? ( n3053 ) : ( n38573 ) ;
assign n38575 =  ( n162 ) ? ( n3052 ) : ( n38574 ) ;
assign n38576 =  ( n3032 ) ? ( VREG_17_0 ) : ( n38575 ) ;
assign n38577 =  ( n3051 ) ? ( n38576 ) : ( VREG_17_0 ) ;
assign n38578 =  ( n3040 ) ? ( n38570 ) : ( n38577 ) ;
assign n38579 =  ( n192 ) ? ( VREG_17_0 ) : ( VREG_17_0 ) ;
assign n38580 =  ( n157 ) ? ( n38578 ) : ( n38579 ) ;
assign n38581 =  ( n6 ) ? ( n38565 ) : ( n38580 ) ;
assign n38582 =  ( n373 ) ? ( n38581 ) : ( VREG_17_0 ) ;
assign n38583 =  ( n148 ) ? ( n4113 ) : ( VREG_17_1 ) ;
assign n38584 =  ( n146 ) ? ( n4112 ) : ( n38583 ) ;
assign n38585 =  ( n144 ) ? ( n4111 ) : ( n38584 ) ;
assign n38586 =  ( n142 ) ? ( n4110 ) : ( n38585 ) ;
assign n38587 =  ( n10 ) ? ( n4109 ) : ( n38586 ) ;
assign n38588 =  ( n148 ) ? ( n5147 ) : ( VREG_17_1 ) ;
assign n38589 =  ( n146 ) ? ( n5146 ) : ( n38588 ) ;
assign n38590 =  ( n144 ) ? ( n5145 ) : ( n38589 ) ;
assign n38591 =  ( n142 ) ? ( n5144 ) : ( n38590 ) ;
assign n38592 =  ( n10 ) ? ( n5143 ) : ( n38591 ) ;
assign n38593 =  ( n5154 ) ? ( VREG_17_1 ) : ( n38587 ) ;
assign n38594 =  ( n5154 ) ? ( VREG_17_1 ) : ( n38592 ) ;
assign n38595 =  ( n3034 ) ? ( n38594 ) : ( VREG_17_1 ) ;
assign n38596 =  ( n2965 ) ? ( n38593 ) : ( n38595 ) ;
assign n38597 =  ( n1930 ) ? ( n38592 ) : ( n38596 ) ;
assign n38598 =  ( n879 ) ? ( n38587 ) : ( n38597 ) ;
assign n38599 =  ( n172 ) ? ( n5165 ) : ( VREG_17_1 ) ;
assign n38600 =  ( n170 ) ? ( n5164 ) : ( n38599 ) ;
assign n38601 =  ( n168 ) ? ( n5163 ) : ( n38600 ) ;
assign n38602 =  ( n166 ) ? ( n5162 ) : ( n38601 ) ;
assign n38603 =  ( n162 ) ? ( n5161 ) : ( n38602 ) ;
assign n38604 =  ( n172 ) ? ( n5175 ) : ( VREG_17_1 ) ;
assign n38605 =  ( n170 ) ? ( n5174 ) : ( n38604 ) ;
assign n38606 =  ( n168 ) ? ( n5173 ) : ( n38605 ) ;
assign n38607 =  ( n166 ) ? ( n5172 ) : ( n38606 ) ;
assign n38608 =  ( n162 ) ? ( n5171 ) : ( n38607 ) ;
assign n38609 =  ( n5154 ) ? ( VREG_17_1 ) : ( n38608 ) ;
assign n38610 =  ( n3051 ) ? ( n38609 ) : ( VREG_17_1 ) ;
assign n38611 =  ( n3040 ) ? ( n38603 ) : ( n38610 ) ;
assign n38612 =  ( n192 ) ? ( VREG_17_1 ) : ( VREG_17_1 ) ;
assign n38613 =  ( n157 ) ? ( n38611 ) : ( n38612 ) ;
assign n38614 =  ( n6 ) ? ( n38598 ) : ( n38613 ) ;
assign n38615 =  ( n373 ) ? ( n38614 ) : ( VREG_17_1 ) ;
assign n38616 =  ( n148 ) ? ( n6232 ) : ( VREG_17_10 ) ;
assign n38617 =  ( n146 ) ? ( n6231 ) : ( n38616 ) ;
assign n38618 =  ( n144 ) ? ( n6230 ) : ( n38617 ) ;
assign n38619 =  ( n142 ) ? ( n6229 ) : ( n38618 ) ;
assign n38620 =  ( n10 ) ? ( n6228 ) : ( n38619 ) ;
assign n38621 =  ( n148 ) ? ( n7266 ) : ( VREG_17_10 ) ;
assign n38622 =  ( n146 ) ? ( n7265 ) : ( n38621 ) ;
assign n38623 =  ( n144 ) ? ( n7264 ) : ( n38622 ) ;
assign n38624 =  ( n142 ) ? ( n7263 ) : ( n38623 ) ;
assign n38625 =  ( n10 ) ? ( n7262 ) : ( n38624 ) ;
assign n38626 =  ( n7273 ) ? ( VREG_17_10 ) : ( n38620 ) ;
assign n38627 =  ( n7273 ) ? ( VREG_17_10 ) : ( n38625 ) ;
assign n38628 =  ( n3034 ) ? ( n38627 ) : ( VREG_17_10 ) ;
assign n38629 =  ( n2965 ) ? ( n38626 ) : ( n38628 ) ;
assign n38630 =  ( n1930 ) ? ( n38625 ) : ( n38629 ) ;
assign n38631 =  ( n879 ) ? ( n38620 ) : ( n38630 ) ;
assign n38632 =  ( n172 ) ? ( n7284 ) : ( VREG_17_10 ) ;
assign n38633 =  ( n170 ) ? ( n7283 ) : ( n38632 ) ;
assign n38634 =  ( n168 ) ? ( n7282 ) : ( n38633 ) ;
assign n38635 =  ( n166 ) ? ( n7281 ) : ( n38634 ) ;
assign n38636 =  ( n162 ) ? ( n7280 ) : ( n38635 ) ;
assign n38637 =  ( n172 ) ? ( n7294 ) : ( VREG_17_10 ) ;
assign n38638 =  ( n170 ) ? ( n7293 ) : ( n38637 ) ;
assign n38639 =  ( n168 ) ? ( n7292 ) : ( n38638 ) ;
assign n38640 =  ( n166 ) ? ( n7291 ) : ( n38639 ) ;
assign n38641 =  ( n162 ) ? ( n7290 ) : ( n38640 ) ;
assign n38642 =  ( n7273 ) ? ( VREG_17_10 ) : ( n38641 ) ;
assign n38643 =  ( n3051 ) ? ( n38642 ) : ( VREG_17_10 ) ;
assign n38644 =  ( n3040 ) ? ( n38636 ) : ( n38643 ) ;
assign n38645 =  ( n192 ) ? ( VREG_17_10 ) : ( VREG_17_10 ) ;
assign n38646 =  ( n157 ) ? ( n38644 ) : ( n38645 ) ;
assign n38647 =  ( n6 ) ? ( n38631 ) : ( n38646 ) ;
assign n38648 =  ( n373 ) ? ( n38647 ) : ( VREG_17_10 ) ;
assign n38649 =  ( n148 ) ? ( n8351 ) : ( VREG_17_11 ) ;
assign n38650 =  ( n146 ) ? ( n8350 ) : ( n38649 ) ;
assign n38651 =  ( n144 ) ? ( n8349 ) : ( n38650 ) ;
assign n38652 =  ( n142 ) ? ( n8348 ) : ( n38651 ) ;
assign n38653 =  ( n10 ) ? ( n8347 ) : ( n38652 ) ;
assign n38654 =  ( n148 ) ? ( n9385 ) : ( VREG_17_11 ) ;
assign n38655 =  ( n146 ) ? ( n9384 ) : ( n38654 ) ;
assign n38656 =  ( n144 ) ? ( n9383 ) : ( n38655 ) ;
assign n38657 =  ( n142 ) ? ( n9382 ) : ( n38656 ) ;
assign n38658 =  ( n10 ) ? ( n9381 ) : ( n38657 ) ;
assign n38659 =  ( n9392 ) ? ( VREG_17_11 ) : ( n38653 ) ;
assign n38660 =  ( n9392 ) ? ( VREG_17_11 ) : ( n38658 ) ;
assign n38661 =  ( n3034 ) ? ( n38660 ) : ( VREG_17_11 ) ;
assign n38662 =  ( n2965 ) ? ( n38659 ) : ( n38661 ) ;
assign n38663 =  ( n1930 ) ? ( n38658 ) : ( n38662 ) ;
assign n38664 =  ( n879 ) ? ( n38653 ) : ( n38663 ) ;
assign n38665 =  ( n172 ) ? ( n9403 ) : ( VREG_17_11 ) ;
assign n38666 =  ( n170 ) ? ( n9402 ) : ( n38665 ) ;
assign n38667 =  ( n168 ) ? ( n9401 ) : ( n38666 ) ;
assign n38668 =  ( n166 ) ? ( n9400 ) : ( n38667 ) ;
assign n38669 =  ( n162 ) ? ( n9399 ) : ( n38668 ) ;
assign n38670 =  ( n172 ) ? ( n9413 ) : ( VREG_17_11 ) ;
assign n38671 =  ( n170 ) ? ( n9412 ) : ( n38670 ) ;
assign n38672 =  ( n168 ) ? ( n9411 ) : ( n38671 ) ;
assign n38673 =  ( n166 ) ? ( n9410 ) : ( n38672 ) ;
assign n38674 =  ( n162 ) ? ( n9409 ) : ( n38673 ) ;
assign n38675 =  ( n9392 ) ? ( VREG_17_11 ) : ( n38674 ) ;
assign n38676 =  ( n3051 ) ? ( n38675 ) : ( VREG_17_11 ) ;
assign n38677 =  ( n3040 ) ? ( n38669 ) : ( n38676 ) ;
assign n38678 =  ( n192 ) ? ( VREG_17_11 ) : ( VREG_17_11 ) ;
assign n38679 =  ( n157 ) ? ( n38677 ) : ( n38678 ) ;
assign n38680 =  ( n6 ) ? ( n38664 ) : ( n38679 ) ;
assign n38681 =  ( n373 ) ? ( n38680 ) : ( VREG_17_11 ) ;
assign n38682 =  ( n148 ) ? ( n10470 ) : ( VREG_17_12 ) ;
assign n38683 =  ( n146 ) ? ( n10469 ) : ( n38682 ) ;
assign n38684 =  ( n144 ) ? ( n10468 ) : ( n38683 ) ;
assign n38685 =  ( n142 ) ? ( n10467 ) : ( n38684 ) ;
assign n38686 =  ( n10 ) ? ( n10466 ) : ( n38685 ) ;
assign n38687 =  ( n148 ) ? ( n11504 ) : ( VREG_17_12 ) ;
assign n38688 =  ( n146 ) ? ( n11503 ) : ( n38687 ) ;
assign n38689 =  ( n144 ) ? ( n11502 ) : ( n38688 ) ;
assign n38690 =  ( n142 ) ? ( n11501 ) : ( n38689 ) ;
assign n38691 =  ( n10 ) ? ( n11500 ) : ( n38690 ) ;
assign n38692 =  ( n11511 ) ? ( VREG_17_12 ) : ( n38686 ) ;
assign n38693 =  ( n11511 ) ? ( VREG_17_12 ) : ( n38691 ) ;
assign n38694 =  ( n3034 ) ? ( n38693 ) : ( VREG_17_12 ) ;
assign n38695 =  ( n2965 ) ? ( n38692 ) : ( n38694 ) ;
assign n38696 =  ( n1930 ) ? ( n38691 ) : ( n38695 ) ;
assign n38697 =  ( n879 ) ? ( n38686 ) : ( n38696 ) ;
assign n38698 =  ( n172 ) ? ( n11522 ) : ( VREG_17_12 ) ;
assign n38699 =  ( n170 ) ? ( n11521 ) : ( n38698 ) ;
assign n38700 =  ( n168 ) ? ( n11520 ) : ( n38699 ) ;
assign n38701 =  ( n166 ) ? ( n11519 ) : ( n38700 ) ;
assign n38702 =  ( n162 ) ? ( n11518 ) : ( n38701 ) ;
assign n38703 =  ( n172 ) ? ( n11532 ) : ( VREG_17_12 ) ;
assign n38704 =  ( n170 ) ? ( n11531 ) : ( n38703 ) ;
assign n38705 =  ( n168 ) ? ( n11530 ) : ( n38704 ) ;
assign n38706 =  ( n166 ) ? ( n11529 ) : ( n38705 ) ;
assign n38707 =  ( n162 ) ? ( n11528 ) : ( n38706 ) ;
assign n38708 =  ( n11511 ) ? ( VREG_17_12 ) : ( n38707 ) ;
assign n38709 =  ( n3051 ) ? ( n38708 ) : ( VREG_17_12 ) ;
assign n38710 =  ( n3040 ) ? ( n38702 ) : ( n38709 ) ;
assign n38711 =  ( n192 ) ? ( VREG_17_12 ) : ( VREG_17_12 ) ;
assign n38712 =  ( n157 ) ? ( n38710 ) : ( n38711 ) ;
assign n38713 =  ( n6 ) ? ( n38697 ) : ( n38712 ) ;
assign n38714 =  ( n373 ) ? ( n38713 ) : ( VREG_17_12 ) ;
assign n38715 =  ( n148 ) ? ( n12589 ) : ( VREG_17_13 ) ;
assign n38716 =  ( n146 ) ? ( n12588 ) : ( n38715 ) ;
assign n38717 =  ( n144 ) ? ( n12587 ) : ( n38716 ) ;
assign n38718 =  ( n142 ) ? ( n12586 ) : ( n38717 ) ;
assign n38719 =  ( n10 ) ? ( n12585 ) : ( n38718 ) ;
assign n38720 =  ( n148 ) ? ( n13623 ) : ( VREG_17_13 ) ;
assign n38721 =  ( n146 ) ? ( n13622 ) : ( n38720 ) ;
assign n38722 =  ( n144 ) ? ( n13621 ) : ( n38721 ) ;
assign n38723 =  ( n142 ) ? ( n13620 ) : ( n38722 ) ;
assign n38724 =  ( n10 ) ? ( n13619 ) : ( n38723 ) ;
assign n38725 =  ( n13630 ) ? ( VREG_17_13 ) : ( n38719 ) ;
assign n38726 =  ( n13630 ) ? ( VREG_17_13 ) : ( n38724 ) ;
assign n38727 =  ( n3034 ) ? ( n38726 ) : ( VREG_17_13 ) ;
assign n38728 =  ( n2965 ) ? ( n38725 ) : ( n38727 ) ;
assign n38729 =  ( n1930 ) ? ( n38724 ) : ( n38728 ) ;
assign n38730 =  ( n879 ) ? ( n38719 ) : ( n38729 ) ;
assign n38731 =  ( n172 ) ? ( n13641 ) : ( VREG_17_13 ) ;
assign n38732 =  ( n170 ) ? ( n13640 ) : ( n38731 ) ;
assign n38733 =  ( n168 ) ? ( n13639 ) : ( n38732 ) ;
assign n38734 =  ( n166 ) ? ( n13638 ) : ( n38733 ) ;
assign n38735 =  ( n162 ) ? ( n13637 ) : ( n38734 ) ;
assign n38736 =  ( n172 ) ? ( n13651 ) : ( VREG_17_13 ) ;
assign n38737 =  ( n170 ) ? ( n13650 ) : ( n38736 ) ;
assign n38738 =  ( n168 ) ? ( n13649 ) : ( n38737 ) ;
assign n38739 =  ( n166 ) ? ( n13648 ) : ( n38738 ) ;
assign n38740 =  ( n162 ) ? ( n13647 ) : ( n38739 ) ;
assign n38741 =  ( n13630 ) ? ( VREG_17_13 ) : ( n38740 ) ;
assign n38742 =  ( n3051 ) ? ( n38741 ) : ( VREG_17_13 ) ;
assign n38743 =  ( n3040 ) ? ( n38735 ) : ( n38742 ) ;
assign n38744 =  ( n192 ) ? ( VREG_17_13 ) : ( VREG_17_13 ) ;
assign n38745 =  ( n157 ) ? ( n38743 ) : ( n38744 ) ;
assign n38746 =  ( n6 ) ? ( n38730 ) : ( n38745 ) ;
assign n38747 =  ( n373 ) ? ( n38746 ) : ( VREG_17_13 ) ;
assign n38748 =  ( n148 ) ? ( n14708 ) : ( VREG_17_14 ) ;
assign n38749 =  ( n146 ) ? ( n14707 ) : ( n38748 ) ;
assign n38750 =  ( n144 ) ? ( n14706 ) : ( n38749 ) ;
assign n38751 =  ( n142 ) ? ( n14705 ) : ( n38750 ) ;
assign n38752 =  ( n10 ) ? ( n14704 ) : ( n38751 ) ;
assign n38753 =  ( n148 ) ? ( n15742 ) : ( VREG_17_14 ) ;
assign n38754 =  ( n146 ) ? ( n15741 ) : ( n38753 ) ;
assign n38755 =  ( n144 ) ? ( n15740 ) : ( n38754 ) ;
assign n38756 =  ( n142 ) ? ( n15739 ) : ( n38755 ) ;
assign n38757 =  ( n10 ) ? ( n15738 ) : ( n38756 ) ;
assign n38758 =  ( n15749 ) ? ( VREG_17_14 ) : ( n38752 ) ;
assign n38759 =  ( n15749 ) ? ( VREG_17_14 ) : ( n38757 ) ;
assign n38760 =  ( n3034 ) ? ( n38759 ) : ( VREG_17_14 ) ;
assign n38761 =  ( n2965 ) ? ( n38758 ) : ( n38760 ) ;
assign n38762 =  ( n1930 ) ? ( n38757 ) : ( n38761 ) ;
assign n38763 =  ( n879 ) ? ( n38752 ) : ( n38762 ) ;
assign n38764 =  ( n172 ) ? ( n15760 ) : ( VREG_17_14 ) ;
assign n38765 =  ( n170 ) ? ( n15759 ) : ( n38764 ) ;
assign n38766 =  ( n168 ) ? ( n15758 ) : ( n38765 ) ;
assign n38767 =  ( n166 ) ? ( n15757 ) : ( n38766 ) ;
assign n38768 =  ( n162 ) ? ( n15756 ) : ( n38767 ) ;
assign n38769 =  ( n172 ) ? ( n15770 ) : ( VREG_17_14 ) ;
assign n38770 =  ( n170 ) ? ( n15769 ) : ( n38769 ) ;
assign n38771 =  ( n168 ) ? ( n15768 ) : ( n38770 ) ;
assign n38772 =  ( n166 ) ? ( n15767 ) : ( n38771 ) ;
assign n38773 =  ( n162 ) ? ( n15766 ) : ( n38772 ) ;
assign n38774 =  ( n15749 ) ? ( VREG_17_14 ) : ( n38773 ) ;
assign n38775 =  ( n3051 ) ? ( n38774 ) : ( VREG_17_14 ) ;
assign n38776 =  ( n3040 ) ? ( n38768 ) : ( n38775 ) ;
assign n38777 =  ( n192 ) ? ( VREG_17_14 ) : ( VREG_17_14 ) ;
assign n38778 =  ( n157 ) ? ( n38776 ) : ( n38777 ) ;
assign n38779 =  ( n6 ) ? ( n38763 ) : ( n38778 ) ;
assign n38780 =  ( n373 ) ? ( n38779 ) : ( VREG_17_14 ) ;
assign n38781 =  ( n148 ) ? ( n16827 ) : ( VREG_17_15 ) ;
assign n38782 =  ( n146 ) ? ( n16826 ) : ( n38781 ) ;
assign n38783 =  ( n144 ) ? ( n16825 ) : ( n38782 ) ;
assign n38784 =  ( n142 ) ? ( n16824 ) : ( n38783 ) ;
assign n38785 =  ( n10 ) ? ( n16823 ) : ( n38784 ) ;
assign n38786 =  ( n148 ) ? ( n17861 ) : ( VREG_17_15 ) ;
assign n38787 =  ( n146 ) ? ( n17860 ) : ( n38786 ) ;
assign n38788 =  ( n144 ) ? ( n17859 ) : ( n38787 ) ;
assign n38789 =  ( n142 ) ? ( n17858 ) : ( n38788 ) ;
assign n38790 =  ( n10 ) ? ( n17857 ) : ( n38789 ) ;
assign n38791 =  ( n17868 ) ? ( VREG_17_15 ) : ( n38785 ) ;
assign n38792 =  ( n17868 ) ? ( VREG_17_15 ) : ( n38790 ) ;
assign n38793 =  ( n3034 ) ? ( n38792 ) : ( VREG_17_15 ) ;
assign n38794 =  ( n2965 ) ? ( n38791 ) : ( n38793 ) ;
assign n38795 =  ( n1930 ) ? ( n38790 ) : ( n38794 ) ;
assign n38796 =  ( n879 ) ? ( n38785 ) : ( n38795 ) ;
assign n38797 =  ( n172 ) ? ( n17879 ) : ( VREG_17_15 ) ;
assign n38798 =  ( n170 ) ? ( n17878 ) : ( n38797 ) ;
assign n38799 =  ( n168 ) ? ( n17877 ) : ( n38798 ) ;
assign n38800 =  ( n166 ) ? ( n17876 ) : ( n38799 ) ;
assign n38801 =  ( n162 ) ? ( n17875 ) : ( n38800 ) ;
assign n38802 =  ( n172 ) ? ( n17889 ) : ( VREG_17_15 ) ;
assign n38803 =  ( n170 ) ? ( n17888 ) : ( n38802 ) ;
assign n38804 =  ( n168 ) ? ( n17887 ) : ( n38803 ) ;
assign n38805 =  ( n166 ) ? ( n17886 ) : ( n38804 ) ;
assign n38806 =  ( n162 ) ? ( n17885 ) : ( n38805 ) ;
assign n38807 =  ( n17868 ) ? ( VREG_17_15 ) : ( n38806 ) ;
assign n38808 =  ( n3051 ) ? ( n38807 ) : ( VREG_17_15 ) ;
assign n38809 =  ( n3040 ) ? ( n38801 ) : ( n38808 ) ;
assign n38810 =  ( n192 ) ? ( VREG_17_15 ) : ( VREG_17_15 ) ;
assign n38811 =  ( n157 ) ? ( n38809 ) : ( n38810 ) ;
assign n38812 =  ( n6 ) ? ( n38796 ) : ( n38811 ) ;
assign n38813 =  ( n373 ) ? ( n38812 ) : ( VREG_17_15 ) ;
assign n38814 =  ( n148 ) ? ( n18946 ) : ( VREG_17_2 ) ;
assign n38815 =  ( n146 ) ? ( n18945 ) : ( n38814 ) ;
assign n38816 =  ( n144 ) ? ( n18944 ) : ( n38815 ) ;
assign n38817 =  ( n142 ) ? ( n18943 ) : ( n38816 ) ;
assign n38818 =  ( n10 ) ? ( n18942 ) : ( n38817 ) ;
assign n38819 =  ( n148 ) ? ( n19980 ) : ( VREG_17_2 ) ;
assign n38820 =  ( n146 ) ? ( n19979 ) : ( n38819 ) ;
assign n38821 =  ( n144 ) ? ( n19978 ) : ( n38820 ) ;
assign n38822 =  ( n142 ) ? ( n19977 ) : ( n38821 ) ;
assign n38823 =  ( n10 ) ? ( n19976 ) : ( n38822 ) ;
assign n38824 =  ( n19987 ) ? ( VREG_17_2 ) : ( n38818 ) ;
assign n38825 =  ( n19987 ) ? ( VREG_17_2 ) : ( n38823 ) ;
assign n38826 =  ( n3034 ) ? ( n38825 ) : ( VREG_17_2 ) ;
assign n38827 =  ( n2965 ) ? ( n38824 ) : ( n38826 ) ;
assign n38828 =  ( n1930 ) ? ( n38823 ) : ( n38827 ) ;
assign n38829 =  ( n879 ) ? ( n38818 ) : ( n38828 ) ;
assign n38830 =  ( n172 ) ? ( n19998 ) : ( VREG_17_2 ) ;
assign n38831 =  ( n170 ) ? ( n19997 ) : ( n38830 ) ;
assign n38832 =  ( n168 ) ? ( n19996 ) : ( n38831 ) ;
assign n38833 =  ( n166 ) ? ( n19995 ) : ( n38832 ) ;
assign n38834 =  ( n162 ) ? ( n19994 ) : ( n38833 ) ;
assign n38835 =  ( n172 ) ? ( n20008 ) : ( VREG_17_2 ) ;
assign n38836 =  ( n170 ) ? ( n20007 ) : ( n38835 ) ;
assign n38837 =  ( n168 ) ? ( n20006 ) : ( n38836 ) ;
assign n38838 =  ( n166 ) ? ( n20005 ) : ( n38837 ) ;
assign n38839 =  ( n162 ) ? ( n20004 ) : ( n38838 ) ;
assign n38840 =  ( n19987 ) ? ( VREG_17_2 ) : ( n38839 ) ;
assign n38841 =  ( n3051 ) ? ( n38840 ) : ( VREG_17_2 ) ;
assign n38842 =  ( n3040 ) ? ( n38834 ) : ( n38841 ) ;
assign n38843 =  ( n192 ) ? ( VREG_17_2 ) : ( VREG_17_2 ) ;
assign n38844 =  ( n157 ) ? ( n38842 ) : ( n38843 ) ;
assign n38845 =  ( n6 ) ? ( n38829 ) : ( n38844 ) ;
assign n38846 =  ( n373 ) ? ( n38845 ) : ( VREG_17_2 ) ;
assign n38847 =  ( n148 ) ? ( n21065 ) : ( VREG_17_3 ) ;
assign n38848 =  ( n146 ) ? ( n21064 ) : ( n38847 ) ;
assign n38849 =  ( n144 ) ? ( n21063 ) : ( n38848 ) ;
assign n38850 =  ( n142 ) ? ( n21062 ) : ( n38849 ) ;
assign n38851 =  ( n10 ) ? ( n21061 ) : ( n38850 ) ;
assign n38852 =  ( n148 ) ? ( n22099 ) : ( VREG_17_3 ) ;
assign n38853 =  ( n146 ) ? ( n22098 ) : ( n38852 ) ;
assign n38854 =  ( n144 ) ? ( n22097 ) : ( n38853 ) ;
assign n38855 =  ( n142 ) ? ( n22096 ) : ( n38854 ) ;
assign n38856 =  ( n10 ) ? ( n22095 ) : ( n38855 ) ;
assign n38857 =  ( n22106 ) ? ( VREG_17_3 ) : ( n38851 ) ;
assign n38858 =  ( n22106 ) ? ( VREG_17_3 ) : ( n38856 ) ;
assign n38859 =  ( n3034 ) ? ( n38858 ) : ( VREG_17_3 ) ;
assign n38860 =  ( n2965 ) ? ( n38857 ) : ( n38859 ) ;
assign n38861 =  ( n1930 ) ? ( n38856 ) : ( n38860 ) ;
assign n38862 =  ( n879 ) ? ( n38851 ) : ( n38861 ) ;
assign n38863 =  ( n172 ) ? ( n22117 ) : ( VREG_17_3 ) ;
assign n38864 =  ( n170 ) ? ( n22116 ) : ( n38863 ) ;
assign n38865 =  ( n168 ) ? ( n22115 ) : ( n38864 ) ;
assign n38866 =  ( n166 ) ? ( n22114 ) : ( n38865 ) ;
assign n38867 =  ( n162 ) ? ( n22113 ) : ( n38866 ) ;
assign n38868 =  ( n172 ) ? ( n22127 ) : ( VREG_17_3 ) ;
assign n38869 =  ( n170 ) ? ( n22126 ) : ( n38868 ) ;
assign n38870 =  ( n168 ) ? ( n22125 ) : ( n38869 ) ;
assign n38871 =  ( n166 ) ? ( n22124 ) : ( n38870 ) ;
assign n38872 =  ( n162 ) ? ( n22123 ) : ( n38871 ) ;
assign n38873 =  ( n22106 ) ? ( VREG_17_3 ) : ( n38872 ) ;
assign n38874 =  ( n3051 ) ? ( n38873 ) : ( VREG_17_3 ) ;
assign n38875 =  ( n3040 ) ? ( n38867 ) : ( n38874 ) ;
assign n38876 =  ( n192 ) ? ( VREG_17_3 ) : ( VREG_17_3 ) ;
assign n38877 =  ( n157 ) ? ( n38875 ) : ( n38876 ) ;
assign n38878 =  ( n6 ) ? ( n38862 ) : ( n38877 ) ;
assign n38879 =  ( n373 ) ? ( n38878 ) : ( VREG_17_3 ) ;
assign n38880 =  ( n148 ) ? ( n23184 ) : ( VREG_17_4 ) ;
assign n38881 =  ( n146 ) ? ( n23183 ) : ( n38880 ) ;
assign n38882 =  ( n144 ) ? ( n23182 ) : ( n38881 ) ;
assign n38883 =  ( n142 ) ? ( n23181 ) : ( n38882 ) ;
assign n38884 =  ( n10 ) ? ( n23180 ) : ( n38883 ) ;
assign n38885 =  ( n148 ) ? ( n24218 ) : ( VREG_17_4 ) ;
assign n38886 =  ( n146 ) ? ( n24217 ) : ( n38885 ) ;
assign n38887 =  ( n144 ) ? ( n24216 ) : ( n38886 ) ;
assign n38888 =  ( n142 ) ? ( n24215 ) : ( n38887 ) ;
assign n38889 =  ( n10 ) ? ( n24214 ) : ( n38888 ) ;
assign n38890 =  ( n24225 ) ? ( VREG_17_4 ) : ( n38884 ) ;
assign n38891 =  ( n24225 ) ? ( VREG_17_4 ) : ( n38889 ) ;
assign n38892 =  ( n3034 ) ? ( n38891 ) : ( VREG_17_4 ) ;
assign n38893 =  ( n2965 ) ? ( n38890 ) : ( n38892 ) ;
assign n38894 =  ( n1930 ) ? ( n38889 ) : ( n38893 ) ;
assign n38895 =  ( n879 ) ? ( n38884 ) : ( n38894 ) ;
assign n38896 =  ( n172 ) ? ( n24236 ) : ( VREG_17_4 ) ;
assign n38897 =  ( n170 ) ? ( n24235 ) : ( n38896 ) ;
assign n38898 =  ( n168 ) ? ( n24234 ) : ( n38897 ) ;
assign n38899 =  ( n166 ) ? ( n24233 ) : ( n38898 ) ;
assign n38900 =  ( n162 ) ? ( n24232 ) : ( n38899 ) ;
assign n38901 =  ( n172 ) ? ( n24246 ) : ( VREG_17_4 ) ;
assign n38902 =  ( n170 ) ? ( n24245 ) : ( n38901 ) ;
assign n38903 =  ( n168 ) ? ( n24244 ) : ( n38902 ) ;
assign n38904 =  ( n166 ) ? ( n24243 ) : ( n38903 ) ;
assign n38905 =  ( n162 ) ? ( n24242 ) : ( n38904 ) ;
assign n38906 =  ( n24225 ) ? ( VREG_17_4 ) : ( n38905 ) ;
assign n38907 =  ( n3051 ) ? ( n38906 ) : ( VREG_17_4 ) ;
assign n38908 =  ( n3040 ) ? ( n38900 ) : ( n38907 ) ;
assign n38909 =  ( n192 ) ? ( VREG_17_4 ) : ( VREG_17_4 ) ;
assign n38910 =  ( n157 ) ? ( n38908 ) : ( n38909 ) ;
assign n38911 =  ( n6 ) ? ( n38895 ) : ( n38910 ) ;
assign n38912 =  ( n373 ) ? ( n38911 ) : ( VREG_17_4 ) ;
assign n38913 =  ( n148 ) ? ( n25303 ) : ( VREG_17_5 ) ;
assign n38914 =  ( n146 ) ? ( n25302 ) : ( n38913 ) ;
assign n38915 =  ( n144 ) ? ( n25301 ) : ( n38914 ) ;
assign n38916 =  ( n142 ) ? ( n25300 ) : ( n38915 ) ;
assign n38917 =  ( n10 ) ? ( n25299 ) : ( n38916 ) ;
assign n38918 =  ( n148 ) ? ( n26337 ) : ( VREG_17_5 ) ;
assign n38919 =  ( n146 ) ? ( n26336 ) : ( n38918 ) ;
assign n38920 =  ( n144 ) ? ( n26335 ) : ( n38919 ) ;
assign n38921 =  ( n142 ) ? ( n26334 ) : ( n38920 ) ;
assign n38922 =  ( n10 ) ? ( n26333 ) : ( n38921 ) ;
assign n38923 =  ( n26344 ) ? ( VREG_17_5 ) : ( n38917 ) ;
assign n38924 =  ( n26344 ) ? ( VREG_17_5 ) : ( n38922 ) ;
assign n38925 =  ( n3034 ) ? ( n38924 ) : ( VREG_17_5 ) ;
assign n38926 =  ( n2965 ) ? ( n38923 ) : ( n38925 ) ;
assign n38927 =  ( n1930 ) ? ( n38922 ) : ( n38926 ) ;
assign n38928 =  ( n879 ) ? ( n38917 ) : ( n38927 ) ;
assign n38929 =  ( n172 ) ? ( n26355 ) : ( VREG_17_5 ) ;
assign n38930 =  ( n170 ) ? ( n26354 ) : ( n38929 ) ;
assign n38931 =  ( n168 ) ? ( n26353 ) : ( n38930 ) ;
assign n38932 =  ( n166 ) ? ( n26352 ) : ( n38931 ) ;
assign n38933 =  ( n162 ) ? ( n26351 ) : ( n38932 ) ;
assign n38934 =  ( n172 ) ? ( n26365 ) : ( VREG_17_5 ) ;
assign n38935 =  ( n170 ) ? ( n26364 ) : ( n38934 ) ;
assign n38936 =  ( n168 ) ? ( n26363 ) : ( n38935 ) ;
assign n38937 =  ( n166 ) ? ( n26362 ) : ( n38936 ) ;
assign n38938 =  ( n162 ) ? ( n26361 ) : ( n38937 ) ;
assign n38939 =  ( n26344 ) ? ( VREG_17_5 ) : ( n38938 ) ;
assign n38940 =  ( n3051 ) ? ( n38939 ) : ( VREG_17_5 ) ;
assign n38941 =  ( n3040 ) ? ( n38933 ) : ( n38940 ) ;
assign n38942 =  ( n192 ) ? ( VREG_17_5 ) : ( VREG_17_5 ) ;
assign n38943 =  ( n157 ) ? ( n38941 ) : ( n38942 ) ;
assign n38944 =  ( n6 ) ? ( n38928 ) : ( n38943 ) ;
assign n38945 =  ( n373 ) ? ( n38944 ) : ( VREG_17_5 ) ;
assign n38946 =  ( n148 ) ? ( n27422 ) : ( VREG_17_6 ) ;
assign n38947 =  ( n146 ) ? ( n27421 ) : ( n38946 ) ;
assign n38948 =  ( n144 ) ? ( n27420 ) : ( n38947 ) ;
assign n38949 =  ( n142 ) ? ( n27419 ) : ( n38948 ) ;
assign n38950 =  ( n10 ) ? ( n27418 ) : ( n38949 ) ;
assign n38951 =  ( n148 ) ? ( n28456 ) : ( VREG_17_6 ) ;
assign n38952 =  ( n146 ) ? ( n28455 ) : ( n38951 ) ;
assign n38953 =  ( n144 ) ? ( n28454 ) : ( n38952 ) ;
assign n38954 =  ( n142 ) ? ( n28453 ) : ( n38953 ) ;
assign n38955 =  ( n10 ) ? ( n28452 ) : ( n38954 ) ;
assign n38956 =  ( n28463 ) ? ( VREG_17_6 ) : ( n38950 ) ;
assign n38957 =  ( n28463 ) ? ( VREG_17_6 ) : ( n38955 ) ;
assign n38958 =  ( n3034 ) ? ( n38957 ) : ( VREG_17_6 ) ;
assign n38959 =  ( n2965 ) ? ( n38956 ) : ( n38958 ) ;
assign n38960 =  ( n1930 ) ? ( n38955 ) : ( n38959 ) ;
assign n38961 =  ( n879 ) ? ( n38950 ) : ( n38960 ) ;
assign n38962 =  ( n172 ) ? ( n28474 ) : ( VREG_17_6 ) ;
assign n38963 =  ( n170 ) ? ( n28473 ) : ( n38962 ) ;
assign n38964 =  ( n168 ) ? ( n28472 ) : ( n38963 ) ;
assign n38965 =  ( n166 ) ? ( n28471 ) : ( n38964 ) ;
assign n38966 =  ( n162 ) ? ( n28470 ) : ( n38965 ) ;
assign n38967 =  ( n172 ) ? ( n28484 ) : ( VREG_17_6 ) ;
assign n38968 =  ( n170 ) ? ( n28483 ) : ( n38967 ) ;
assign n38969 =  ( n168 ) ? ( n28482 ) : ( n38968 ) ;
assign n38970 =  ( n166 ) ? ( n28481 ) : ( n38969 ) ;
assign n38971 =  ( n162 ) ? ( n28480 ) : ( n38970 ) ;
assign n38972 =  ( n28463 ) ? ( VREG_17_6 ) : ( n38971 ) ;
assign n38973 =  ( n3051 ) ? ( n38972 ) : ( VREG_17_6 ) ;
assign n38974 =  ( n3040 ) ? ( n38966 ) : ( n38973 ) ;
assign n38975 =  ( n192 ) ? ( VREG_17_6 ) : ( VREG_17_6 ) ;
assign n38976 =  ( n157 ) ? ( n38974 ) : ( n38975 ) ;
assign n38977 =  ( n6 ) ? ( n38961 ) : ( n38976 ) ;
assign n38978 =  ( n373 ) ? ( n38977 ) : ( VREG_17_6 ) ;
assign n38979 =  ( n148 ) ? ( n29541 ) : ( VREG_17_7 ) ;
assign n38980 =  ( n146 ) ? ( n29540 ) : ( n38979 ) ;
assign n38981 =  ( n144 ) ? ( n29539 ) : ( n38980 ) ;
assign n38982 =  ( n142 ) ? ( n29538 ) : ( n38981 ) ;
assign n38983 =  ( n10 ) ? ( n29537 ) : ( n38982 ) ;
assign n38984 =  ( n148 ) ? ( n30575 ) : ( VREG_17_7 ) ;
assign n38985 =  ( n146 ) ? ( n30574 ) : ( n38984 ) ;
assign n38986 =  ( n144 ) ? ( n30573 ) : ( n38985 ) ;
assign n38987 =  ( n142 ) ? ( n30572 ) : ( n38986 ) ;
assign n38988 =  ( n10 ) ? ( n30571 ) : ( n38987 ) ;
assign n38989 =  ( n30582 ) ? ( VREG_17_7 ) : ( n38983 ) ;
assign n38990 =  ( n30582 ) ? ( VREG_17_7 ) : ( n38988 ) ;
assign n38991 =  ( n3034 ) ? ( n38990 ) : ( VREG_17_7 ) ;
assign n38992 =  ( n2965 ) ? ( n38989 ) : ( n38991 ) ;
assign n38993 =  ( n1930 ) ? ( n38988 ) : ( n38992 ) ;
assign n38994 =  ( n879 ) ? ( n38983 ) : ( n38993 ) ;
assign n38995 =  ( n172 ) ? ( n30593 ) : ( VREG_17_7 ) ;
assign n38996 =  ( n170 ) ? ( n30592 ) : ( n38995 ) ;
assign n38997 =  ( n168 ) ? ( n30591 ) : ( n38996 ) ;
assign n38998 =  ( n166 ) ? ( n30590 ) : ( n38997 ) ;
assign n38999 =  ( n162 ) ? ( n30589 ) : ( n38998 ) ;
assign n39000 =  ( n172 ) ? ( n30603 ) : ( VREG_17_7 ) ;
assign n39001 =  ( n170 ) ? ( n30602 ) : ( n39000 ) ;
assign n39002 =  ( n168 ) ? ( n30601 ) : ( n39001 ) ;
assign n39003 =  ( n166 ) ? ( n30600 ) : ( n39002 ) ;
assign n39004 =  ( n162 ) ? ( n30599 ) : ( n39003 ) ;
assign n39005 =  ( n30582 ) ? ( VREG_17_7 ) : ( n39004 ) ;
assign n39006 =  ( n3051 ) ? ( n39005 ) : ( VREG_17_7 ) ;
assign n39007 =  ( n3040 ) ? ( n38999 ) : ( n39006 ) ;
assign n39008 =  ( n192 ) ? ( VREG_17_7 ) : ( VREG_17_7 ) ;
assign n39009 =  ( n157 ) ? ( n39007 ) : ( n39008 ) ;
assign n39010 =  ( n6 ) ? ( n38994 ) : ( n39009 ) ;
assign n39011 =  ( n373 ) ? ( n39010 ) : ( VREG_17_7 ) ;
assign n39012 =  ( n148 ) ? ( n31660 ) : ( VREG_17_8 ) ;
assign n39013 =  ( n146 ) ? ( n31659 ) : ( n39012 ) ;
assign n39014 =  ( n144 ) ? ( n31658 ) : ( n39013 ) ;
assign n39015 =  ( n142 ) ? ( n31657 ) : ( n39014 ) ;
assign n39016 =  ( n10 ) ? ( n31656 ) : ( n39015 ) ;
assign n39017 =  ( n148 ) ? ( n32694 ) : ( VREG_17_8 ) ;
assign n39018 =  ( n146 ) ? ( n32693 ) : ( n39017 ) ;
assign n39019 =  ( n144 ) ? ( n32692 ) : ( n39018 ) ;
assign n39020 =  ( n142 ) ? ( n32691 ) : ( n39019 ) ;
assign n39021 =  ( n10 ) ? ( n32690 ) : ( n39020 ) ;
assign n39022 =  ( n32701 ) ? ( VREG_17_8 ) : ( n39016 ) ;
assign n39023 =  ( n32701 ) ? ( VREG_17_8 ) : ( n39021 ) ;
assign n39024 =  ( n3034 ) ? ( n39023 ) : ( VREG_17_8 ) ;
assign n39025 =  ( n2965 ) ? ( n39022 ) : ( n39024 ) ;
assign n39026 =  ( n1930 ) ? ( n39021 ) : ( n39025 ) ;
assign n39027 =  ( n879 ) ? ( n39016 ) : ( n39026 ) ;
assign n39028 =  ( n172 ) ? ( n32712 ) : ( VREG_17_8 ) ;
assign n39029 =  ( n170 ) ? ( n32711 ) : ( n39028 ) ;
assign n39030 =  ( n168 ) ? ( n32710 ) : ( n39029 ) ;
assign n39031 =  ( n166 ) ? ( n32709 ) : ( n39030 ) ;
assign n39032 =  ( n162 ) ? ( n32708 ) : ( n39031 ) ;
assign n39033 =  ( n172 ) ? ( n32722 ) : ( VREG_17_8 ) ;
assign n39034 =  ( n170 ) ? ( n32721 ) : ( n39033 ) ;
assign n39035 =  ( n168 ) ? ( n32720 ) : ( n39034 ) ;
assign n39036 =  ( n166 ) ? ( n32719 ) : ( n39035 ) ;
assign n39037 =  ( n162 ) ? ( n32718 ) : ( n39036 ) ;
assign n39038 =  ( n32701 ) ? ( VREG_17_8 ) : ( n39037 ) ;
assign n39039 =  ( n3051 ) ? ( n39038 ) : ( VREG_17_8 ) ;
assign n39040 =  ( n3040 ) ? ( n39032 ) : ( n39039 ) ;
assign n39041 =  ( n192 ) ? ( VREG_17_8 ) : ( VREG_17_8 ) ;
assign n39042 =  ( n157 ) ? ( n39040 ) : ( n39041 ) ;
assign n39043 =  ( n6 ) ? ( n39027 ) : ( n39042 ) ;
assign n39044 =  ( n373 ) ? ( n39043 ) : ( VREG_17_8 ) ;
assign n39045 =  ( n148 ) ? ( n33779 ) : ( VREG_17_9 ) ;
assign n39046 =  ( n146 ) ? ( n33778 ) : ( n39045 ) ;
assign n39047 =  ( n144 ) ? ( n33777 ) : ( n39046 ) ;
assign n39048 =  ( n142 ) ? ( n33776 ) : ( n39047 ) ;
assign n39049 =  ( n10 ) ? ( n33775 ) : ( n39048 ) ;
assign n39050 =  ( n148 ) ? ( n34813 ) : ( VREG_17_9 ) ;
assign n39051 =  ( n146 ) ? ( n34812 ) : ( n39050 ) ;
assign n39052 =  ( n144 ) ? ( n34811 ) : ( n39051 ) ;
assign n39053 =  ( n142 ) ? ( n34810 ) : ( n39052 ) ;
assign n39054 =  ( n10 ) ? ( n34809 ) : ( n39053 ) ;
assign n39055 =  ( n34820 ) ? ( VREG_17_9 ) : ( n39049 ) ;
assign n39056 =  ( n34820 ) ? ( VREG_17_9 ) : ( n39054 ) ;
assign n39057 =  ( n3034 ) ? ( n39056 ) : ( VREG_17_9 ) ;
assign n39058 =  ( n2965 ) ? ( n39055 ) : ( n39057 ) ;
assign n39059 =  ( n1930 ) ? ( n39054 ) : ( n39058 ) ;
assign n39060 =  ( n879 ) ? ( n39049 ) : ( n39059 ) ;
assign n39061 =  ( n172 ) ? ( n34831 ) : ( VREG_17_9 ) ;
assign n39062 =  ( n170 ) ? ( n34830 ) : ( n39061 ) ;
assign n39063 =  ( n168 ) ? ( n34829 ) : ( n39062 ) ;
assign n39064 =  ( n166 ) ? ( n34828 ) : ( n39063 ) ;
assign n39065 =  ( n162 ) ? ( n34827 ) : ( n39064 ) ;
assign n39066 =  ( n172 ) ? ( n34841 ) : ( VREG_17_9 ) ;
assign n39067 =  ( n170 ) ? ( n34840 ) : ( n39066 ) ;
assign n39068 =  ( n168 ) ? ( n34839 ) : ( n39067 ) ;
assign n39069 =  ( n166 ) ? ( n34838 ) : ( n39068 ) ;
assign n39070 =  ( n162 ) ? ( n34837 ) : ( n39069 ) ;
assign n39071 =  ( n34820 ) ? ( VREG_17_9 ) : ( n39070 ) ;
assign n39072 =  ( n3051 ) ? ( n39071 ) : ( VREG_17_9 ) ;
assign n39073 =  ( n3040 ) ? ( n39065 ) : ( n39072 ) ;
assign n39074 =  ( n192 ) ? ( VREG_17_9 ) : ( VREG_17_9 ) ;
assign n39075 =  ( n157 ) ? ( n39073 ) : ( n39074 ) ;
assign n39076 =  ( n6 ) ? ( n39060 ) : ( n39075 ) ;
assign n39077 =  ( n373 ) ? ( n39076 ) : ( VREG_17_9 ) ;
assign n39078 =  ( n148 ) ? ( n1924 ) : ( VREG_18_0 ) ;
assign n39079 =  ( n146 ) ? ( n1923 ) : ( n39078 ) ;
assign n39080 =  ( n144 ) ? ( n1922 ) : ( n39079 ) ;
assign n39081 =  ( n142 ) ? ( n1921 ) : ( n39080 ) ;
assign n39082 =  ( n10 ) ? ( n1920 ) : ( n39081 ) ;
assign n39083 =  ( n148 ) ? ( n2959 ) : ( VREG_18_0 ) ;
assign n39084 =  ( n146 ) ? ( n2958 ) : ( n39083 ) ;
assign n39085 =  ( n144 ) ? ( n2957 ) : ( n39084 ) ;
assign n39086 =  ( n142 ) ? ( n2956 ) : ( n39085 ) ;
assign n39087 =  ( n10 ) ? ( n2955 ) : ( n39086 ) ;
assign n39088 =  ( n3032 ) ? ( VREG_18_0 ) : ( n39082 ) ;
assign n39089 =  ( n3032 ) ? ( VREG_18_0 ) : ( n39087 ) ;
assign n39090 =  ( n3034 ) ? ( n39089 ) : ( VREG_18_0 ) ;
assign n39091 =  ( n2965 ) ? ( n39088 ) : ( n39090 ) ;
assign n39092 =  ( n1930 ) ? ( n39087 ) : ( n39091 ) ;
assign n39093 =  ( n879 ) ? ( n39082 ) : ( n39092 ) ;
assign n39094 =  ( n172 ) ? ( n3045 ) : ( VREG_18_0 ) ;
assign n39095 =  ( n170 ) ? ( n3044 ) : ( n39094 ) ;
assign n39096 =  ( n168 ) ? ( n3043 ) : ( n39095 ) ;
assign n39097 =  ( n166 ) ? ( n3042 ) : ( n39096 ) ;
assign n39098 =  ( n162 ) ? ( n3041 ) : ( n39097 ) ;
assign n39099 =  ( n172 ) ? ( n3056 ) : ( VREG_18_0 ) ;
assign n39100 =  ( n170 ) ? ( n3055 ) : ( n39099 ) ;
assign n39101 =  ( n168 ) ? ( n3054 ) : ( n39100 ) ;
assign n39102 =  ( n166 ) ? ( n3053 ) : ( n39101 ) ;
assign n39103 =  ( n162 ) ? ( n3052 ) : ( n39102 ) ;
assign n39104 =  ( n3032 ) ? ( VREG_18_0 ) : ( n39103 ) ;
assign n39105 =  ( n3051 ) ? ( n39104 ) : ( VREG_18_0 ) ;
assign n39106 =  ( n3040 ) ? ( n39098 ) : ( n39105 ) ;
assign n39107 =  ( n192 ) ? ( VREG_18_0 ) : ( VREG_18_0 ) ;
assign n39108 =  ( n157 ) ? ( n39106 ) : ( n39107 ) ;
assign n39109 =  ( n6 ) ? ( n39093 ) : ( n39108 ) ;
assign n39110 =  ( n395 ) ? ( n39109 ) : ( VREG_18_0 ) ;
assign n39111 =  ( n148 ) ? ( n4113 ) : ( VREG_18_1 ) ;
assign n39112 =  ( n146 ) ? ( n4112 ) : ( n39111 ) ;
assign n39113 =  ( n144 ) ? ( n4111 ) : ( n39112 ) ;
assign n39114 =  ( n142 ) ? ( n4110 ) : ( n39113 ) ;
assign n39115 =  ( n10 ) ? ( n4109 ) : ( n39114 ) ;
assign n39116 =  ( n148 ) ? ( n5147 ) : ( VREG_18_1 ) ;
assign n39117 =  ( n146 ) ? ( n5146 ) : ( n39116 ) ;
assign n39118 =  ( n144 ) ? ( n5145 ) : ( n39117 ) ;
assign n39119 =  ( n142 ) ? ( n5144 ) : ( n39118 ) ;
assign n39120 =  ( n10 ) ? ( n5143 ) : ( n39119 ) ;
assign n39121 =  ( n5154 ) ? ( VREG_18_1 ) : ( n39115 ) ;
assign n39122 =  ( n5154 ) ? ( VREG_18_1 ) : ( n39120 ) ;
assign n39123 =  ( n3034 ) ? ( n39122 ) : ( VREG_18_1 ) ;
assign n39124 =  ( n2965 ) ? ( n39121 ) : ( n39123 ) ;
assign n39125 =  ( n1930 ) ? ( n39120 ) : ( n39124 ) ;
assign n39126 =  ( n879 ) ? ( n39115 ) : ( n39125 ) ;
assign n39127 =  ( n172 ) ? ( n5165 ) : ( VREG_18_1 ) ;
assign n39128 =  ( n170 ) ? ( n5164 ) : ( n39127 ) ;
assign n39129 =  ( n168 ) ? ( n5163 ) : ( n39128 ) ;
assign n39130 =  ( n166 ) ? ( n5162 ) : ( n39129 ) ;
assign n39131 =  ( n162 ) ? ( n5161 ) : ( n39130 ) ;
assign n39132 =  ( n172 ) ? ( n5175 ) : ( VREG_18_1 ) ;
assign n39133 =  ( n170 ) ? ( n5174 ) : ( n39132 ) ;
assign n39134 =  ( n168 ) ? ( n5173 ) : ( n39133 ) ;
assign n39135 =  ( n166 ) ? ( n5172 ) : ( n39134 ) ;
assign n39136 =  ( n162 ) ? ( n5171 ) : ( n39135 ) ;
assign n39137 =  ( n5154 ) ? ( VREG_18_1 ) : ( n39136 ) ;
assign n39138 =  ( n3051 ) ? ( n39137 ) : ( VREG_18_1 ) ;
assign n39139 =  ( n3040 ) ? ( n39131 ) : ( n39138 ) ;
assign n39140 =  ( n192 ) ? ( VREG_18_1 ) : ( VREG_18_1 ) ;
assign n39141 =  ( n157 ) ? ( n39139 ) : ( n39140 ) ;
assign n39142 =  ( n6 ) ? ( n39126 ) : ( n39141 ) ;
assign n39143 =  ( n395 ) ? ( n39142 ) : ( VREG_18_1 ) ;
assign n39144 =  ( n148 ) ? ( n6232 ) : ( VREG_18_10 ) ;
assign n39145 =  ( n146 ) ? ( n6231 ) : ( n39144 ) ;
assign n39146 =  ( n144 ) ? ( n6230 ) : ( n39145 ) ;
assign n39147 =  ( n142 ) ? ( n6229 ) : ( n39146 ) ;
assign n39148 =  ( n10 ) ? ( n6228 ) : ( n39147 ) ;
assign n39149 =  ( n148 ) ? ( n7266 ) : ( VREG_18_10 ) ;
assign n39150 =  ( n146 ) ? ( n7265 ) : ( n39149 ) ;
assign n39151 =  ( n144 ) ? ( n7264 ) : ( n39150 ) ;
assign n39152 =  ( n142 ) ? ( n7263 ) : ( n39151 ) ;
assign n39153 =  ( n10 ) ? ( n7262 ) : ( n39152 ) ;
assign n39154 =  ( n7273 ) ? ( VREG_18_10 ) : ( n39148 ) ;
assign n39155 =  ( n7273 ) ? ( VREG_18_10 ) : ( n39153 ) ;
assign n39156 =  ( n3034 ) ? ( n39155 ) : ( VREG_18_10 ) ;
assign n39157 =  ( n2965 ) ? ( n39154 ) : ( n39156 ) ;
assign n39158 =  ( n1930 ) ? ( n39153 ) : ( n39157 ) ;
assign n39159 =  ( n879 ) ? ( n39148 ) : ( n39158 ) ;
assign n39160 =  ( n172 ) ? ( n7284 ) : ( VREG_18_10 ) ;
assign n39161 =  ( n170 ) ? ( n7283 ) : ( n39160 ) ;
assign n39162 =  ( n168 ) ? ( n7282 ) : ( n39161 ) ;
assign n39163 =  ( n166 ) ? ( n7281 ) : ( n39162 ) ;
assign n39164 =  ( n162 ) ? ( n7280 ) : ( n39163 ) ;
assign n39165 =  ( n172 ) ? ( n7294 ) : ( VREG_18_10 ) ;
assign n39166 =  ( n170 ) ? ( n7293 ) : ( n39165 ) ;
assign n39167 =  ( n168 ) ? ( n7292 ) : ( n39166 ) ;
assign n39168 =  ( n166 ) ? ( n7291 ) : ( n39167 ) ;
assign n39169 =  ( n162 ) ? ( n7290 ) : ( n39168 ) ;
assign n39170 =  ( n7273 ) ? ( VREG_18_10 ) : ( n39169 ) ;
assign n39171 =  ( n3051 ) ? ( n39170 ) : ( VREG_18_10 ) ;
assign n39172 =  ( n3040 ) ? ( n39164 ) : ( n39171 ) ;
assign n39173 =  ( n192 ) ? ( VREG_18_10 ) : ( VREG_18_10 ) ;
assign n39174 =  ( n157 ) ? ( n39172 ) : ( n39173 ) ;
assign n39175 =  ( n6 ) ? ( n39159 ) : ( n39174 ) ;
assign n39176 =  ( n395 ) ? ( n39175 ) : ( VREG_18_10 ) ;
assign n39177 =  ( n148 ) ? ( n8351 ) : ( VREG_18_11 ) ;
assign n39178 =  ( n146 ) ? ( n8350 ) : ( n39177 ) ;
assign n39179 =  ( n144 ) ? ( n8349 ) : ( n39178 ) ;
assign n39180 =  ( n142 ) ? ( n8348 ) : ( n39179 ) ;
assign n39181 =  ( n10 ) ? ( n8347 ) : ( n39180 ) ;
assign n39182 =  ( n148 ) ? ( n9385 ) : ( VREG_18_11 ) ;
assign n39183 =  ( n146 ) ? ( n9384 ) : ( n39182 ) ;
assign n39184 =  ( n144 ) ? ( n9383 ) : ( n39183 ) ;
assign n39185 =  ( n142 ) ? ( n9382 ) : ( n39184 ) ;
assign n39186 =  ( n10 ) ? ( n9381 ) : ( n39185 ) ;
assign n39187 =  ( n9392 ) ? ( VREG_18_11 ) : ( n39181 ) ;
assign n39188 =  ( n9392 ) ? ( VREG_18_11 ) : ( n39186 ) ;
assign n39189 =  ( n3034 ) ? ( n39188 ) : ( VREG_18_11 ) ;
assign n39190 =  ( n2965 ) ? ( n39187 ) : ( n39189 ) ;
assign n39191 =  ( n1930 ) ? ( n39186 ) : ( n39190 ) ;
assign n39192 =  ( n879 ) ? ( n39181 ) : ( n39191 ) ;
assign n39193 =  ( n172 ) ? ( n9403 ) : ( VREG_18_11 ) ;
assign n39194 =  ( n170 ) ? ( n9402 ) : ( n39193 ) ;
assign n39195 =  ( n168 ) ? ( n9401 ) : ( n39194 ) ;
assign n39196 =  ( n166 ) ? ( n9400 ) : ( n39195 ) ;
assign n39197 =  ( n162 ) ? ( n9399 ) : ( n39196 ) ;
assign n39198 =  ( n172 ) ? ( n9413 ) : ( VREG_18_11 ) ;
assign n39199 =  ( n170 ) ? ( n9412 ) : ( n39198 ) ;
assign n39200 =  ( n168 ) ? ( n9411 ) : ( n39199 ) ;
assign n39201 =  ( n166 ) ? ( n9410 ) : ( n39200 ) ;
assign n39202 =  ( n162 ) ? ( n9409 ) : ( n39201 ) ;
assign n39203 =  ( n9392 ) ? ( VREG_18_11 ) : ( n39202 ) ;
assign n39204 =  ( n3051 ) ? ( n39203 ) : ( VREG_18_11 ) ;
assign n39205 =  ( n3040 ) ? ( n39197 ) : ( n39204 ) ;
assign n39206 =  ( n192 ) ? ( VREG_18_11 ) : ( VREG_18_11 ) ;
assign n39207 =  ( n157 ) ? ( n39205 ) : ( n39206 ) ;
assign n39208 =  ( n6 ) ? ( n39192 ) : ( n39207 ) ;
assign n39209 =  ( n395 ) ? ( n39208 ) : ( VREG_18_11 ) ;
assign n39210 =  ( n148 ) ? ( n10470 ) : ( VREG_18_12 ) ;
assign n39211 =  ( n146 ) ? ( n10469 ) : ( n39210 ) ;
assign n39212 =  ( n144 ) ? ( n10468 ) : ( n39211 ) ;
assign n39213 =  ( n142 ) ? ( n10467 ) : ( n39212 ) ;
assign n39214 =  ( n10 ) ? ( n10466 ) : ( n39213 ) ;
assign n39215 =  ( n148 ) ? ( n11504 ) : ( VREG_18_12 ) ;
assign n39216 =  ( n146 ) ? ( n11503 ) : ( n39215 ) ;
assign n39217 =  ( n144 ) ? ( n11502 ) : ( n39216 ) ;
assign n39218 =  ( n142 ) ? ( n11501 ) : ( n39217 ) ;
assign n39219 =  ( n10 ) ? ( n11500 ) : ( n39218 ) ;
assign n39220 =  ( n11511 ) ? ( VREG_18_12 ) : ( n39214 ) ;
assign n39221 =  ( n11511 ) ? ( VREG_18_12 ) : ( n39219 ) ;
assign n39222 =  ( n3034 ) ? ( n39221 ) : ( VREG_18_12 ) ;
assign n39223 =  ( n2965 ) ? ( n39220 ) : ( n39222 ) ;
assign n39224 =  ( n1930 ) ? ( n39219 ) : ( n39223 ) ;
assign n39225 =  ( n879 ) ? ( n39214 ) : ( n39224 ) ;
assign n39226 =  ( n172 ) ? ( n11522 ) : ( VREG_18_12 ) ;
assign n39227 =  ( n170 ) ? ( n11521 ) : ( n39226 ) ;
assign n39228 =  ( n168 ) ? ( n11520 ) : ( n39227 ) ;
assign n39229 =  ( n166 ) ? ( n11519 ) : ( n39228 ) ;
assign n39230 =  ( n162 ) ? ( n11518 ) : ( n39229 ) ;
assign n39231 =  ( n172 ) ? ( n11532 ) : ( VREG_18_12 ) ;
assign n39232 =  ( n170 ) ? ( n11531 ) : ( n39231 ) ;
assign n39233 =  ( n168 ) ? ( n11530 ) : ( n39232 ) ;
assign n39234 =  ( n166 ) ? ( n11529 ) : ( n39233 ) ;
assign n39235 =  ( n162 ) ? ( n11528 ) : ( n39234 ) ;
assign n39236 =  ( n11511 ) ? ( VREG_18_12 ) : ( n39235 ) ;
assign n39237 =  ( n3051 ) ? ( n39236 ) : ( VREG_18_12 ) ;
assign n39238 =  ( n3040 ) ? ( n39230 ) : ( n39237 ) ;
assign n39239 =  ( n192 ) ? ( VREG_18_12 ) : ( VREG_18_12 ) ;
assign n39240 =  ( n157 ) ? ( n39238 ) : ( n39239 ) ;
assign n39241 =  ( n6 ) ? ( n39225 ) : ( n39240 ) ;
assign n39242 =  ( n395 ) ? ( n39241 ) : ( VREG_18_12 ) ;
assign n39243 =  ( n148 ) ? ( n12589 ) : ( VREG_18_13 ) ;
assign n39244 =  ( n146 ) ? ( n12588 ) : ( n39243 ) ;
assign n39245 =  ( n144 ) ? ( n12587 ) : ( n39244 ) ;
assign n39246 =  ( n142 ) ? ( n12586 ) : ( n39245 ) ;
assign n39247 =  ( n10 ) ? ( n12585 ) : ( n39246 ) ;
assign n39248 =  ( n148 ) ? ( n13623 ) : ( VREG_18_13 ) ;
assign n39249 =  ( n146 ) ? ( n13622 ) : ( n39248 ) ;
assign n39250 =  ( n144 ) ? ( n13621 ) : ( n39249 ) ;
assign n39251 =  ( n142 ) ? ( n13620 ) : ( n39250 ) ;
assign n39252 =  ( n10 ) ? ( n13619 ) : ( n39251 ) ;
assign n39253 =  ( n13630 ) ? ( VREG_18_13 ) : ( n39247 ) ;
assign n39254 =  ( n13630 ) ? ( VREG_18_13 ) : ( n39252 ) ;
assign n39255 =  ( n3034 ) ? ( n39254 ) : ( VREG_18_13 ) ;
assign n39256 =  ( n2965 ) ? ( n39253 ) : ( n39255 ) ;
assign n39257 =  ( n1930 ) ? ( n39252 ) : ( n39256 ) ;
assign n39258 =  ( n879 ) ? ( n39247 ) : ( n39257 ) ;
assign n39259 =  ( n172 ) ? ( n13641 ) : ( VREG_18_13 ) ;
assign n39260 =  ( n170 ) ? ( n13640 ) : ( n39259 ) ;
assign n39261 =  ( n168 ) ? ( n13639 ) : ( n39260 ) ;
assign n39262 =  ( n166 ) ? ( n13638 ) : ( n39261 ) ;
assign n39263 =  ( n162 ) ? ( n13637 ) : ( n39262 ) ;
assign n39264 =  ( n172 ) ? ( n13651 ) : ( VREG_18_13 ) ;
assign n39265 =  ( n170 ) ? ( n13650 ) : ( n39264 ) ;
assign n39266 =  ( n168 ) ? ( n13649 ) : ( n39265 ) ;
assign n39267 =  ( n166 ) ? ( n13648 ) : ( n39266 ) ;
assign n39268 =  ( n162 ) ? ( n13647 ) : ( n39267 ) ;
assign n39269 =  ( n13630 ) ? ( VREG_18_13 ) : ( n39268 ) ;
assign n39270 =  ( n3051 ) ? ( n39269 ) : ( VREG_18_13 ) ;
assign n39271 =  ( n3040 ) ? ( n39263 ) : ( n39270 ) ;
assign n39272 =  ( n192 ) ? ( VREG_18_13 ) : ( VREG_18_13 ) ;
assign n39273 =  ( n157 ) ? ( n39271 ) : ( n39272 ) ;
assign n39274 =  ( n6 ) ? ( n39258 ) : ( n39273 ) ;
assign n39275 =  ( n395 ) ? ( n39274 ) : ( VREG_18_13 ) ;
assign n39276 =  ( n148 ) ? ( n14708 ) : ( VREG_18_14 ) ;
assign n39277 =  ( n146 ) ? ( n14707 ) : ( n39276 ) ;
assign n39278 =  ( n144 ) ? ( n14706 ) : ( n39277 ) ;
assign n39279 =  ( n142 ) ? ( n14705 ) : ( n39278 ) ;
assign n39280 =  ( n10 ) ? ( n14704 ) : ( n39279 ) ;
assign n39281 =  ( n148 ) ? ( n15742 ) : ( VREG_18_14 ) ;
assign n39282 =  ( n146 ) ? ( n15741 ) : ( n39281 ) ;
assign n39283 =  ( n144 ) ? ( n15740 ) : ( n39282 ) ;
assign n39284 =  ( n142 ) ? ( n15739 ) : ( n39283 ) ;
assign n39285 =  ( n10 ) ? ( n15738 ) : ( n39284 ) ;
assign n39286 =  ( n15749 ) ? ( VREG_18_14 ) : ( n39280 ) ;
assign n39287 =  ( n15749 ) ? ( VREG_18_14 ) : ( n39285 ) ;
assign n39288 =  ( n3034 ) ? ( n39287 ) : ( VREG_18_14 ) ;
assign n39289 =  ( n2965 ) ? ( n39286 ) : ( n39288 ) ;
assign n39290 =  ( n1930 ) ? ( n39285 ) : ( n39289 ) ;
assign n39291 =  ( n879 ) ? ( n39280 ) : ( n39290 ) ;
assign n39292 =  ( n172 ) ? ( n15760 ) : ( VREG_18_14 ) ;
assign n39293 =  ( n170 ) ? ( n15759 ) : ( n39292 ) ;
assign n39294 =  ( n168 ) ? ( n15758 ) : ( n39293 ) ;
assign n39295 =  ( n166 ) ? ( n15757 ) : ( n39294 ) ;
assign n39296 =  ( n162 ) ? ( n15756 ) : ( n39295 ) ;
assign n39297 =  ( n172 ) ? ( n15770 ) : ( VREG_18_14 ) ;
assign n39298 =  ( n170 ) ? ( n15769 ) : ( n39297 ) ;
assign n39299 =  ( n168 ) ? ( n15768 ) : ( n39298 ) ;
assign n39300 =  ( n166 ) ? ( n15767 ) : ( n39299 ) ;
assign n39301 =  ( n162 ) ? ( n15766 ) : ( n39300 ) ;
assign n39302 =  ( n15749 ) ? ( VREG_18_14 ) : ( n39301 ) ;
assign n39303 =  ( n3051 ) ? ( n39302 ) : ( VREG_18_14 ) ;
assign n39304 =  ( n3040 ) ? ( n39296 ) : ( n39303 ) ;
assign n39305 =  ( n192 ) ? ( VREG_18_14 ) : ( VREG_18_14 ) ;
assign n39306 =  ( n157 ) ? ( n39304 ) : ( n39305 ) ;
assign n39307 =  ( n6 ) ? ( n39291 ) : ( n39306 ) ;
assign n39308 =  ( n395 ) ? ( n39307 ) : ( VREG_18_14 ) ;
assign n39309 =  ( n148 ) ? ( n16827 ) : ( VREG_18_15 ) ;
assign n39310 =  ( n146 ) ? ( n16826 ) : ( n39309 ) ;
assign n39311 =  ( n144 ) ? ( n16825 ) : ( n39310 ) ;
assign n39312 =  ( n142 ) ? ( n16824 ) : ( n39311 ) ;
assign n39313 =  ( n10 ) ? ( n16823 ) : ( n39312 ) ;
assign n39314 =  ( n148 ) ? ( n17861 ) : ( VREG_18_15 ) ;
assign n39315 =  ( n146 ) ? ( n17860 ) : ( n39314 ) ;
assign n39316 =  ( n144 ) ? ( n17859 ) : ( n39315 ) ;
assign n39317 =  ( n142 ) ? ( n17858 ) : ( n39316 ) ;
assign n39318 =  ( n10 ) ? ( n17857 ) : ( n39317 ) ;
assign n39319 =  ( n17868 ) ? ( VREG_18_15 ) : ( n39313 ) ;
assign n39320 =  ( n17868 ) ? ( VREG_18_15 ) : ( n39318 ) ;
assign n39321 =  ( n3034 ) ? ( n39320 ) : ( VREG_18_15 ) ;
assign n39322 =  ( n2965 ) ? ( n39319 ) : ( n39321 ) ;
assign n39323 =  ( n1930 ) ? ( n39318 ) : ( n39322 ) ;
assign n39324 =  ( n879 ) ? ( n39313 ) : ( n39323 ) ;
assign n39325 =  ( n172 ) ? ( n17879 ) : ( VREG_18_15 ) ;
assign n39326 =  ( n170 ) ? ( n17878 ) : ( n39325 ) ;
assign n39327 =  ( n168 ) ? ( n17877 ) : ( n39326 ) ;
assign n39328 =  ( n166 ) ? ( n17876 ) : ( n39327 ) ;
assign n39329 =  ( n162 ) ? ( n17875 ) : ( n39328 ) ;
assign n39330 =  ( n172 ) ? ( n17889 ) : ( VREG_18_15 ) ;
assign n39331 =  ( n170 ) ? ( n17888 ) : ( n39330 ) ;
assign n39332 =  ( n168 ) ? ( n17887 ) : ( n39331 ) ;
assign n39333 =  ( n166 ) ? ( n17886 ) : ( n39332 ) ;
assign n39334 =  ( n162 ) ? ( n17885 ) : ( n39333 ) ;
assign n39335 =  ( n17868 ) ? ( VREG_18_15 ) : ( n39334 ) ;
assign n39336 =  ( n3051 ) ? ( n39335 ) : ( VREG_18_15 ) ;
assign n39337 =  ( n3040 ) ? ( n39329 ) : ( n39336 ) ;
assign n39338 =  ( n192 ) ? ( VREG_18_15 ) : ( VREG_18_15 ) ;
assign n39339 =  ( n157 ) ? ( n39337 ) : ( n39338 ) ;
assign n39340 =  ( n6 ) ? ( n39324 ) : ( n39339 ) ;
assign n39341 =  ( n395 ) ? ( n39340 ) : ( VREG_18_15 ) ;
assign n39342 =  ( n148 ) ? ( n18946 ) : ( VREG_18_2 ) ;
assign n39343 =  ( n146 ) ? ( n18945 ) : ( n39342 ) ;
assign n39344 =  ( n144 ) ? ( n18944 ) : ( n39343 ) ;
assign n39345 =  ( n142 ) ? ( n18943 ) : ( n39344 ) ;
assign n39346 =  ( n10 ) ? ( n18942 ) : ( n39345 ) ;
assign n39347 =  ( n148 ) ? ( n19980 ) : ( VREG_18_2 ) ;
assign n39348 =  ( n146 ) ? ( n19979 ) : ( n39347 ) ;
assign n39349 =  ( n144 ) ? ( n19978 ) : ( n39348 ) ;
assign n39350 =  ( n142 ) ? ( n19977 ) : ( n39349 ) ;
assign n39351 =  ( n10 ) ? ( n19976 ) : ( n39350 ) ;
assign n39352 =  ( n19987 ) ? ( VREG_18_2 ) : ( n39346 ) ;
assign n39353 =  ( n19987 ) ? ( VREG_18_2 ) : ( n39351 ) ;
assign n39354 =  ( n3034 ) ? ( n39353 ) : ( VREG_18_2 ) ;
assign n39355 =  ( n2965 ) ? ( n39352 ) : ( n39354 ) ;
assign n39356 =  ( n1930 ) ? ( n39351 ) : ( n39355 ) ;
assign n39357 =  ( n879 ) ? ( n39346 ) : ( n39356 ) ;
assign n39358 =  ( n172 ) ? ( n19998 ) : ( VREG_18_2 ) ;
assign n39359 =  ( n170 ) ? ( n19997 ) : ( n39358 ) ;
assign n39360 =  ( n168 ) ? ( n19996 ) : ( n39359 ) ;
assign n39361 =  ( n166 ) ? ( n19995 ) : ( n39360 ) ;
assign n39362 =  ( n162 ) ? ( n19994 ) : ( n39361 ) ;
assign n39363 =  ( n172 ) ? ( n20008 ) : ( VREG_18_2 ) ;
assign n39364 =  ( n170 ) ? ( n20007 ) : ( n39363 ) ;
assign n39365 =  ( n168 ) ? ( n20006 ) : ( n39364 ) ;
assign n39366 =  ( n166 ) ? ( n20005 ) : ( n39365 ) ;
assign n39367 =  ( n162 ) ? ( n20004 ) : ( n39366 ) ;
assign n39368 =  ( n19987 ) ? ( VREG_18_2 ) : ( n39367 ) ;
assign n39369 =  ( n3051 ) ? ( n39368 ) : ( VREG_18_2 ) ;
assign n39370 =  ( n3040 ) ? ( n39362 ) : ( n39369 ) ;
assign n39371 =  ( n192 ) ? ( VREG_18_2 ) : ( VREG_18_2 ) ;
assign n39372 =  ( n157 ) ? ( n39370 ) : ( n39371 ) ;
assign n39373 =  ( n6 ) ? ( n39357 ) : ( n39372 ) ;
assign n39374 =  ( n395 ) ? ( n39373 ) : ( VREG_18_2 ) ;
assign n39375 =  ( n148 ) ? ( n21065 ) : ( VREG_18_3 ) ;
assign n39376 =  ( n146 ) ? ( n21064 ) : ( n39375 ) ;
assign n39377 =  ( n144 ) ? ( n21063 ) : ( n39376 ) ;
assign n39378 =  ( n142 ) ? ( n21062 ) : ( n39377 ) ;
assign n39379 =  ( n10 ) ? ( n21061 ) : ( n39378 ) ;
assign n39380 =  ( n148 ) ? ( n22099 ) : ( VREG_18_3 ) ;
assign n39381 =  ( n146 ) ? ( n22098 ) : ( n39380 ) ;
assign n39382 =  ( n144 ) ? ( n22097 ) : ( n39381 ) ;
assign n39383 =  ( n142 ) ? ( n22096 ) : ( n39382 ) ;
assign n39384 =  ( n10 ) ? ( n22095 ) : ( n39383 ) ;
assign n39385 =  ( n22106 ) ? ( VREG_18_3 ) : ( n39379 ) ;
assign n39386 =  ( n22106 ) ? ( VREG_18_3 ) : ( n39384 ) ;
assign n39387 =  ( n3034 ) ? ( n39386 ) : ( VREG_18_3 ) ;
assign n39388 =  ( n2965 ) ? ( n39385 ) : ( n39387 ) ;
assign n39389 =  ( n1930 ) ? ( n39384 ) : ( n39388 ) ;
assign n39390 =  ( n879 ) ? ( n39379 ) : ( n39389 ) ;
assign n39391 =  ( n172 ) ? ( n22117 ) : ( VREG_18_3 ) ;
assign n39392 =  ( n170 ) ? ( n22116 ) : ( n39391 ) ;
assign n39393 =  ( n168 ) ? ( n22115 ) : ( n39392 ) ;
assign n39394 =  ( n166 ) ? ( n22114 ) : ( n39393 ) ;
assign n39395 =  ( n162 ) ? ( n22113 ) : ( n39394 ) ;
assign n39396 =  ( n172 ) ? ( n22127 ) : ( VREG_18_3 ) ;
assign n39397 =  ( n170 ) ? ( n22126 ) : ( n39396 ) ;
assign n39398 =  ( n168 ) ? ( n22125 ) : ( n39397 ) ;
assign n39399 =  ( n166 ) ? ( n22124 ) : ( n39398 ) ;
assign n39400 =  ( n162 ) ? ( n22123 ) : ( n39399 ) ;
assign n39401 =  ( n22106 ) ? ( VREG_18_3 ) : ( n39400 ) ;
assign n39402 =  ( n3051 ) ? ( n39401 ) : ( VREG_18_3 ) ;
assign n39403 =  ( n3040 ) ? ( n39395 ) : ( n39402 ) ;
assign n39404 =  ( n192 ) ? ( VREG_18_3 ) : ( VREG_18_3 ) ;
assign n39405 =  ( n157 ) ? ( n39403 ) : ( n39404 ) ;
assign n39406 =  ( n6 ) ? ( n39390 ) : ( n39405 ) ;
assign n39407 =  ( n395 ) ? ( n39406 ) : ( VREG_18_3 ) ;
assign n39408 =  ( n148 ) ? ( n23184 ) : ( VREG_18_4 ) ;
assign n39409 =  ( n146 ) ? ( n23183 ) : ( n39408 ) ;
assign n39410 =  ( n144 ) ? ( n23182 ) : ( n39409 ) ;
assign n39411 =  ( n142 ) ? ( n23181 ) : ( n39410 ) ;
assign n39412 =  ( n10 ) ? ( n23180 ) : ( n39411 ) ;
assign n39413 =  ( n148 ) ? ( n24218 ) : ( VREG_18_4 ) ;
assign n39414 =  ( n146 ) ? ( n24217 ) : ( n39413 ) ;
assign n39415 =  ( n144 ) ? ( n24216 ) : ( n39414 ) ;
assign n39416 =  ( n142 ) ? ( n24215 ) : ( n39415 ) ;
assign n39417 =  ( n10 ) ? ( n24214 ) : ( n39416 ) ;
assign n39418 =  ( n24225 ) ? ( VREG_18_4 ) : ( n39412 ) ;
assign n39419 =  ( n24225 ) ? ( VREG_18_4 ) : ( n39417 ) ;
assign n39420 =  ( n3034 ) ? ( n39419 ) : ( VREG_18_4 ) ;
assign n39421 =  ( n2965 ) ? ( n39418 ) : ( n39420 ) ;
assign n39422 =  ( n1930 ) ? ( n39417 ) : ( n39421 ) ;
assign n39423 =  ( n879 ) ? ( n39412 ) : ( n39422 ) ;
assign n39424 =  ( n172 ) ? ( n24236 ) : ( VREG_18_4 ) ;
assign n39425 =  ( n170 ) ? ( n24235 ) : ( n39424 ) ;
assign n39426 =  ( n168 ) ? ( n24234 ) : ( n39425 ) ;
assign n39427 =  ( n166 ) ? ( n24233 ) : ( n39426 ) ;
assign n39428 =  ( n162 ) ? ( n24232 ) : ( n39427 ) ;
assign n39429 =  ( n172 ) ? ( n24246 ) : ( VREG_18_4 ) ;
assign n39430 =  ( n170 ) ? ( n24245 ) : ( n39429 ) ;
assign n39431 =  ( n168 ) ? ( n24244 ) : ( n39430 ) ;
assign n39432 =  ( n166 ) ? ( n24243 ) : ( n39431 ) ;
assign n39433 =  ( n162 ) ? ( n24242 ) : ( n39432 ) ;
assign n39434 =  ( n24225 ) ? ( VREG_18_4 ) : ( n39433 ) ;
assign n39435 =  ( n3051 ) ? ( n39434 ) : ( VREG_18_4 ) ;
assign n39436 =  ( n3040 ) ? ( n39428 ) : ( n39435 ) ;
assign n39437 =  ( n192 ) ? ( VREG_18_4 ) : ( VREG_18_4 ) ;
assign n39438 =  ( n157 ) ? ( n39436 ) : ( n39437 ) ;
assign n39439 =  ( n6 ) ? ( n39423 ) : ( n39438 ) ;
assign n39440 =  ( n395 ) ? ( n39439 ) : ( VREG_18_4 ) ;
assign n39441 =  ( n148 ) ? ( n25303 ) : ( VREG_18_5 ) ;
assign n39442 =  ( n146 ) ? ( n25302 ) : ( n39441 ) ;
assign n39443 =  ( n144 ) ? ( n25301 ) : ( n39442 ) ;
assign n39444 =  ( n142 ) ? ( n25300 ) : ( n39443 ) ;
assign n39445 =  ( n10 ) ? ( n25299 ) : ( n39444 ) ;
assign n39446 =  ( n148 ) ? ( n26337 ) : ( VREG_18_5 ) ;
assign n39447 =  ( n146 ) ? ( n26336 ) : ( n39446 ) ;
assign n39448 =  ( n144 ) ? ( n26335 ) : ( n39447 ) ;
assign n39449 =  ( n142 ) ? ( n26334 ) : ( n39448 ) ;
assign n39450 =  ( n10 ) ? ( n26333 ) : ( n39449 ) ;
assign n39451 =  ( n26344 ) ? ( VREG_18_5 ) : ( n39445 ) ;
assign n39452 =  ( n26344 ) ? ( VREG_18_5 ) : ( n39450 ) ;
assign n39453 =  ( n3034 ) ? ( n39452 ) : ( VREG_18_5 ) ;
assign n39454 =  ( n2965 ) ? ( n39451 ) : ( n39453 ) ;
assign n39455 =  ( n1930 ) ? ( n39450 ) : ( n39454 ) ;
assign n39456 =  ( n879 ) ? ( n39445 ) : ( n39455 ) ;
assign n39457 =  ( n172 ) ? ( n26355 ) : ( VREG_18_5 ) ;
assign n39458 =  ( n170 ) ? ( n26354 ) : ( n39457 ) ;
assign n39459 =  ( n168 ) ? ( n26353 ) : ( n39458 ) ;
assign n39460 =  ( n166 ) ? ( n26352 ) : ( n39459 ) ;
assign n39461 =  ( n162 ) ? ( n26351 ) : ( n39460 ) ;
assign n39462 =  ( n172 ) ? ( n26365 ) : ( VREG_18_5 ) ;
assign n39463 =  ( n170 ) ? ( n26364 ) : ( n39462 ) ;
assign n39464 =  ( n168 ) ? ( n26363 ) : ( n39463 ) ;
assign n39465 =  ( n166 ) ? ( n26362 ) : ( n39464 ) ;
assign n39466 =  ( n162 ) ? ( n26361 ) : ( n39465 ) ;
assign n39467 =  ( n26344 ) ? ( VREG_18_5 ) : ( n39466 ) ;
assign n39468 =  ( n3051 ) ? ( n39467 ) : ( VREG_18_5 ) ;
assign n39469 =  ( n3040 ) ? ( n39461 ) : ( n39468 ) ;
assign n39470 =  ( n192 ) ? ( VREG_18_5 ) : ( VREG_18_5 ) ;
assign n39471 =  ( n157 ) ? ( n39469 ) : ( n39470 ) ;
assign n39472 =  ( n6 ) ? ( n39456 ) : ( n39471 ) ;
assign n39473 =  ( n395 ) ? ( n39472 ) : ( VREG_18_5 ) ;
assign n39474 =  ( n148 ) ? ( n27422 ) : ( VREG_18_6 ) ;
assign n39475 =  ( n146 ) ? ( n27421 ) : ( n39474 ) ;
assign n39476 =  ( n144 ) ? ( n27420 ) : ( n39475 ) ;
assign n39477 =  ( n142 ) ? ( n27419 ) : ( n39476 ) ;
assign n39478 =  ( n10 ) ? ( n27418 ) : ( n39477 ) ;
assign n39479 =  ( n148 ) ? ( n28456 ) : ( VREG_18_6 ) ;
assign n39480 =  ( n146 ) ? ( n28455 ) : ( n39479 ) ;
assign n39481 =  ( n144 ) ? ( n28454 ) : ( n39480 ) ;
assign n39482 =  ( n142 ) ? ( n28453 ) : ( n39481 ) ;
assign n39483 =  ( n10 ) ? ( n28452 ) : ( n39482 ) ;
assign n39484 =  ( n28463 ) ? ( VREG_18_6 ) : ( n39478 ) ;
assign n39485 =  ( n28463 ) ? ( VREG_18_6 ) : ( n39483 ) ;
assign n39486 =  ( n3034 ) ? ( n39485 ) : ( VREG_18_6 ) ;
assign n39487 =  ( n2965 ) ? ( n39484 ) : ( n39486 ) ;
assign n39488 =  ( n1930 ) ? ( n39483 ) : ( n39487 ) ;
assign n39489 =  ( n879 ) ? ( n39478 ) : ( n39488 ) ;
assign n39490 =  ( n172 ) ? ( n28474 ) : ( VREG_18_6 ) ;
assign n39491 =  ( n170 ) ? ( n28473 ) : ( n39490 ) ;
assign n39492 =  ( n168 ) ? ( n28472 ) : ( n39491 ) ;
assign n39493 =  ( n166 ) ? ( n28471 ) : ( n39492 ) ;
assign n39494 =  ( n162 ) ? ( n28470 ) : ( n39493 ) ;
assign n39495 =  ( n172 ) ? ( n28484 ) : ( VREG_18_6 ) ;
assign n39496 =  ( n170 ) ? ( n28483 ) : ( n39495 ) ;
assign n39497 =  ( n168 ) ? ( n28482 ) : ( n39496 ) ;
assign n39498 =  ( n166 ) ? ( n28481 ) : ( n39497 ) ;
assign n39499 =  ( n162 ) ? ( n28480 ) : ( n39498 ) ;
assign n39500 =  ( n28463 ) ? ( VREG_18_6 ) : ( n39499 ) ;
assign n39501 =  ( n3051 ) ? ( n39500 ) : ( VREG_18_6 ) ;
assign n39502 =  ( n3040 ) ? ( n39494 ) : ( n39501 ) ;
assign n39503 =  ( n192 ) ? ( VREG_18_6 ) : ( VREG_18_6 ) ;
assign n39504 =  ( n157 ) ? ( n39502 ) : ( n39503 ) ;
assign n39505 =  ( n6 ) ? ( n39489 ) : ( n39504 ) ;
assign n39506 =  ( n395 ) ? ( n39505 ) : ( VREG_18_6 ) ;
assign n39507 =  ( n148 ) ? ( n29541 ) : ( VREG_18_7 ) ;
assign n39508 =  ( n146 ) ? ( n29540 ) : ( n39507 ) ;
assign n39509 =  ( n144 ) ? ( n29539 ) : ( n39508 ) ;
assign n39510 =  ( n142 ) ? ( n29538 ) : ( n39509 ) ;
assign n39511 =  ( n10 ) ? ( n29537 ) : ( n39510 ) ;
assign n39512 =  ( n148 ) ? ( n30575 ) : ( VREG_18_7 ) ;
assign n39513 =  ( n146 ) ? ( n30574 ) : ( n39512 ) ;
assign n39514 =  ( n144 ) ? ( n30573 ) : ( n39513 ) ;
assign n39515 =  ( n142 ) ? ( n30572 ) : ( n39514 ) ;
assign n39516 =  ( n10 ) ? ( n30571 ) : ( n39515 ) ;
assign n39517 =  ( n30582 ) ? ( VREG_18_7 ) : ( n39511 ) ;
assign n39518 =  ( n30582 ) ? ( VREG_18_7 ) : ( n39516 ) ;
assign n39519 =  ( n3034 ) ? ( n39518 ) : ( VREG_18_7 ) ;
assign n39520 =  ( n2965 ) ? ( n39517 ) : ( n39519 ) ;
assign n39521 =  ( n1930 ) ? ( n39516 ) : ( n39520 ) ;
assign n39522 =  ( n879 ) ? ( n39511 ) : ( n39521 ) ;
assign n39523 =  ( n172 ) ? ( n30593 ) : ( VREG_18_7 ) ;
assign n39524 =  ( n170 ) ? ( n30592 ) : ( n39523 ) ;
assign n39525 =  ( n168 ) ? ( n30591 ) : ( n39524 ) ;
assign n39526 =  ( n166 ) ? ( n30590 ) : ( n39525 ) ;
assign n39527 =  ( n162 ) ? ( n30589 ) : ( n39526 ) ;
assign n39528 =  ( n172 ) ? ( n30603 ) : ( VREG_18_7 ) ;
assign n39529 =  ( n170 ) ? ( n30602 ) : ( n39528 ) ;
assign n39530 =  ( n168 ) ? ( n30601 ) : ( n39529 ) ;
assign n39531 =  ( n166 ) ? ( n30600 ) : ( n39530 ) ;
assign n39532 =  ( n162 ) ? ( n30599 ) : ( n39531 ) ;
assign n39533 =  ( n30582 ) ? ( VREG_18_7 ) : ( n39532 ) ;
assign n39534 =  ( n3051 ) ? ( n39533 ) : ( VREG_18_7 ) ;
assign n39535 =  ( n3040 ) ? ( n39527 ) : ( n39534 ) ;
assign n39536 =  ( n192 ) ? ( VREG_18_7 ) : ( VREG_18_7 ) ;
assign n39537 =  ( n157 ) ? ( n39535 ) : ( n39536 ) ;
assign n39538 =  ( n6 ) ? ( n39522 ) : ( n39537 ) ;
assign n39539 =  ( n395 ) ? ( n39538 ) : ( VREG_18_7 ) ;
assign n39540 =  ( n148 ) ? ( n31660 ) : ( VREG_18_8 ) ;
assign n39541 =  ( n146 ) ? ( n31659 ) : ( n39540 ) ;
assign n39542 =  ( n144 ) ? ( n31658 ) : ( n39541 ) ;
assign n39543 =  ( n142 ) ? ( n31657 ) : ( n39542 ) ;
assign n39544 =  ( n10 ) ? ( n31656 ) : ( n39543 ) ;
assign n39545 =  ( n148 ) ? ( n32694 ) : ( VREG_18_8 ) ;
assign n39546 =  ( n146 ) ? ( n32693 ) : ( n39545 ) ;
assign n39547 =  ( n144 ) ? ( n32692 ) : ( n39546 ) ;
assign n39548 =  ( n142 ) ? ( n32691 ) : ( n39547 ) ;
assign n39549 =  ( n10 ) ? ( n32690 ) : ( n39548 ) ;
assign n39550 =  ( n32701 ) ? ( VREG_18_8 ) : ( n39544 ) ;
assign n39551 =  ( n32701 ) ? ( VREG_18_8 ) : ( n39549 ) ;
assign n39552 =  ( n3034 ) ? ( n39551 ) : ( VREG_18_8 ) ;
assign n39553 =  ( n2965 ) ? ( n39550 ) : ( n39552 ) ;
assign n39554 =  ( n1930 ) ? ( n39549 ) : ( n39553 ) ;
assign n39555 =  ( n879 ) ? ( n39544 ) : ( n39554 ) ;
assign n39556 =  ( n172 ) ? ( n32712 ) : ( VREG_18_8 ) ;
assign n39557 =  ( n170 ) ? ( n32711 ) : ( n39556 ) ;
assign n39558 =  ( n168 ) ? ( n32710 ) : ( n39557 ) ;
assign n39559 =  ( n166 ) ? ( n32709 ) : ( n39558 ) ;
assign n39560 =  ( n162 ) ? ( n32708 ) : ( n39559 ) ;
assign n39561 =  ( n172 ) ? ( n32722 ) : ( VREG_18_8 ) ;
assign n39562 =  ( n170 ) ? ( n32721 ) : ( n39561 ) ;
assign n39563 =  ( n168 ) ? ( n32720 ) : ( n39562 ) ;
assign n39564 =  ( n166 ) ? ( n32719 ) : ( n39563 ) ;
assign n39565 =  ( n162 ) ? ( n32718 ) : ( n39564 ) ;
assign n39566 =  ( n32701 ) ? ( VREG_18_8 ) : ( n39565 ) ;
assign n39567 =  ( n3051 ) ? ( n39566 ) : ( VREG_18_8 ) ;
assign n39568 =  ( n3040 ) ? ( n39560 ) : ( n39567 ) ;
assign n39569 =  ( n192 ) ? ( VREG_18_8 ) : ( VREG_18_8 ) ;
assign n39570 =  ( n157 ) ? ( n39568 ) : ( n39569 ) ;
assign n39571 =  ( n6 ) ? ( n39555 ) : ( n39570 ) ;
assign n39572 =  ( n395 ) ? ( n39571 ) : ( VREG_18_8 ) ;
assign n39573 =  ( n148 ) ? ( n33779 ) : ( VREG_18_9 ) ;
assign n39574 =  ( n146 ) ? ( n33778 ) : ( n39573 ) ;
assign n39575 =  ( n144 ) ? ( n33777 ) : ( n39574 ) ;
assign n39576 =  ( n142 ) ? ( n33776 ) : ( n39575 ) ;
assign n39577 =  ( n10 ) ? ( n33775 ) : ( n39576 ) ;
assign n39578 =  ( n148 ) ? ( n34813 ) : ( VREG_18_9 ) ;
assign n39579 =  ( n146 ) ? ( n34812 ) : ( n39578 ) ;
assign n39580 =  ( n144 ) ? ( n34811 ) : ( n39579 ) ;
assign n39581 =  ( n142 ) ? ( n34810 ) : ( n39580 ) ;
assign n39582 =  ( n10 ) ? ( n34809 ) : ( n39581 ) ;
assign n39583 =  ( n34820 ) ? ( VREG_18_9 ) : ( n39577 ) ;
assign n39584 =  ( n34820 ) ? ( VREG_18_9 ) : ( n39582 ) ;
assign n39585 =  ( n3034 ) ? ( n39584 ) : ( VREG_18_9 ) ;
assign n39586 =  ( n2965 ) ? ( n39583 ) : ( n39585 ) ;
assign n39587 =  ( n1930 ) ? ( n39582 ) : ( n39586 ) ;
assign n39588 =  ( n879 ) ? ( n39577 ) : ( n39587 ) ;
assign n39589 =  ( n172 ) ? ( n34831 ) : ( VREG_18_9 ) ;
assign n39590 =  ( n170 ) ? ( n34830 ) : ( n39589 ) ;
assign n39591 =  ( n168 ) ? ( n34829 ) : ( n39590 ) ;
assign n39592 =  ( n166 ) ? ( n34828 ) : ( n39591 ) ;
assign n39593 =  ( n162 ) ? ( n34827 ) : ( n39592 ) ;
assign n39594 =  ( n172 ) ? ( n34841 ) : ( VREG_18_9 ) ;
assign n39595 =  ( n170 ) ? ( n34840 ) : ( n39594 ) ;
assign n39596 =  ( n168 ) ? ( n34839 ) : ( n39595 ) ;
assign n39597 =  ( n166 ) ? ( n34838 ) : ( n39596 ) ;
assign n39598 =  ( n162 ) ? ( n34837 ) : ( n39597 ) ;
assign n39599 =  ( n34820 ) ? ( VREG_18_9 ) : ( n39598 ) ;
assign n39600 =  ( n3051 ) ? ( n39599 ) : ( VREG_18_9 ) ;
assign n39601 =  ( n3040 ) ? ( n39593 ) : ( n39600 ) ;
assign n39602 =  ( n192 ) ? ( VREG_18_9 ) : ( VREG_18_9 ) ;
assign n39603 =  ( n157 ) ? ( n39601 ) : ( n39602 ) ;
assign n39604 =  ( n6 ) ? ( n39588 ) : ( n39603 ) ;
assign n39605 =  ( n395 ) ? ( n39604 ) : ( VREG_18_9 ) ;
assign n39606 =  ( n148 ) ? ( n1924 ) : ( VREG_19_0 ) ;
assign n39607 =  ( n146 ) ? ( n1923 ) : ( n39606 ) ;
assign n39608 =  ( n144 ) ? ( n1922 ) : ( n39607 ) ;
assign n39609 =  ( n142 ) ? ( n1921 ) : ( n39608 ) ;
assign n39610 =  ( n10 ) ? ( n1920 ) : ( n39609 ) ;
assign n39611 =  ( n148 ) ? ( n2959 ) : ( VREG_19_0 ) ;
assign n39612 =  ( n146 ) ? ( n2958 ) : ( n39611 ) ;
assign n39613 =  ( n144 ) ? ( n2957 ) : ( n39612 ) ;
assign n39614 =  ( n142 ) ? ( n2956 ) : ( n39613 ) ;
assign n39615 =  ( n10 ) ? ( n2955 ) : ( n39614 ) ;
assign n39616 =  ( n3032 ) ? ( VREG_19_0 ) : ( n39610 ) ;
assign n39617 =  ( n3032 ) ? ( VREG_19_0 ) : ( n39615 ) ;
assign n39618 =  ( n3034 ) ? ( n39617 ) : ( VREG_19_0 ) ;
assign n39619 =  ( n2965 ) ? ( n39616 ) : ( n39618 ) ;
assign n39620 =  ( n1930 ) ? ( n39615 ) : ( n39619 ) ;
assign n39621 =  ( n879 ) ? ( n39610 ) : ( n39620 ) ;
assign n39622 =  ( n172 ) ? ( n3045 ) : ( VREG_19_0 ) ;
assign n39623 =  ( n170 ) ? ( n3044 ) : ( n39622 ) ;
assign n39624 =  ( n168 ) ? ( n3043 ) : ( n39623 ) ;
assign n39625 =  ( n166 ) ? ( n3042 ) : ( n39624 ) ;
assign n39626 =  ( n162 ) ? ( n3041 ) : ( n39625 ) ;
assign n39627 =  ( n172 ) ? ( n3056 ) : ( VREG_19_0 ) ;
assign n39628 =  ( n170 ) ? ( n3055 ) : ( n39627 ) ;
assign n39629 =  ( n168 ) ? ( n3054 ) : ( n39628 ) ;
assign n39630 =  ( n166 ) ? ( n3053 ) : ( n39629 ) ;
assign n39631 =  ( n162 ) ? ( n3052 ) : ( n39630 ) ;
assign n39632 =  ( n3032 ) ? ( VREG_19_0 ) : ( n39631 ) ;
assign n39633 =  ( n3051 ) ? ( n39632 ) : ( VREG_19_0 ) ;
assign n39634 =  ( n3040 ) ? ( n39626 ) : ( n39633 ) ;
assign n39635 =  ( n192 ) ? ( VREG_19_0 ) : ( VREG_19_0 ) ;
assign n39636 =  ( n157 ) ? ( n39634 ) : ( n39635 ) ;
assign n39637 =  ( n6 ) ? ( n39621 ) : ( n39636 ) ;
assign n39638 =  ( n417 ) ? ( n39637 ) : ( VREG_19_0 ) ;
assign n39639 =  ( n148 ) ? ( n4113 ) : ( VREG_19_1 ) ;
assign n39640 =  ( n146 ) ? ( n4112 ) : ( n39639 ) ;
assign n39641 =  ( n144 ) ? ( n4111 ) : ( n39640 ) ;
assign n39642 =  ( n142 ) ? ( n4110 ) : ( n39641 ) ;
assign n39643 =  ( n10 ) ? ( n4109 ) : ( n39642 ) ;
assign n39644 =  ( n148 ) ? ( n5147 ) : ( VREG_19_1 ) ;
assign n39645 =  ( n146 ) ? ( n5146 ) : ( n39644 ) ;
assign n39646 =  ( n144 ) ? ( n5145 ) : ( n39645 ) ;
assign n39647 =  ( n142 ) ? ( n5144 ) : ( n39646 ) ;
assign n39648 =  ( n10 ) ? ( n5143 ) : ( n39647 ) ;
assign n39649 =  ( n5154 ) ? ( VREG_19_1 ) : ( n39643 ) ;
assign n39650 =  ( n5154 ) ? ( VREG_19_1 ) : ( n39648 ) ;
assign n39651 =  ( n3034 ) ? ( n39650 ) : ( VREG_19_1 ) ;
assign n39652 =  ( n2965 ) ? ( n39649 ) : ( n39651 ) ;
assign n39653 =  ( n1930 ) ? ( n39648 ) : ( n39652 ) ;
assign n39654 =  ( n879 ) ? ( n39643 ) : ( n39653 ) ;
assign n39655 =  ( n172 ) ? ( n5165 ) : ( VREG_19_1 ) ;
assign n39656 =  ( n170 ) ? ( n5164 ) : ( n39655 ) ;
assign n39657 =  ( n168 ) ? ( n5163 ) : ( n39656 ) ;
assign n39658 =  ( n166 ) ? ( n5162 ) : ( n39657 ) ;
assign n39659 =  ( n162 ) ? ( n5161 ) : ( n39658 ) ;
assign n39660 =  ( n172 ) ? ( n5175 ) : ( VREG_19_1 ) ;
assign n39661 =  ( n170 ) ? ( n5174 ) : ( n39660 ) ;
assign n39662 =  ( n168 ) ? ( n5173 ) : ( n39661 ) ;
assign n39663 =  ( n166 ) ? ( n5172 ) : ( n39662 ) ;
assign n39664 =  ( n162 ) ? ( n5171 ) : ( n39663 ) ;
assign n39665 =  ( n5154 ) ? ( VREG_19_1 ) : ( n39664 ) ;
assign n39666 =  ( n3051 ) ? ( n39665 ) : ( VREG_19_1 ) ;
assign n39667 =  ( n3040 ) ? ( n39659 ) : ( n39666 ) ;
assign n39668 =  ( n192 ) ? ( VREG_19_1 ) : ( VREG_19_1 ) ;
assign n39669 =  ( n157 ) ? ( n39667 ) : ( n39668 ) ;
assign n39670 =  ( n6 ) ? ( n39654 ) : ( n39669 ) ;
assign n39671 =  ( n417 ) ? ( n39670 ) : ( VREG_19_1 ) ;
assign n39672 =  ( n148 ) ? ( n6232 ) : ( VREG_19_10 ) ;
assign n39673 =  ( n146 ) ? ( n6231 ) : ( n39672 ) ;
assign n39674 =  ( n144 ) ? ( n6230 ) : ( n39673 ) ;
assign n39675 =  ( n142 ) ? ( n6229 ) : ( n39674 ) ;
assign n39676 =  ( n10 ) ? ( n6228 ) : ( n39675 ) ;
assign n39677 =  ( n148 ) ? ( n7266 ) : ( VREG_19_10 ) ;
assign n39678 =  ( n146 ) ? ( n7265 ) : ( n39677 ) ;
assign n39679 =  ( n144 ) ? ( n7264 ) : ( n39678 ) ;
assign n39680 =  ( n142 ) ? ( n7263 ) : ( n39679 ) ;
assign n39681 =  ( n10 ) ? ( n7262 ) : ( n39680 ) ;
assign n39682 =  ( n7273 ) ? ( VREG_19_10 ) : ( n39676 ) ;
assign n39683 =  ( n7273 ) ? ( VREG_19_10 ) : ( n39681 ) ;
assign n39684 =  ( n3034 ) ? ( n39683 ) : ( VREG_19_10 ) ;
assign n39685 =  ( n2965 ) ? ( n39682 ) : ( n39684 ) ;
assign n39686 =  ( n1930 ) ? ( n39681 ) : ( n39685 ) ;
assign n39687 =  ( n879 ) ? ( n39676 ) : ( n39686 ) ;
assign n39688 =  ( n172 ) ? ( n7284 ) : ( VREG_19_10 ) ;
assign n39689 =  ( n170 ) ? ( n7283 ) : ( n39688 ) ;
assign n39690 =  ( n168 ) ? ( n7282 ) : ( n39689 ) ;
assign n39691 =  ( n166 ) ? ( n7281 ) : ( n39690 ) ;
assign n39692 =  ( n162 ) ? ( n7280 ) : ( n39691 ) ;
assign n39693 =  ( n172 ) ? ( n7294 ) : ( VREG_19_10 ) ;
assign n39694 =  ( n170 ) ? ( n7293 ) : ( n39693 ) ;
assign n39695 =  ( n168 ) ? ( n7292 ) : ( n39694 ) ;
assign n39696 =  ( n166 ) ? ( n7291 ) : ( n39695 ) ;
assign n39697 =  ( n162 ) ? ( n7290 ) : ( n39696 ) ;
assign n39698 =  ( n7273 ) ? ( VREG_19_10 ) : ( n39697 ) ;
assign n39699 =  ( n3051 ) ? ( n39698 ) : ( VREG_19_10 ) ;
assign n39700 =  ( n3040 ) ? ( n39692 ) : ( n39699 ) ;
assign n39701 =  ( n192 ) ? ( VREG_19_10 ) : ( VREG_19_10 ) ;
assign n39702 =  ( n157 ) ? ( n39700 ) : ( n39701 ) ;
assign n39703 =  ( n6 ) ? ( n39687 ) : ( n39702 ) ;
assign n39704 =  ( n417 ) ? ( n39703 ) : ( VREG_19_10 ) ;
assign n39705 =  ( n148 ) ? ( n8351 ) : ( VREG_19_11 ) ;
assign n39706 =  ( n146 ) ? ( n8350 ) : ( n39705 ) ;
assign n39707 =  ( n144 ) ? ( n8349 ) : ( n39706 ) ;
assign n39708 =  ( n142 ) ? ( n8348 ) : ( n39707 ) ;
assign n39709 =  ( n10 ) ? ( n8347 ) : ( n39708 ) ;
assign n39710 =  ( n148 ) ? ( n9385 ) : ( VREG_19_11 ) ;
assign n39711 =  ( n146 ) ? ( n9384 ) : ( n39710 ) ;
assign n39712 =  ( n144 ) ? ( n9383 ) : ( n39711 ) ;
assign n39713 =  ( n142 ) ? ( n9382 ) : ( n39712 ) ;
assign n39714 =  ( n10 ) ? ( n9381 ) : ( n39713 ) ;
assign n39715 =  ( n9392 ) ? ( VREG_19_11 ) : ( n39709 ) ;
assign n39716 =  ( n9392 ) ? ( VREG_19_11 ) : ( n39714 ) ;
assign n39717 =  ( n3034 ) ? ( n39716 ) : ( VREG_19_11 ) ;
assign n39718 =  ( n2965 ) ? ( n39715 ) : ( n39717 ) ;
assign n39719 =  ( n1930 ) ? ( n39714 ) : ( n39718 ) ;
assign n39720 =  ( n879 ) ? ( n39709 ) : ( n39719 ) ;
assign n39721 =  ( n172 ) ? ( n9403 ) : ( VREG_19_11 ) ;
assign n39722 =  ( n170 ) ? ( n9402 ) : ( n39721 ) ;
assign n39723 =  ( n168 ) ? ( n9401 ) : ( n39722 ) ;
assign n39724 =  ( n166 ) ? ( n9400 ) : ( n39723 ) ;
assign n39725 =  ( n162 ) ? ( n9399 ) : ( n39724 ) ;
assign n39726 =  ( n172 ) ? ( n9413 ) : ( VREG_19_11 ) ;
assign n39727 =  ( n170 ) ? ( n9412 ) : ( n39726 ) ;
assign n39728 =  ( n168 ) ? ( n9411 ) : ( n39727 ) ;
assign n39729 =  ( n166 ) ? ( n9410 ) : ( n39728 ) ;
assign n39730 =  ( n162 ) ? ( n9409 ) : ( n39729 ) ;
assign n39731 =  ( n9392 ) ? ( VREG_19_11 ) : ( n39730 ) ;
assign n39732 =  ( n3051 ) ? ( n39731 ) : ( VREG_19_11 ) ;
assign n39733 =  ( n3040 ) ? ( n39725 ) : ( n39732 ) ;
assign n39734 =  ( n192 ) ? ( VREG_19_11 ) : ( VREG_19_11 ) ;
assign n39735 =  ( n157 ) ? ( n39733 ) : ( n39734 ) ;
assign n39736 =  ( n6 ) ? ( n39720 ) : ( n39735 ) ;
assign n39737 =  ( n417 ) ? ( n39736 ) : ( VREG_19_11 ) ;
assign n39738 =  ( n148 ) ? ( n10470 ) : ( VREG_19_12 ) ;
assign n39739 =  ( n146 ) ? ( n10469 ) : ( n39738 ) ;
assign n39740 =  ( n144 ) ? ( n10468 ) : ( n39739 ) ;
assign n39741 =  ( n142 ) ? ( n10467 ) : ( n39740 ) ;
assign n39742 =  ( n10 ) ? ( n10466 ) : ( n39741 ) ;
assign n39743 =  ( n148 ) ? ( n11504 ) : ( VREG_19_12 ) ;
assign n39744 =  ( n146 ) ? ( n11503 ) : ( n39743 ) ;
assign n39745 =  ( n144 ) ? ( n11502 ) : ( n39744 ) ;
assign n39746 =  ( n142 ) ? ( n11501 ) : ( n39745 ) ;
assign n39747 =  ( n10 ) ? ( n11500 ) : ( n39746 ) ;
assign n39748 =  ( n11511 ) ? ( VREG_19_12 ) : ( n39742 ) ;
assign n39749 =  ( n11511 ) ? ( VREG_19_12 ) : ( n39747 ) ;
assign n39750 =  ( n3034 ) ? ( n39749 ) : ( VREG_19_12 ) ;
assign n39751 =  ( n2965 ) ? ( n39748 ) : ( n39750 ) ;
assign n39752 =  ( n1930 ) ? ( n39747 ) : ( n39751 ) ;
assign n39753 =  ( n879 ) ? ( n39742 ) : ( n39752 ) ;
assign n39754 =  ( n172 ) ? ( n11522 ) : ( VREG_19_12 ) ;
assign n39755 =  ( n170 ) ? ( n11521 ) : ( n39754 ) ;
assign n39756 =  ( n168 ) ? ( n11520 ) : ( n39755 ) ;
assign n39757 =  ( n166 ) ? ( n11519 ) : ( n39756 ) ;
assign n39758 =  ( n162 ) ? ( n11518 ) : ( n39757 ) ;
assign n39759 =  ( n172 ) ? ( n11532 ) : ( VREG_19_12 ) ;
assign n39760 =  ( n170 ) ? ( n11531 ) : ( n39759 ) ;
assign n39761 =  ( n168 ) ? ( n11530 ) : ( n39760 ) ;
assign n39762 =  ( n166 ) ? ( n11529 ) : ( n39761 ) ;
assign n39763 =  ( n162 ) ? ( n11528 ) : ( n39762 ) ;
assign n39764 =  ( n11511 ) ? ( VREG_19_12 ) : ( n39763 ) ;
assign n39765 =  ( n3051 ) ? ( n39764 ) : ( VREG_19_12 ) ;
assign n39766 =  ( n3040 ) ? ( n39758 ) : ( n39765 ) ;
assign n39767 =  ( n192 ) ? ( VREG_19_12 ) : ( VREG_19_12 ) ;
assign n39768 =  ( n157 ) ? ( n39766 ) : ( n39767 ) ;
assign n39769 =  ( n6 ) ? ( n39753 ) : ( n39768 ) ;
assign n39770 =  ( n417 ) ? ( n39769 ) : ( VREG_19_12 ) ;
assign n39771 =  ( n148 ) ? ( n12589 ) : ( VREG_19_13 ) ;
assign n39772 =  ( n146 ) ? ( n12588 ) : ( n39771 ) ;
assign n39773 =  ( n144 ) ? ( n12587 ) : ( n39772 ) ;
assign n39774 =  ( n142 ) ? ( n12586 ) : ( n39773 ) ;
assign n39775 =  ( n10 ) ? ( n12585 ) : ( n39774 ) ;
assign n39776 =  ( n148 ) ? ( n13623 ) : ( VREG_19_13 ) ;
assign n39777 =  ( n146 ) ? ( n13622 ) : ( n39776 ) ;
assign n39778 =  ( n144 ) ? ( n13621 ) : ( n39777 ) ;
assign n39779 =  ( n142 ) ? ( n13620 ) : ( n39778 ) ;
assign n39780 =  ( n10 ) ? ( n13619 ) : ( n39779 ) ;
assign n39781 =  ( n13630 ) ? ( VREG_19_13 ) : ( n39775 ) ;
assign n39782 =  ( n13630 ) ? ( VREG_19_13 ) : ( n39780 ) ;
assign n39783 =  ( n3034 ) ? ( n39782 ) : ( VREG_19_13 ) ;
assign n39784 =  ( n2965 ) ? ( n39781 ) : ( n39783 ) ;
assign n39785 =  ( n1930 ) ? ( n39780 ) : ( n39784 ) ;
assign n39786 =  ( n879 ) ? ( n39775 ) : ( n39785 ) ;
assign n39787 =  ( n172 ) ? ( n13641 ) : ( VREG_19_13 ) ;
assign n39788 =  ( n170 ) ? ( n13640 ) : ( n39787 ) ;
assign n39789 =  ( n168 ) ? ( n13639 ) : ( n39788 ) ;
assign n39790 =  ( n166 ) ? ( n13638 ) : ( n39789 ) ;
assign n39791 =  ( n162 ) ? ( n13637 ) : ( n39790 ) ;
assign n39792 =  ( n172 ) ? ( n13651 ) : ( VREG_19_13 ) ;
assign n39793 =  ( n170 ) ? ( n13650 ) : ( n39792 ) ;
assign n39794 =  ( n168 ) ? ( n13649 ) : ( n39793 ) ;
assign n39795 =  ( n166 ) ? ( n13648 ) : ( n39794 ) ;
assign n39796 =  ( n162 ) ? ( n13647 ) : ( n39795 ) ;
assign n39797 =  ( n13630 ) ? ( VREG_19_13 ) : ( n39796 ) ;
assign n39798 =  ( n3051 ) ? ( n39797 ) : ( VREG_19_13 ) ;
assign n39799 =  ( n3040 ) ? ( n39791 ) : ( n39798 ) ;
assign n39800 =  ( n192 ) ? ( VREG_19_13 ) : ( VREG_19_13 ) ;
assign n39801 =  ( n157 ) ? ( n39799 ) : ( n39800 ) ;
assign n39802 =  ( n6 ) ? ( n39786 ) : ( n39801 ) ;
assign n39803 =  ( n417 ) ? ( n39802 ) : ( VREG_19_13 ) ;
assign n39804 =  ( n148 ) ? ( n14708 ) : ( VREG_19_14 ) ;
assign n39805 =  ( n146 ) ? ( n14707 ) : ( n39804 ) ;
assign n39806 =  ( n144 ) ? ( n14706 ) : ( n39805 ) ;
assign n39807 =  ( n142 ) ? ( n14705 ) : ( n39806 ) ;
assign n39808 =  ( n10 ) ? ( n14704 ) : ( n39807 ) ;
assign n39809 =  ( n148 ) ? ( n15742 ) : ( VREG_19_14 ) ;
assign n39810 =  ( n146 ) ? ( n15741 ) : ( n39809 ) ;
assign n39811 =  ( n144 ) ? ( n15740 ) : ( n39810 ) ;
assign n39812 =  ( n142 ) ? ( n15739 ) : ( n39811 ) ;
assign n39813 =  ( n10 ) ? ( n15738 ) : ( n39812 ) ;
assign n39814 =  ( n15749 ) ? ( VREG_19_14 ) : ( n39808 ) ;
assign n39815 =  ( n15749 ) ? ( VREG_19_14 ) : ( n39813 ) ;
assign n39816 =  ( n3034 ) ? ( n39815 ) : ( VREG_19_14 ) ;
assign n39817 =  ( n2965 ) ? ( n39814 ) : ( n39816 ) ;
assign n39818 =  ( n1930 ) ? ( n39813 ) : ( n39817 ) ;
assign n39819 =  ( n879 ) ? ( n39808 ) : ( n39818 ) ;
assign n39820 =  ( n172 ) ? ( n15760 ) : ( VREG_19_14 ) ;
assign n39821 =  ( n170 ) ? ( n15759 ) : ( n39820 ) ;
assign n39822 =  ( n168 ) ? ( n15758 ) : ( n39821 ) ;
assign n39823 =  ( n166 ) ? ( n15757 ) : ( n39822 ) ;
assign n39824 =  ( n162 ) ? ( n15756 ) : ( n39823 ) ;
assign n39825 =  ( n172 ) ? ( n15770 ) : ( VREG_19_14 ) ;
assign n39826 =  ( n170 ) ? ( n15769 ) : ( n39825 ) ;
assign n39827 =  ( n168 ) ? ( n15768 ) : ( n39826 ) ;
assign n39828 =  ( n166 ) ? ( n15767 ) : ( n39827 ) ;
assign n39829 =  ( n162 ) ? ( n15766 ) : ( n39828 ) ;
assign n39830 =  ( n15749 ) ? ( VREG_19_14 ) : ( n39829 ) ;
assign n39831 =  ( n3051 ) ? ( n39830 ) : ( VREG_19_14 ) ;
assign n39832 =  ( n3040 ) ? ( n39824 ) : ( n39831 ) ;
assign n39833 =  ( n192 ) ? ( VREG_19_14 ) : ( VREG_19_14 ) ;
assign n39834 =  ( n157 ) ? ( n39832 ) : ( n39833 ) ;
assign n39835 =  ( n6 ) ? ( n39819 ) : ( n39834 ) ;
assign n39836 =  ( n417 ) ? ( n39835 ) : ( VREG_19_14 ) ;
assign n39837 =  ( n148 ) ? ( n16827 ) : ( VREG_19_15 ) ;
assign n39838 =  ( n146 ) ? ( n16826 ) : ( n39837 ) ;
assign n39839 =  ( n144 ) ? ( n16825 ) : ( n39838 ) ;
assign n39840 =  ( n142 ) ? ( n16824 ) : ( n39839 ) ;
assign n39841 =  ( n10 ) ? ( n16823 ) : ( n39840 ) ;
assign n39842 =  ( n148 ) ? ( n17861 ) : ( VREG_19_15 ) ;
assign n39843 =  ( n146 ) ? ( n17860 ) : ( n39842 ) ;
assign n39844 =  ( n144 ) ? ( n17859 ) : ( n39843 ) ;
assign n39845 =  ( n142 ) ? ( n17858 ) : ( n39844 ) ;
assign n39846 =  ( n10 ) ? ( n17857 ) : ( n39845 ) ;
assign n39847 =  ( n17868 ) ? ( VREG_19_15 ) : ( n39841 ) ;
assign n39848 =  ( n17868 ) ? ( VREG_19_15 ) : ( n39846 ) ;
assign n39849 =  ( n3034 ) ? ( n39848 ) : ( VREG_19_15 ) ;
assign n39850 =  ( n2965 ) ? ( n39847 ) : ( n39849 ) ;
assign n39851 =  ( n1930 ) ? ( n39846 ) : ( n39850 ) ;
assign n39852 =  ( n879 ) ? ( n39841 ) : ( n39851 ) ;
assign n39853 =  ( n172 ) ? ( n17879 ) : ( VREG_19_15 ) ;
assign n39854 =  ( n170 ) ? ( n17878 ) : ( n39853 ) ;
assign n39855 =  ( n168 ) ? ( n17877 ) : ( n39854 ) ;
assign n39856 =  ( n166 ) ? ( n17876 ) : ( n39855 ) ;
assign n39857 =  ( n162 ) ? ( n17875 ) : ( n39856 ) ;
assign n39858 =  ( n172 ) ? ( n17889 ) : ( VREG_19_15 ) ;
assign n39859 =  ( n170 ) ? ( n17888 ) : ( n39858 ) ;
assign n39860 =  ( n168 ) ? ( n17887 ) : ( n39859 ) ;
assign n39861 =  ( n166 ) ? ( n17886 ) : ( n39860 ) ;
assign n39862 =  ( n162 ) ? ( n17885 ) : ( n39861 ) ;
assign n39863 =  ( n17868 ) ? ( VREG_19_15 ) : ( n39862 ) ;
assign n39864 =  ( n3051 ) ? ( n39863 ) : ( VREG_19_15 ) ;
assign n39865 =  ( n3040 ) ? ( n39857 ) : ( n39864 ) ;
assign n39866 =  ( n192 ) ? ( VREG_19_15 ) : ( VREG_19_15 ) ;
assign n39867 =  ( n157 ) ? ( n39865 ) : ( n39866 ) ;
assign n39868 =  ( n6 ) ? ( n39852 ) : ( n39867 ) ;
assign n39869 =  ( n417 ) ? ( n39868 ) : ( VREG_19_15 ) ;
assign n39870 =  ( n148 ) ? ( n18946 ) : ( VREG_19_2 ) ;
assign n39871 =  ( n146 ) ? ( n18945 ) : ( n39870 ) ;
assign n39872 =  ( n144 ) ? ( n18944 ) : ( n39871 ) ;
assign n39873 =  ( n142 ) ? ( n18943 ) : ( n39872 ) ;
assign n39874 =  ( n10 ) ? ( n18942 ) : ( n39873 ) ;
assign n39875 =  ( n148 ) ? ( n19980 ) : ( VREG_19_2 ) ;
assign n39876 =  ( n146 ) ? ( n19979 ) : ( n39875 ) ;
assign n39877 =  ( n144 ) ? ( n19978 ) : ( n39876 ) ;
assign n39878 =  ( n142 ) ? ( n19977 ) : ( n39877 ) ;
assign n39879 =  ( n10 ) ? ( n19976 ) : ( n39878 ) ;
assign n39880 =  ( n19987 ) ? ( VREG_19_2 ) : ( n39874 ) ;
assign n39881 =  ( n19987 ) ? ( VREG_19_2 ) : ( n39879 ) ;
assign n39882 =  ( n3034 ) ? ( n39881 ) : ( VREG_19_2 ) ;
assign n39883 =  ( n2965 ) ? ( n39880 ) : ( n39882 ) ;
assign n39884 =  ( n1930 ) ? ( n39879 ) : ( n39883 ) ;
assign n39885 =  ( n879 ) ? ( n39874 ) : ( n39884 ) ;
assign n39886 =  ( n172 ) ? ( n19998 ) : ( VREG_19_2 ) ;
assign n39887 =  ( n170 ) ? ( n19997 ) : ( n39886 ) ;
assign n39888 =  ( n168 ) ? ( n19996 ) : ( n39887 ) ;
assign n39889 =  ( n166 ) ? ( n19995 ) : ( n39888 ) ;
assign n39890 =  ( n162 ) ? ( n19994 ) : ( n39889 ) ;
assign n39891 =  ( n172 ) ? ( n20008 ) : ( VREG_19_2 ) ;
assign n39892 =  ( n170 ) ? ( n20007 ) : ( n39891 ) ;
assign n39893 =  ( n168 ) ? ( n20006 ) : ( n39892 ) ;
assign n39894 =  ( n166 ) ? ( n20005 ) : ( n39893 ) ;
assign n39895 =  ( n162 ) ? ( n20004 ) : ( n39894 ) ;
assign n39896 =  ( n19987 ) ? ( VREG_19_2 ) : ( n39895 ) ;
assign n39897 =  ( n3051 ) ? ( n39896 ) : ( VREG_19_2 ) ;
assign n39898 =  ( n3040 ) ? ( n39890 ) : ( n39897 ) ;
assign n39899 =  ( n192 ) ? ( VREG_19_2 ) : ( VREG_19_2 ) ;
assign n39900 =  ( n157 ) ? ( n39898 ) : ( n39899 ) ;
assign n39901 =  ( n6 ) ? ( n39885 ) : ( n39900 ) ;
assign n39902 =  ( n417 ) ? ( n39901 ) : ( VREG_19_2 ) ;
assign n39903 =  ( n148 ) ? ( n21065 ) : ( VREG_19_3 ) ;
assign n39904 =  ( n146 ) ? ( n21064 ) : ( n39903 ) ;
assign n39905 =  ( n144 ) ? ( n21063 ) : ( n39904 ) ;
assign n39906 =  ( n142 ) ? ( n21062 ) : ( n39905 ) ;
assign n39907 =  ( n10 ) ? ( n21061 ) : ( n39906 ) ;
assign n39908 =  ( n148 ) ? ( n22099 ) : ( VREG_19_3 ) ;
assign n39909 =  ( n146 ) ? ( n22098 ) : ( n39908 ) ;
assign n39910 =  ( n144 ) ? ( n22097 ) : ( n39909 ) ;
assign n39911 =  ( n142 ) ? ( n22096 ) : ( n39910 ) ;
assign n39912 =  ( n10 ) ? ( n22095 ) : ( n39911 ) ;
assign n39913 =  ( n22106 ) ? ( VREG_19_3 ) : ( n39907 ) ;
assign n39914 =  ( n22106 ) ? ( VREG_19_3 ) : ( n39912 ) ;
assign n39915 =  ( n3034 ) ? ( n39914 ) : ( VREG_19_3 ) ;
assign n39916 =  ( n2965 ) ? ( n39913 ) : ( n39915 ) ;
assign n39917 =  ( n1930 ) ? ( n39912 ) : ( n39916 ) ;
assign n39918 =  ( n879 ) ? ( n39907 ) : ( n39917 ) ;
assign n39919 =  ( n172 ) ? ( n22117 ) : ( VREG_19_3 ) ;
assign n39920 =  ( n170 ) ? ( n22116 ) : ( n39919 ) ;
assign n39921 =  ( n168 ) ? ( n22115 ) : ( n39920 ) ;
assign n39922 =  ( n166 ) ? ( n22114 ) : ( n39921 ) ;
assign n39923 =  ( n162 ) ? ( n22113 ) : ( n39922 ) ;
assign n39924 =  ( n172 ) ? ( n22127 ) : ( VREG_19_3 ) ;
assign n39925 =  ( n170 ) ? ( n22126 ) : ( n39924 ) ;
assign n39926 =  ( n168 ) ? ( n22125 ) : ( n39925 ) ;
assign n39927 =  ( n166 ) ? ( n22124 ) : ( n39926 ) ;
assign n39928 =  ( n162 ) ? ( n22123 ) : ( n39927 ) ;
assign n39929 =  ( n22106 ) ? ( VREG_19_3 ) : ( n39928 ) ;
assign n39930 =  ( n3051 ) ? ( n39929 ) : ( VREG_19_3 ) ;
assign n39931 =  ( n3040 ) ? ( n39923 ) : ( n39930 ) ;
assign n39932 =  ( n192 ) ? ( VREG_19_3 ) : ( VREG_19_3 ) ;
assign n39933 =  ( n157 ) ? ( n39931 ) : ( n39932 ) ;
assign n39934 =  ( n6 ) ? ( n39918 ) : ( n39933 ) ;
assign n39935 =  ( n417 ) ? ( n39934 ) : ( VREG_19_3 ) ;
assign n39936 =  ( n148 ) ? ( n23184 ) : ( VREG_19_4 ) ;
assign n39937 =  ( n146 ) ? ( n23183 ) : ( n39936 ) ;
assign n39938 =  ( n144 ) ? ( n23182 ) : ( n39937 ) ;
assign n39939 =  ( n142 ) ? ( n23181 ) : ( n39938 ) ;
assign n39940 =  ( n10 ) ? ( n23180 ) : ( n39939 ) ;
assign n39941 =  ( n148 ) ? ( n24218 ) : ( VREG_19_4 ) ;
assign n39942 =  ( n146 ) ? ( n24217 ) : ( n39941 ) ;
assign n39943 =  ( n144 ) ? ( n24216 ) : ( n39942 ) ;
assign n39944 =  ( n142 ) ? ( n24215 ) : ( n39943 ) ;
assign n39945 =  ( n10 ) ? ( n24214 ) : ( n39944 ) ;
assign n39946 =  ( n24225 ) ? ( VREG_19_4 ) : ( n39940 ) ;
assign n39947 =  ( n24225 ) ? ( VREG_19_4 ) : ( n39945 ) ;
assign n39948 =  ( n3034 ) ? ( n39947 ) : ( VREG_19_4 ) ;
assign n39949 =  ( n2965 ) ? ( n39946 ) : ( n39948 ) ;
assign n39950 =  ( n1930 ) ? ( n39945 ) : ( n39949 ) ;
assign n39951 =  ( n879 ) ? ( n39940 ) : ( n39950 ) ;
assign n39952 =  ( n172 ) ? ( n24236 ) : ( VREG_19_4 ) ;
assign n39953 =  ( n170 ) ? ( n24235 ) : ( n39952 ) ;
assign n39954 =  ( n168 ) ? ( n24234 ) : ( n39953 ) ;
assign n39955 =  ( n166 ) ? ( n24233 ) : ( n39954 ) ;
assign n39956 =  ( n162 ) ? ( n24232 ) : ( n39955 ) ;
assign n39957 =  ( n172 ) ? ( n24246 ) : ( VREG_19_4 ) ;
assign n39958 =  ( n170 ) ? ( n24245 ) : ( n39957 ) ;
assign n39959 =  ( n168 ) ? ( n24244 ) : ( n39958 ) ;
assign n39960 =  ( n166 ) ? ( n24243 ) : ( n39959 ) ;
assign n39961 =  ( n162 ) ? ( n24242 ) : ( n39960 ) ;
assign n39962 =  ( n24225 ) ? ( VREG_19_4 ) : ( n39961 ) ;
assign n39963 =  ( n3051 ) ? ( n39962 ) : ( VREG_19_4 ) ;
assign n39964 =  ( n3040 ) ? ( n39956 ) : ( n39963 ) ;
assign n39965 =  ( n192 ) ? ( VREG_19_4 ) : ( VREG_19_4 ) ;
assign n39966 =  ( n157 ) ? ( n39964 ) : ( n39965 ) ;
assign n39967 =  ( n6 ) ? ( n39951 ) : ( n39966 ) ;
assign n39968 =  ( n417 ) ? ( n39967 ) : ( VREG_19_4 ) ;
assign n39969 =  ( n148 ) ? ( n25303 ) : ( VREG_19_5 ) ;
assign n39970 =  ( n146 ) ? ( n25302 ) : ( n39969 ) ;
assign n39971 =  ( n144 ) ? ( n25301 ) : ( n39970 ) ;
assign n39972 =  ( n142 ) ? ( n25300 ) : ( n39971 ) ;
assign n39973 =  ( n10 ) ? ( n25299 ) : ( n39972 ) ;
assign n39974 =  ( n148 ) ? ( n26337 ) : ( VREG_19_5 ) ;
assign n39975 =  ( n146 ) ? ( n26336 ) : ( n39974 ) ;
assign n39976 =  ( n144 ) ? ( n26335 ) : ( n39975 ) ;
assign n39977 =  ( n142 ) ? ( n26334 ) : ( n39976 ) ;
assign n39978 =  ( n10 ) ? ( n26333 ) : ( n39977 ) ;
assign n39979 =  ( n26344 ) ? ( VREG_19_5 ) : ( n39973 ) ;
assign n39980 =  ( n26344 ) ? ( VREG_19_5 ) : ( n39978 ) ;
assign n39981 =  ( n3034 ) ? ( n39980 ) : ( VREG_19_5 ) ;
assign n39982 =  ( n2965 ) ? ( n39979 ) : ( n39981 ) ;
assign n39983 =  ( n1930 ) ? ( n39978 ) : ( n39982 ) ;
assign n39984 =  ( n879 ) ? ( n39973 ) : ( n39983 ) ;
assign n39985 =  ( n172 ) ? ( n26355 ) : ( VREG_19_5 ) ;
assign n39986 =  ( n170 ) ? ( n26354 ) : ( n39985 ) ;
assign n39987 =  ( n168 ) ? ( n26353 ) : ( n39986 ) ;
assign n39988 =  ( n166 ) ? ( n26352 ) : ( n39987 ) ;
assign n39989 =  ( n162 ) ? ( n26351 ) : ( n39988 ) ;
assign n39990 =  ( n172 ) ? ( n26365 ) : ( VREG_19_5 ) ;
assign n39991 =  ( n170 ) ? ( n26364 ) : ( n39990 ) ;
assign n39992 =  ( n168 ) ? ( n26363 ) : ( n39991 ) ;
assign n39993 =  ( n166 ) ? ( n26362 ) : ( n39992 ) ;
assign n39994 =  ( n162 ) ? ( n26361 ) : ( n39993 ) ;
assign n39995 =  ( n26344 ) ? ( VREG_19_5 ) : ( n39994 ) ;
assign n39996 =  ( n3051 ) ? ( n39995 ) : ( VREG_19_5 ) ;
assign n39997 =  ( n3040 ) ? ( n39989 ) : ( n39996 ) ;
assign n39998 =  ( n192 ) ? ( VREG_19_5 ) : ( VREG_19_5 ) ;
assign n39999 =  ( n157 ) ? ( n39997 ) : ( n39998 ) ;
assign n40000 =  ( n6 ) ? ( n39984 ) : ( n39999 ) ;
assign n40001 =  ( n417 ) ? ( n40000 ) : ( VREG_19_5 ) ;
assign n40002 =  ( n148 ) ? ( n27422 ) : ( VREG_19_6 ) ;
assign n40003 =  ( n146 ) ? ( n27421 ) : ( n40002 ) ;
assign n40004 =  ( n144 ) ? ( n27420 ) : ( n40003 ) ;
assign n40005 =  ( n142 ) ? ( n27419 ) : ( n40004 ) ;
assign n40006 =  ( n10 ) ? ( n27418 ) : ( n40005 ) ;
assign n40007 =  ( n148 ) ? ( n28456 ) : ( VREG_19_6 ) ;
assign n40008 =  ( n146 ) ? ( n28455 ) : ( n40007 ) ;
assign n40009 =  ( n144 ) ? ( n28454 ) : ( n40008 ) ;
assign n40010 =  ( n142 ) ? ( n28453 ) : ( n40009 ) ;
assign n40011 =  ( n10 ) ? ( n28452 ) : ( n40010 ) ;
assign n40012 =  ( n28463 ) ? ( VREG_19_6 ) : ( n40006 ) ;
assign n40013 =  ( n28463 ) ? ( VREG_19_6 ) : ( n40011 ) ;
assign n40014 =  ( n3034 ) ? ( n40013 ) : ( VREG_19_6 ) ;
assign n40015 =  ( n2965 ) ? ( n40012 ) : ( n40014 ) ;
assign n40016 =  ( n1930 ) ? ( n40011 ) : ( n40015 ) ;
assign n40017 =  ( n879 ) ? ( n40006 ) : ( n40016 ) ;
assign n40018 =  ( n172 ) ? ( n28474 ) : ( VREG_19_6 ) ;
assign n40019 =  ( n170 ) ? ( n28473 ) : ( n40018 ) ;
assign n40020 =  ( n168 ) ? ( n28472 ) : ( n40019 ) ;
assign n40021 =  ( n166 ) ? ( n28471 ) : ( n40020 ) ;
assign n40022 =  ( n162 ) ? ( n28470 ) : ( n40021 ) ;
assign n40023 =  ( n172 ) ? ( n28484 ) : ( VREG_19_6 ) ;
assign n40024 =  ( n170 ) ? ( n28483 ) : ( n40023 ) ;
assign n40025 =  ( n168 ) ? ( n28482 ) : ( n40024 ) ;
assign n40026 =  ( n166 ) ? ( n28481 ) : ( n40025 ) ;
assign n40027 =  ( n162 ) ? ( n28480 ) : ( n40026 ) ;
assign n40028 =  ( n28463 ) ? ( VREG_19_6 ) : ( n40027 ) ;
assign n40029 =  ( n3051 ) ? ( n40028 ) : ( VREG_19_6 ) ;
assign n40030 =  ( n3040 ) ? ( n40022 ) : ( n40029 ) ;
assign n40031 =  ( n192 ) ? ( VREG_19_6 ) : ( VREG_19_6 ) ;
assign n40032 =  ( n157 ) ? ( n40030 ) : ( n40031 ) ;
assign n40033 =  ( n6 ) ? ( n40017 ) : ( n40032 ) ;
assign n40034 =  ( n417 ) ? ( n40033 ) : ( VREG_19_6 ) ;
assign n40035 =  ( n148 ) ? ( n29541 ) : ( VREG_19_7 ) ;
assign n40036 =  ( n146 ) ? ( n29540 ) : ( n40035 ) ;
assign n40037 =  ( n144 ) ? ( n29539 ) : ( n40036 ) ;
assign n40038 =  ( n142 ) ? ( n29538 ) : ( n40037 ) ;
assign n40039 =  ( n10 ) ? ( n29537 ) : ( n40038 ) ;
assign n40040 =  ( n148 ) ? ( n30575 ) : ( VREG_19_7 ) ;
assign n40041 =  ( n146 ) ? ( n30574 ) : ( n40040 ) ;
assign n40042 =  ( n144 ) ? ( n30573 ) : ( n40041 ) ;
assign n40043 =  ( n142 ) ? ( n30572 ) : ( n40042 ) ;
assign n40044 =  ( n10 ) ? ( n30571 ) : ( n40043 ) ;
assign n40045 =  ( n30582 ) ? ( VREG_19_7 ) : ( n40039 ) ;
assign n40046 =  ( n30582 ) ? ( VREG_19_7 ) : ( n40044 ) ;
assign n40047 =  ( n3034 ) ? ( n40046 ) : ( VREG_19_7 ) ;
assign n40048 =  ( n2965 ) ? ( n40045 ) : ( n40047 ) ;
assign n40049 =  ( n1930 ) ? ( n40044 ) : ( n40048 ) ;
assign n40050 =  ( n879 ) ? ( n40039 ) : ( n40049 ) ;
assign n40051 =  ( n172 ) ? ( n30593 ) : ( VREG_19_7 ) ;
assign n40052 =  ( n170 ) ? ( n30592 ) : ( n40051 ) ;
assign n40053 =  ( n168 ) ? ( n30591 ) : ( n40052 ) ;
assign n40054 =  ( n166 ) ? ( n30590 ) : ( n40053 ) ;
assign n40055 =  ( n162 ) ? ( n30589 ) : ( n40054 ) ;
assign n40056 =  ( n172 ) ? ( n30603 ) : ( VREG_19_7 ) ;
assign n40057 =  ( n170 ) ? ( n30602 ) : ( n40056 ) ;
assign n40058 =  ( n168 ) ? ( n30601 ) : ( n40057 ) ;
assign n40059 =  ( n166 ) ? ( n30600 ) : ( n40058 ) ;
assign n40060 =  ( n162 ) ? ( n30599 ) : ( n40059 ) ;
assign n40061 =  ( n30582 ) ? ( VREG_19_7 ) : ( n40060 ) ;
assign n40062 =  ( n3051 ) ? ( n40061 ) : ( VREG_19_7 ) ;
assign n40063 =  ( n3040 ) ? ( n40055 ) : ( n40062 ) ;
assign n40064 =  ( n192 ) ? ( VREG_19_7 ) : ( VREG_19_7 ) ;
assign n40065 =  ( n157 ) ? ( n40063 ) : ( n40064 ) ;
assign n40066 =  ( n6 ) ? ( n40050 ) : ( n40065 ) ;
assign n40067 =  ( n417 ) ? ( n40066 ) : ( VREG_19_7 ) ;
assign n40068 =  ( n148 ) ? ( n31660 ) : ( VREG_19_8 ) ;
assign n40069 =  ( n146 ) ? ( n31659 ) : ( n40068 ) ;
assign n40070 =  ( n144 ) ? ( n31658 ) : ( n40069 ) ;
assign n40071 =  ( n142 ) ? ( n31657 ) : ( n40070 ) ;
assign n40072 =  ( n10 ) ? ( n31656 ) : ( n40071 ) ;
assign n40073 =  ( n148 ) ? ( n32694 ) : ( VREG_19_8 ) ;
assign n40074 =  ( n146 ) ? ( n32693 ) : ( n40073 ) ;
assign n40075 =  ( n144 ) ? ( n32692 ) : ( n40074 ) ;
assign n40076 =  ( n142 ) ? ( n32691 ) : ( n40075 ) ;
assign n40077 =  ( n10 ) ? ( n32690 ) : ( n40076 ) ;
assign n40078 =  ( n32701 ) ? ( VREG_19_8 ) : ( n40072 ) ;
assign n40079 =  ( n32701 ) ? ( VREG_19_8 ) : ( n40077 ) ;
assign n40080 =  ( n3034 ) ? ( n40079 ) : ( VREG_19_8 ) ;
assign n40081 =  ( n2965 ) ? ( n40078 ) : ( n40080 ) ;
assign n40082 =  ( n1930 ) ? ( n40077 ) : ( n40081 ) ;
assign n40083 =  ( n879 ) ? ( n40072 ) : ( n40082 ) ;
assign n40084 =  ( n172 ) ? ( n32712 ) : ( VREG_19_8 ) ;
assign n40085 =  ( n170 ) ? ( n32711 ) : ( n40084 ) ;
assign n40086 =  ( n168 ) ? ( n32710 ) : ( n40085 ) ;
assign n40087 =  ( n166 ) ? ( n32709 ) : ( n40086 ) ;
assign n40088 =  ( n162 ) ? ( n32708 ) : ( n40087 ) ;
assign n40089 =  ( n172 ) ? ( n32722 ) : ( VREG_19_8 ) ;
assign n40090 =  ( n170 ) ? ( n32721 ) : ( n40089 ) ;
assign n40091 =  ( n168 ) ? ( n32720 ) : ( n40090 ) ;
assign n40092 =  ( n166 ) ? ( n32719 ) : ( n40091 ) ;
assign n40093 =  ( n162 ) ? ( n32718 ) : ( n40092 ) ;
assign n40094 =  ( n32701 ) ? ( VREG_19_8 ) : ( n40093 ) ;
assign n40095 =  ( n3051 ) ? ( n40094 ) : ( VREG_19_8 ) ;
assign n40096 =  ( n3040 ) ? ( n40088 ) : ( n40095 ) ;
assign n40097 =  ( n192 ) ? ( VREG_19_8 ) : ( VREG_19_8 ) ;
assign n40098 =  ( n157 ) ? ( n40096 ) : ( n40097 ) ;
assign n40099 =  ( n6 ) ? ( n40083 ) : ( n40098 ) ;
assign n40100 =  ( n417 ) ? ( n40099 ) : ( VREG_19_8 ) ;
assign n40101 =  ( n148 ) ? ( n33779 ) : ( VREG_19_9 ) ;
assign n40102 =  ( n146 ) ? ( n33778 ) : ( n40101 ) ;
assign n40103 =  ( n144 ) ? ( n33777 ) : ( n40102 ) ;
assign n40104 =  ( n142 ) ? ( n33776 ) : ( n40103 ) ;
assign n40105 =  ( n10 ) ? ( n33775 ) : ( n40104 ) ;
assign n40106 =  ( n148 ) ? ( n34813 ) : ( VREG_19_9 ) ;
assign n40107 =  ( n146 ) ? ( n34812 ) : ( n40106 ) ;
assign n40108 =  ( n144 ) ? ( n34811 ) : ( n40107 ) ;
assign n40109 =  ( n142 ) ? ( n34810 ) : ( n40108 ) ;
assign n40110 =  ( n10 ) ? ( n34809 ) : ( n40109 ) ;
assign n40111 =  ( n34820 ) ? ( VREG_19_9 ) : ( n40105 ) ;
assign n40112 =  ( n34820 ) ? ( VREG_19_9 ) : ( n40110 ) ;
assign n40113 =  ( n3034 ) ? ( n40112 ) : ( VREG_19_9 ) ;
assign n40114 =  ( n2965 ) ? ( n40111 ) : ( n40113 ) ;
assign n40115 =  ( n1930 ) ? ( n40110 ) : ( n40114 ) ;
assign n40116 =  ( n879 ) ? ( n40105 ) : ( n40115 ) ;
assign n40117 =  ( n172 ) ? ( n34831 ) : ( VREG_19_9 ) ;
assign n40118 =  ( n170 ) ? ( n34830 ) : ( n40117 ) ;
assign n40119 =  ( n168 ) ? ( n34829 ) : ( n40118 ) ;
assign n40120 =  ( n166 ) ? ( n34828 ) : ( n40119 ) ;
assign n40121 =  ( n162 ) ? ( n34827 ) : ( n40120 ) ;
assign n40122 =  ( n172 ) ? ( n34841 ) : ( VREG_19_9 ) ;
assign n40123 =  ( n170 ) ? ( n34840 ) : ( n40122 ) ;
assign n40124 =  ( n168 ) ? ( n34839 ) : ( n40123 ) ;
assign n40125 =  ( n166 ) ? ( n34838 ) : ( n40124 ) ;
assign n40126 =  ( n162 ) ? ( n34837 ) : ( n40125 ) ;
assign n40127 =  ( n34820 ) ? ( VREG_19_9 ) : ( n40126 ) ;
assign n40128 =  ( n3051 ) ? ( n40127 ) : ( VREG_19_9 ) ;
assign n40129 =  ( n3040 ) ? ( n40121 ) : ( n40128 ) ;
assign n40130 =  ( n192 ) ? ( VREG_19_9 ) : ( VREG_19_9 ) ;
assign n40131 =  ( n157 ) ? ( n40129 ) : ( n40130 ) ;
assign n40132 =  ( n6 ) ? ( n40116 ) : ( n40131 ) ;
assign n40133 =  ( n417 ) ? ( n40132 ) : ( VREG_19_9 ) ;
assign n40134 =  ( n148 ) ? ( n1924 ) : ( VREG_1_0 ) ;
assign n40135 =  ( n146 ) ? ( n1923 ) : ( n40134 ) ;
assign n40136 =  ( n144 ) ? ( n1922 ) : ( n40135 ) ;
assign n40137 =  ( n142 ) ? ( n1921 ) : ( n40136 ) ;
assign n40138 =  ( n10 ) ? ( n1920 ) : ( n40137 ) ;
assign n40139 =  ( n148 ) ? ( n2959 ) : ( VREG_1_0 ) ;
assign n40140 =  ( n146 ) ? ( n2958 ) : ( n40139 ) ;
assign n40141 =  ( n144 ) ? ( n2957 ) : ( n40140 ) ;
assign n40142 =  ( n142 ) ? ( n2956 ) : ( n40141 ) ;
assign n40143 =  ( n10 ) ? ( n2955 ) : ( n40142 ) ;
assign n40144 =  ( n3032 ) ? ( VREG_1_0 ) : ( n40138 ) ;
assign n40145 =  ( n3032 ) ? ( VREG_1_0 ) : ( n40143 ) ;
assign n40146 =  ( n3034 ) ? ( n40145 ) : ( VREG_1_0 ) ;
assign n40147 =  ( n2965 ) ? ( n40144 ) : ( n40146 ) ;
assign n40148 =  ( n1930 ) ? ( n40143 ) : ( n40147 ) ;
assign n40149 =  ( n879 ) ? ( n40138 ) : ( n40148 ) ;
assign n40150 =  ( n172 ) ? ( n3045 ) : ( VREG_1_0 ) ;
assign n40151 =  ( n170 ) ? ( n3044 ) : ( n40150 ) ;
assign n40152 =  ( n168 ) ? ( n3043 ) : ( n40151 ) ;
assign n40153 =  ( n166 ) ? ( n3042 ) : ( n40152 ) ;
assign n40154 =  ( n162 ) ? ( n3041 ) : ( n40153 ) ;
assign n40155 =  ( n172 ) ? ( n3056 ) : ( VREG_1_0 ) ;
assign n40156 =  ( n170 ) ? ( n3055 ) : ( n40155 ) ;
assign n40157 =  ( n168 ) ? ( n3054 ) : ( n40156 ) ;
assign n40158 =  ( n166 ) ? ( n3053 ) : ( n40157 ) ;
assign n40159 =  ( n162 ) ? ( n3052 ) : ( n40158 ) ;
assign n40160 =  ( n3032 ) ? ( VREG_1_0 ) : ( n40159 ) ;
assign n40161 =  ( n3051 ) ? ( n40160 ) : ( VREG_1_0 ) ;
assign n40162 =  ( n3040 ) ? ( n40154 ) : ( n40161 ) ;
assign n40163 =  ( n192 ) ? ( VREG_1_0 ) : ( VREG_1_0 ) ;
assign n40164 =  ( n157 ) ? ( n40162 ) : ( n40163 ) ;
assign n40165 =  ( n6 ) ? ( n40149 ) : ( n40164 ) ;
assign n40166 =  ( n197 ) ? ( n40165 ) : ( VREG_1_0 ) ;
assign n40167 =  ( n148 ) ? ( n4113 ) : ( VREG_1_1 ) ;
assign n40168 =  ( n146 ) ? ( n4112 ) : ( n40167 ) ;
assign n40169 =  ( n144 ) ? ( n4111 ) : ( n40168 ) ;
assign n40170 =  ( n142 ) ? ( n4110 ) : ( n40169 ) ;
assign n40171 =  ( n10 ) ? ( n4109 ) : ( n40170 ) ;
assign n40172 =  ( n148 ) ? ( n5147 ) : ( VREG_1_1 ) ;
assign n40173 =  ( n146 ) ? ( n5146 ) : ( n40172 ) ;
assign n40174 =  ( n144 ) ? ( n5145 ) : ( n40173 ) ;
assign n40175 =  ( n142 ) ? ( n5144 ) : ( n40174 ) ;
assign n40176 =  ( n10 ) ? ( n5143 ) : ( n40175 ) ;
assign n40177 =  ( n5154 ) ? ( VREG_1_1 ) : ( n40171 ) ;
assign n40178 =  ( n5154 ) ? ( VREG_1_1 ) : ( n40176 ) ;
assign n40179 =  ( n3034 ) ? ( n40178 ) : ( VREG_1_1 ) ;
assign n40180 =  ( n2965 ) ? ( n40177 ) : ( n40179 ) ;
assign n40181 =  ( n1930 ) ? ( n40176 ) : ( n40180 ) ;
assign n40182 =  ( n879 ) ? ( n40171 ) : ( n40181 ) ;
assign n40183 =  ( n172 ) ? ( n5165 ) : ( VREG_1_1 ) ;
assign n40184 =  ( n170 ) ? ( n5164 ) : ( n40183 ) ;
assign n40185 =  ( n168 ) ? ( n5163 ) : ( n40184 ) ;
assign n40186 =  ( n166 ) ? ( n5162 ) : ( n40185 ) ;
assign n40187 =  ( n162 ) ? ( n5161 ) : ( n40186 ) ;
assign n40188 =  ( n172 ) ? ( n5175 ) : ( VREG_1_1 ) ;
assign n40189 =  ( n170 ) ? ( n5174 ) : ( n40188 ) ;
assign n40190 =  ( n168 ) ? ( n5173 ) : ( n40189 ) ;
assign n40191 =  ( n166 ) ? ( n5172 ) : ( n40190 ) ;
assign n40192 =  ( n162 ) ? ( n5171 ) : ( n40191 ) ;
assign n40193 =  ( n5154 ) ? ( VREG_1_1 ) : ( n40192 ) ;
assign n40194 =  ( n3051 ) ? ( n40193 ) : ( VREG_1_1 ) ;
assign n40195 =  ( n3040 ) ? ( n40187 ) : ( n40194 ) ;
assign n40196 =  ( n192 ) ? ( VREG_1_1 ) : ( VREG_1_1 ) ;
assign n40197 =  ( n157 ) ? ( n40195 ) : ( n40196 ) ;
assign n40198 =  ( n6 ) ? ( n40182 ) : ( n40197 ) ;
assign n40199 =  ( n197 ) ? ( n40198 ) : ( VREG_1_1 ) ;
assign n40200 =  ( n148 ) ? ( n6232 ) : ( VREG_1_10 ) ;
assign n40201 =  ( n146 ) ? ( n6231 ) : ( n40200 ) ;
assign n40202 =  ( n144 ) ? ( n6230 ) : ( n40201 ) ;
assign n40203 =  ( n142 ) ? ( n6229 ) : ( n40202 ) ;
assign n40204 =  ( n10 ) ? ( n6228 ) : ( n40203 ) ;
assign n40205 =  ( n148 ) ? ( n7266 ) : ( VREG_1_10 ) ;
assign n40206 =  ( n146 ) ? ( n7265 ) : ( n40205 ) ;
assign n40207 =  ( n144 ) ? ( n7264 ) : ( n40206 ) ;
assign n40208 =  ( n142 ) ? ( n7263 ) : ( n40207 ) ;
assign n40209 =  ( n10 ) ? ( n7262 ) : ( n40208 ) ;
assign n40210 =  ( n7273 ) ? ( VREG_1_10 ) : ( n40204 ) ;
assign n40211 =  ( n7273 ) ? ( VREG_1_10 ) : ( n40209 ) ;
assign n40212 =  ( n3034 ) ? ( n40211 ) : ( VREG_1_10 ) ;
assign n40213 =  ( n2965 ) ? ( n40210 ) : ( n40212 ) ;
assign n40214 =  ( n1930 ) ? ( n40209 ) : ( n40213 ) ;
assign n40215 =  ( n879 ) ? ( n40204 ) : ( n40214 ) ;
assign n40216 =  ( n172 ) ? ( n7284 ) : ( VREG_1_10 ) ;
assign n40217 =  ( n170 ) ? ( n7283 ) : ( n40216 ) ;
assign n40218 =  ( n168 ) ? ( n7282 ) : ( n40217 ) ;
assign n40219 =  ( n166 ) ? ( n7281 ) : ( n40218 ) ;
assign n40220 =  ( n162 ) ? ( n7280 ) : ( n40219 ) ;
assign n40221 =  ( n172 ) ? ( n7294 ) : ( VREG_1_10 ) ;
assign n40222 =  ( n170 ) ? ( n7293 ) : ( n40221 ) ;
assign n40223 =  ( n168 ) ? ( n7292 ) : ( n40222 ) ;
assign n40224 =  ( n166 ) ? ( n7291 ) : ( n40223 ) ;
assign n40225 =  ( n162 ) ? ( n7290 ) : ( n40224 ) ;
assign n40226 =  ( n7273 ) ? ( VREG_1_10 ) : ( n40225 ) ;
assign n40227 =  ( n3051 ) ? ( n40226 ) : ( VREG_1_10 ) ;
assign n40228 =  ( n3040 ) ? ( n40220 ) : ( n40227 ) ;
assign n40229 =  ( n192 ) ? ( VREG_1_10 ) : ( VREG_1_10 ) ;
assign n40230 =  ( n157 ) ? ( n40228 ) : ( n40229 ) ;
assign n40231 =  ( n6 ) ? ( n40215 ) : ( n40230 ) ;
assign n40232 =  ( n197 ) ? ( n40231 ) : ( VREG_1_10 ) ;
assign n40233 =  ( n148 ) ? ( n8351 ) : ( VREG_1_11 ) ;
assign n40234 =  ( n146 ) ? ( n8350 ) : ( n40233 ) ;
assign n40235 =  ( n144 ) ? ( n8349 ) : ( n40234 ) ;
assign n40236 =  ( n142 ) ? ( n8348 ) : ( n40235 ) ;
assign n40237 =  ( n10 ) ? ( n8347 ) : ( n40236 ) ;
assign n40238 =  ( n148 ) ? ( n9385 ) : ( VREG_1_11 ) ;
assign n40239 =  ( n146 ) ? ( n9384 ) : ( n40238 ) ;
assign n40240 =  ( n144 ) ? ( n9383 ) : ( n40239 ) ;
assign n40241 =  ( n142 ) ? ( n9382 ) : ( n40240 ) ;
assign n40242 =  ( n10 ) ? ( n9381 ) : ( n40241 ) ;
assign n40243 =  ( n9392 ) ? ( VREG_1_11 ) : ( n40237 ) ;
assign n40244 =  ( n9392 ) ? ( VREG_1_11 ) : ( n40242 ) ;
assign n40245 =  ( n3034 ) ? ( n40244 ) : ( VREG_1_11 ) ;
assign n40246 =  ( n2965 ) ? ( n40243 ) : ( n40245 ) ;
assign n40247 =  ( n1930 ) ? ( n40242 ) : ( n40246 ) ;
assign n40248 =  ( n879 ) ? ( n40237 ) : ( n40247 ) ;
assign n40249 =  ( n172 ) ? ( n9403 ) : ( VREG_1_11 ) ;
assign n40250 =  ( n170 ) ? ( n9402 ) : ( n40249 ) ;
assign n40251 =  ( n168 ) ? ( n9401 ) : ( n40250 ) ;
assign n40252 =  ( n166 ) ? ( n9400 ) : ( n40251 ) ;
assign n40253 =  ( n162 ) ? ( n9399 ) : ( n40252 ) ;
assign n40254 =  ( n172 ) ? ( n9413 ) : ( VREG_1_11 ) ;
assign n40255 =  ( n170 ) ? ( n9412 ) : ( n40254 ) ;
assign n40256 =  ( n168 ) ? ( n9411 ) : ( n40255 ) ;
assign n40257 =  ( n166 ) ? ( n9410 ) : ( n40256 ) ;
assign n40258 =  ( n162 ) ? ( n9409 ) : ( n40257 ) ;
assign n40259 =  ( n9392 ) ? ( VREG_1_11 ) : ( n40258 ) ;
assign n40260 =  ( n3051 ) ? ( n40259 ) : ( VREG_1_11 ) ;
assign n40261 =  ( n3040 ) ? ( n40253 ) : ( n40260 ) ;
assign n40262 =  ( n192 ) ? ( VREG_1_11 ) : ( VREG_1_11 ) ;
assign n40263 =  ( n157 ) ? ( n40261 ) : ( n40262 ) ;
assign n40264 =  ( n6 ) ? ( n40248 ) : ( n40263 ) ;
assign n40265 =  ( n197 ) ? ( n40264 ) : ( VREG_1_11 ) ;
assign n40266 =  ( n148 ) ? ( n10470 ) : ( VREG_1_12 ) ;
assign n40267 =  ( n146 ) ? ( n10469 ) : ( n40266 ) ;
assign n40268 =  ( n144 ) ? ( n10468 ) : ( n40267 ) ;
assign n40269 =  ( n142 ) ? ( n10467 ) : ( n40268 ) ;
assign n40270 =  ( n10 ) ? ( n10466 ) : ( n40269 ) ;
assign n40271 =  ( n148 ) ? ( n11504 ) : ( VREG_1_12 ) ;
assign n40272 =  ( n146 ) ? ( n11503 ) : ( n40271 ) ;
assign n40273 =  ( n144 ) ? ( n11502 ) : ( n40272 ) ;
assign n40274 =  ( n142 ) ? ( n11501 ) : ( n40273 ) ;
assign n40275 =  ( n10 ) ? ( n11500 ) : ( n40274 ) ;
assign n40276 =  ( n11511 ) ? ( VREG_1_12 ) : ( n40270 ) ;
assign n40277 =  ( n11511 ) ? ( VREG_1_12 ) : ( n40275 ) ;
assign n40278 =  ( n3034 ) ? ( n40277 ) : ( VREG_1_12 ) ;
assign n40279 =  ( n2965 ) ? ( n40276 ) : ( n40278 ) ;
assign n40280 =  ( n1930 ) ? ( n40275 ) : ( n40279 ) ;
assign n40281 =  ( n879 ) ? ( n40270 ) : ( n40280 ) ;
assign n40282 =  ( n172 ) ? ( n11522 ) : ( VREG_1_12 ) ;
assign n40283 =  ( n170 ) ? ( n11521 ) : ( n40282 ) ;
assign n40284 =  ( n168 ) ? ( n11520 ) : ( n40283 ) ;
assign n40285 =  ( n166 ) ? ( n11519 ) : ( n40284 ) ;
assign n40286 =  ( n162 ) ? ( n11518 ) : ( n40285 ) ;
assign n40287 =  ( n172 ) ? ( n11532 ) : ( VREG_1_12 ) ;
assign n40288 =  ( n170 ) ? ( n11531 ) : ( n40287 ) ;
assign n40289 =  ( n168 ) ? ( n11530 ) : ( n40288 ) ;
assign n40290 =  ( n166 ) ? ( n11529 ) : ( n40289 ) ;
assign n40291 =  ( n162 ) ? ( n11528 ) : ( n40290 ) ;
assign n40292 =  ( n11511 ) ? ( VREG_1_12 ) : ( n40291 ) ;
assign n40293 =  ( n3051 ) ? ( n40292 ) : ( VREG_1_12 ) ;
assign n40294 =  ( n3040 ) ? ( n40286 ) : ( n40293 ) ;
assign n40295 =  ( n192 ) ? ( VREG_1_12 ) : ( VREG_1_12 ) ;
assign n40296 =  ( n157 ) ? ( n40294 ) : ( n40295 ) ;
assign n40297 =  ( n6 ) ? ( n40281 ) : ( n40296 ) ;
assign n40298 =  ( n197 ) ? ( n40297 ) : ( VREG_1_12 ) ;
assign n40299 =  ( n148 ) ? ( n12589 ) : ( VREG_1_13 ) ;
assign n40300 =  ( n146 ) ? ( n12588 ) : ( n40299 ) ;
assign n40301 =  ( n144 ) ? ( n12587 ) : ( n40300 ) ;
assign n40302 =  ( n142 ) ? ( n12586 ) : ( n40301 ) ;
assign n40303 =  ( n10 ) ? ( n12585 ) : ( n40302 ) ;
assign n40304 =  ( n148 ) ? ( n13623 ) : ( VREG_1_13 ) ;
assign n40305 =  ( n146 ) ? ( n13622 ) : ( n40304 ) ;
assign n40306 =  ( n144 ) ? ( n13621 ) : ( n40305 ) ;
assign n40307 =  ( n142 ) ? ( n13620 ) : ( n40306 ) ;
assign n40308 =  ( n10 ) ? ( n13619 ) : ( n40307 ) ;
assign n40309 =  ( n13630 ) ? ( VREG_1_13 ) : ( n40303 ) ;
assign n40310 =  ( n13630 ) ? ( VREG_1_13 ) : ( n40308 ) ;
assign n40311 =  ( n3034 ) ? ( n40310 ) : ( VREG_1_13 ) ;
assign n40312 =  ( n2965 ) ? ( n40309 ) : ( n40311 ) ;
assign n40313 =  ( n1930 ) ? ( n40308 ) : ( n40312 ) ;
assign n40314 =  ( n879 ) ? ( n40303 ) : ( n40313 ) ;
assign n40315 =  ( n172 ) ? ( n13641 ) : ( VREG_1_13 ) ;
assign n40316 =  ( n170 ) ? ( n13640 ) : ( n40315 ) ;
assign n40317 =  ( n168 ) ? ( n13639 ) : ( n40316 ) ;
assign n40318 =  ( n166 ) ? ( n13638 ) : ( n40317 ) ;
assign n40319 =  ( n162 ) ? ( n13637 ) : ( n40318 ) ;
assign n40320 =  ( n172 ) ? ( n13651 ) : ( VREG_1_13 ) ;
assign n40321 =  ( n170 ) ? ( n13650 ) : ( n40320 ) ;
assign n40322 =  ( n168 ) ? ( n13649 ) : ( n40321 ) ;
assign n40323 =  ( n166 ) ? ( n13648 ) : ( n40322 ) ;
assign n40324 =  ( n162 ) ? ( n13647 ) : ( n40323 ) ;
assign n40325 =  ( n13630 ) ? ( VREG_1_13 ) : ( n40324 ) ;
assign n40326 =  ( n3051 ) ? ( n40325 ) : ( VREG_1_13 ) ;
assign n40327 =  ( n3040 ) ? ( n40319 ) : ( n40326 ) ;
assign n40328 =  ( n192 ) ? ( VREG_1_13 ) : ( VREG_1_13 ) ;
assign n40329 =  ( n157 ) ? ( n40327 ) : ( n40328 ) ;
assign n40330 =  ( n6 ) ? ( n40314 ) : ( n40329 ) ;
assign n40331 =  ( n197 ) ? ( n40330 ) : ( VREG_1_13 ) ;
assign n40332 =  ( n148 ) ? ( n14708 ) : ( VREG_1_14 ) ;
assign n40333 =  ( n146 ) ? ( n14707 ) : ( n40332 ) ;
assign n40334 =  ( n144 ) ? ( n14706 ) : ( n40333 ) ;
assign n40335 =  ( n142 ) ? ( n14705 ) : ( n40334 ) ;
assign n40336 =  ( n10 ) ? ( n14704 ) : ( n40335 ) ;
assign n40337 =  ( n148 ) ? ( n15742 ) : ( VREG_1_14 ) ;
assign n40338 =  ( n146 ) ? ( n15741 ) : ( n40337 ) ;
assign n40339 =  ( n144 ) ? ( n15740 ) : ( n40338 ) ;
assign n40340 =  ( n142 ) ? ( n15739 ) : ( n40339 ) ;
assign n40341 =  ( n10 ) ? ( n15738 ) : ( n40340 ) ;
assign n40342 =  ( n15749 ) ? ( VREG_1_14 ) : ( n40336 ) ;
assign n40343 =  ( n15749 ) ? ( VREG_1_14 ) : ( n40341 ) ;
assign n40344 =  ( n3034 ) ? ( n40343 ) : ( VREG_1_14 ) ;
assign n40345 =  ( n2965 ) ? ( n40342 ) : ( n40344 ) ;
assign n40346 =  ( n1930 ) ? ( n40341 ) : ( n40345 ) ;
assign n40347 =  ( n879 ) ? ( n40336 ) : ( n40346 ) ;
assign n40348 =  ( n172 ) ? ( n15760 ) : ( VREG_1_14 ) ;
assign n40349 =  ( n170 ) ? ( n15759 ) : ( n40348 ) ;
assign n40350 =  ( n168 ) ? ( n15758 ) : ( n40349 ) ;
assign n40351 =  ( n166 ) ? ( n15757 ) : ( n40350 ) ;
assign n40352 =  ( n162 ) ? ( n15756 ) : ( n40351 ) ;
assign n40353 =  ( n172 ) ? ( n15770 ) : ( VREG_1_14 ) ;
assign n40354 =  ( n170 ) ? ( n15769 ) : ( n40353 ) ;
assign n40355 =  ( n168 ) ? ( n15768 ) : ( n40354 ) ;
assign n40356 =  ( n166 ) ? ( n15767 ) : ( n40355 ) ;
assign n40357 =  ( n162 ) ? ( n15766 ) : ( n40356 ) ;
assign n40358 =  ( n15749 ) ? ( VREG_1_14 ) : ( n40357 ) ;
assign n40359 =  ( n3051 ) ? ( n40358 ) : ( VREG_1_14 ) ;
assign n40360 =  ( n3040 ) ? ( n40352 ) : ( n40359 ) ;
assign n40361 =  ( n192 ) ? ( VREG_1_14 ) : ( VREG_1_14 ) ;
assign n40362 =  ( n157 ) ? ( n40360 ) : ( n40361 ) ;
assign n40363 =  ( n6 ) ? ( n40347 ) : ( n40362 ) ;
assign n40364 =  ( n197 ) ? ( n40363 ) : ( VREG_1_14 ) ;
assign n40365 =  ( n148 ) ? ( n16827 ) : ( VREG_1_15 ) ;
assign n40366 =  ( n146 ) ? ( n16826 ) : ( n40365 ) ;
assign n40367 =  ( n144 ) ? ( n16825 ) : ( n40366 ) ;
assign n40368 =  ( n142 ) ? ( n16824 ) : ( n40367 ) ;
assign n40369 =  ( n10 ) ? ( n16823 ) : ( n40368 ) ;
assign n40370 =  ( n148 ) ? ( n17861 ) : ( VREG_1_15 ) ;
assign n40371 =  ( n146 ) ? ( n17860 ) : ( n40370 ) ;
assign n40372 =  ( n144 ) ? ( n17859 ) : ( n40371 ) ;
assign n40373 =  ( n142 ) ? ( n17858 ) : ( n40372 ) ;
assign n40374 =  ( n10 ) ? ( n17857 ) : ( n40373 ) ;
assign n40375 =  ( n17868 ) ? ( VREG_1_15 ) : ( n40369 ) ;
assign n40376 =  ( n17868 ) ? ( VREG_1_15 ) : ( n40374 ) ;
assign n40377 =  ( n3034 ) ? ( n40376 ) : ( VREG_1_15 ) ;
assign n40378 =  ( n2965 ) ? ( n40375 ) : ( n40377 ) ;
assign n40379 =  ( n1930 ) ? ( n40374 ) : ( n40378 ) ;
assign n40380 =  ( n879 ) ? ( n40369 ) : ( n40379 ) ;
assign n40381 =  ( n172 ) ? ( n17879 ) : ( VREG_1_15 ) ;
assign n40382 =  ( n170 ) ? ( n17878 ) : ( n40381 ) ;
assign n40383 =  ( n168 ) ? ( n17877 ) : ( n40382 ) ;
assign n40384 =  ( n166 ) ? ( n17876 ) : ( n40383 ) ;
assign n40385 =  ( n162 ) ? ( n17875 ) : ( n40384 ) ;
assign n40386 =  ( n172 ) ? ( n17889 ) : ( VREG_1_15 ) ;
assign n40387 =  ( n170 ) ? ( n17888 ) : ( n40386 ) ;
assign n40388 =  ( n168 ) ? ( n17887 ) : ( n40387 ) ;
assign n40389 =  ( n166 ) ? ( n17886 ) : ( n40388 ) ;
assign n40390 =  ( n162 ) ? ( n17885 ) : ( n40389 ) ;
assign n40391 =  ( n17868 ) ? ( VREG_1_15 ) : ( n40390 ) ;
assign n40392 =  ( n3051 ) ? ( n40391 ) : ( VREG_1_15 ) ;
assign n40393 =  ( n3040 ) ? ( n40385 ) : ( n40392 ) ;
assign n40394 =  ( n192 ) ? ( VREG_1_15 ) : ( VREG_1_15 ) ;
assign n40395 =  ( n157 ) ? ( n40393 ) : ( n40394 ) ;
assign n40396 =  ( n6 ) ? ( n40380 ) : ( n40395 ) ;
assign n40397 =  ( n197 ) ? ( n40396 ) : ( VREG_1_15 ) ;
assign n40398 =  ( n148 ) ? ( n18946 ) : ( VREG_1_2 ) ;
assign n40399 =  ( n146 ) ? ( n18945 ) : ( n40398 ) ;
assign n40400 =  ( n144 ) ? ( n18944 ) : ( n40399 ) ;
assign n40401 =  ( n142 ) ? ( n18943 ) : ( n40400 ) ;
assign n40402 =  ( n10 ) ? ( n18942 ) : ( n40401 ) ;
assign n40403 =  ( n148 ) ? ( n19980 ) : ( VREG_1_2 ) ;
assign n40404 =  ( n146 ) ? ( n19979 ) : ( n40403 ) ;
assign n40405 =  ( n144 ) ? ( n19978 ) : ( n40404 ) ;
assign n40406 =  ( n142 ) ? ( n19977 ) : ( n40405 ) ;
assign n40407 =  ( n10 ) ? ( n19976 ) : ( n40406 ) ;
assign n40408 =  ( n19987 ) ? ( VREG_1_2 ) : ( n40402 ) ;
assign n40409 =  ( n19987 ) ? ( VREG_1_2 ) : ( n40407 ) ;
assign n40410 =  ( n3034 ) ? ( n40409 ) : ( VREG_1_2 ) ;
assign n40411 =  ( n2965 ) ? ( n40408 ) : ( n40410 ) ;
assign n40412 =  ( n1930 ) ? ( n40407 ) : ( n40411 ) ;
assign n40413 =  ( n879 ) ? ( n40402 ) : ( n40412 ) ;
assign n40414 =  ( n172 ) ? ( n19998 ) : ( VREG_1_2 ) ;
assign n40415 =  ( n170 ) ? ( n19997 ) : ( n40414 ) ;
assign n40416 =  ( n168 ) ? ( n19996 ) : ( n40415 ) ;
assign n40417 =  ( n166 ) ? ( n19995 ) : ( n40416 ) ;
assign n40418 =  ( n162 ) ? ( n19994 ) : ( n40417 ) ;
assign n40419 =  ( n172 ) ? ( n20008 ) : ( VREG_1_2 ) ;
assign n40420 =  ( n170 ) ? ( n20007 ) : ( n40419 ) ;
assign n40421 =  ( n168 ) ? ( n20006 ) : ( n40420 ) ;
assign n40422 =  ( n166 ) ? ( n20005 ) : ( n40421 ) ;
assign n40423 =  ( n162 ) ? ( n20004 ) : ( n40422 ) ;
assign n40424 =  ( n19987 ) ? ( VREG_1_2 ) : ( n40423 ) ;
assign n40425 =  ( n3051 ) ? ( n40424 ) : ( VREG_1_2 ) ;
assign n40426 =  ( n3040 ) ? ( n40418 ) : ( n40425 ) ;
assign n40427 =  ( n192 ) ? ( VREG_1_2 ) : ( VREG_1_2 ) ;
assign n40428 =  ( n157 ) ? ( n40426 ) : ( n40427 ) ;
assign n40429 =  ( n6 ) ? ( n40413 ) : ( n40428 ) ;
assign n40430 =  ( n197 ) ? ( n40429 ) : ( VREG_1_2 ) ;
assign n40431 =  ( n148 ) ? ( n21065 ) : ( VREG_1_3 ) ;
assign n40432 =  ( n146 ) ? ( n21064 ) : ( n40431 ) ;
assign n40433 =  ( n144 ) ? ( n21063 ) : ( n40432 ) ;
assign n40434 =  ( n142 ) ? ( n21062 ) : ( n40433 ) ;
assign n40435 =  ( n10 ) ? ( n21061 ) : ( n40434 ) ;
assign n40436 =  ( n148 ) ? ( n22099 ) : ( VREG_1_3 ) ;
assign n40437 =  ( n146 ) ? ( n22098 ) : ( n40436 ) ;
assign n40438 =  ( n144 ) ? ( n22097 ) : ( n40437 ) ;
assign n40439 =  ( n142 ) ? ( n22096 ) : ( n40438 ) ;
assign n40440 =  ( n10 ) ? ( n22095 ) : ( n40439 ) ;
assign n40441 =  ( n22106 ) ? ( VREG_1_3 ) : ( n40435 ) ;
assign n40442 =  ( n22106 ) ? ( VREG_1_3 ) : ( n40440 ) ;
assign n40443 =  ( n3034 ) ? ( n40442 ) : ( VREG_1_3 ) ;
assign n40444 =  ( n2965 ) ? ( n40441 ) : ( n40443 ) ;
assign n40445 =  ( n1930 ) ? ( n40440 ) : ( n40444 ) ;
assign n40446 =  ( n879 ) ? ( n40435 ) : ( n40445 ) ;
assign n40447 =  ( n172 ) ? ( n22117 ) : ( VREG_1_3 ) ;
assign n40448 =  ( n170 ) ? ( n22116 ) : ( n40447 ) ;
assign n40449 =  ( n168 ) ? ( n22115 ) : ( n40448 ) ;
assign n40450 =  ( n166 ) ? ( n22114 ) : ( n40449 ) ;
assign n40451 =  ( n162 ) ? ( n22113 ) : ( n40450 ) ;
assign n40452 =  ( n172 ) ? ( n22127 ) : ( VREG_1_3 ) ;
assign n40453 =  ( n170 ) ? ( n22126 ) : ( n40452 ) ;
assign n40454 =  ( n168 ) ? ( n22125 ) : ( n40453 ) ;
assign n40455 =  ( n166 ) ? ( n22124 ) : ( n40454 ) ;
assign n40456 =  ( n162 ) ? ( n22123 ) : ( n40455 ) ;
assign n40457 =  ( n22106 ) ? ( VREG_1_3 ) : ( n40456 ) ;
assign n40458 =  ( n3051 ) ? ( n40457 ) : ( VREG_1_3 ) ;
assign n40459 =  ( n3040 ) ? ( n40451 ) : ( n40458 ) ;
assign n40460 =  ( n192 ) ? ( VREG_1_3 ) : ( VREG_1_3 ) ;
assign n40461 =  ( n157 ) ? ( n40459 ) : ( n40460 ) ;
assign n40462 =  ( n6 ) ? ( n40446 ) : ( n40461 ) ;
assign n40463 =  ( n197 ) ? ( n40462 ) : ( VREG_1_3 ) ;
assign n40464 =  ( n148 ) ? ( n23184 ) : ( VREG_1_4 ) ;
assign n40465 =  ( n146 ) ? ( n23183 ) : ( n40464 ) ;
assign n40466 =  ( n144 ) ? ( n23182 ) : ( n40465 ) ;
assign n40467 =  ( n142 ) ? ( n23181 ) : ( n40466 ) ;
assign n40468 =  ( n10 ) ? ( n23180 ) : ( n40467 ) ;
assign n40469 =  ( n148 ) ? ( n24218 ) : ( VREG_1_4 ) ;
assign n40470 =  ( n146 ) ? ( n24217 ) : ( n40469 ) ;
assign n40471 =  ( n144 ) ? ( n24216 ) : ( n40470 ) ;
assign n40472 =  ( n142 ) ? ( n24215 ) : ( n40471 ) ;
assign n40473 =  ( n10 ) ? ( n24214 ) : ( n40472 ) ;
assign n40474 =  ( n24225 ) ? ( VREG_1_4 ) : ( n40468 ) ;
assign n40475 =  ( n24225 ) ? ( VREG_1_4 ) : ( n40473 ) ;
assign n40476 =  ( n3034 ) ? ( n40475 ) : ( VREG_1_4 ) ;
assign n40477 =  ( n2965 ) ? ( n40474 ) : ( n40476 ) ;
assign n40478 =  ( n1930 ) ? ( n40473 ) : ( n40477 ) ;
assign n40479 =  ( n879 ) ? ( n40468 ) : ( n40478 ) ;
assign n40480 =  ( n172 ) ? ( n24236 ) : ( VREG_1_4 ) ;
assign n40481 =  ( n170 ) ? ( n24235 ) : ( n40480 ) ;
assign n40482 =  ( n168 ) ? ( n24234 ) : ( n40481 ) ;
assign n40483 =  ( n166 ) ? ( n24233 ) : ( n40482 ) ;
assign n40484 =  ( n162 ) ? ( n24232 ) : ( n40483 ) ;
assign n40485 =  ( n172 ) ? ( n24246 ) : ( VREG_1_4 ) ;
assign n40486 =  ( n170 ) ? ( n24245 ) : ( n40485 ) ;
assign n40487 =  ( n168 ) ? ( n24244 ) : ( n40486 ) ;
assign n40488 =  ( n166 ) ? ( n24243 ) : ( n40487 ) ;
assign n40489 =  ( n162 ) ? ( n24242 ) : ( n40488 ) ;
assign n40490 =  ( n24225 ) ? ( VREG_1_4 ) : ( n40489 ) ;
assign n40491 =  ( n3051 ) ? ( n40490 ) : ( VREG_1_4 ) ;
assign n40492 =  ( n3040 ) ? ( n40484 ) : ( n40491 ) ;
assign n40493 =  ( n192 ) ? ( VREG_1_4 ) : ( VREG_1_4 ) ;
assign n40494 =  ( n157 ) ? ( n40492 ) : ( n40493 ) ;
assign n40495 =  ( n6 ) ? ( n40479 ) : ( n40494 ) ;
assign n40496 =  ( n197 ) ? ( n40495 ) : ( VREG_1_4 ) ;
assign n40497 =  ( n148 ) ? ( n25303 ) : ( VREG_1_5 ) ;
assign n40498 =  ( n146 ) ? ( n25302 ) : ( n40497 ) ;
assign n40499 =  ( n144 ) ? ( n25301 ) : ( n40498 ) ;
assign n40500 =  ( n142 ) ? ( n25300 ) : ( n40499 ) ;
assign n40501 =  ( n10 ) ? ( n25299 ) : ( n40500 ) ;
assign n40502 =  ( n148 ) ? ( n26337 ) : ( VREG_1_5 ) ;
assign n40503 =  ( n146 ) ? ( n26336 ) : ( n40502 ) ;
assign n40504 =  ( n144 ) ? ( n26335 ) : ( n40503 ) ;
assign n40505 =  ( n142 ) ? ( n26334 ) : ( n40504 ) ;
assign n40506 =  ( n10 ) ? ( n26333 ) : ( n40505 ) ;
assign n40507 =  ( n26344 ) ? ( VREG_1_5 ) : ( n40501 ) ;
assign n40508 =  ( n26344 ) ? ( VREG_1_5 ) : ( n40506 ) ;
assign n40509 =  ( n3034 ) ? ( n40508 ) : ( VREG_1_5 ) ;
assign n40510 =  ( n2965 ) ? ( n40507 ) : ( n40509 ) ;
assign n40511 =  ( n1930 ) ? ( n40506 ) : ( n40510 ) ;
assign n40512 =  ( n879 ) ? ( n40501 ) : ( n40511 ) ;
assign n40513 =  ( n172 ) ? ( n26355 ) : ( VREG_1_5 ) ;
assign n40514 =  ( n170 ) ? ( n26354 ) : ( n40513 ) ;
assign n40515 =  ( n168 ) ? ( n26353 ) : ( n40514 ) ;
assign n40516 =  ( n166 ) ? ( n26352 ) : ( n40515 ) ;
assign n40517 =  ( n162 ) ? ( n26351 ) : ( n40516 ) ;
assign n40518 =  ( n172 ) ? ( n26365 ) : ( VREG_1_5 ) ;
assign n40519 =  ( n170 ) ? ( n26364 ) : ( n40518 ) ;
assign n40520 =  ( n168 ) ? ( n26363 ) : ( n40519 ) ;
assign n40521 =  ( n166 ) ? ( n26362 ) : ( n40520 ) ;
assign n40522 =  ( n162 ) ? ( n26361 ) : ( n40521 ) ;
assign n40523 =  ( n26344 ) ? ( VREG_1_5 ) : ( n40522 ) ;
assign n40524 =  ( n3051 ) ? ( n40523 ) : ( VREG_1_5 ) ;
assign n40525 =  ( n3040 ) ? ( n40517 ) : ( n40524 ) ;
assign n40526 =  ( n192 ) ? ( VREG_1_5 ) : ( VREG_1_5 ) ;
assign n40527 =  ( n157 ) ? ( n40525 ) : ( n40526 ) ;
assign n40528 =  ( n6 ) ? ( n40512 ) : ( n40527 ) ;
assign n40529 =  ( n197 ) ? ( n40528 ) : ( VREG_1_5 ) ;
assign n40530 =  ( n148 ) ? ( n27422 ) : ( VREG_1_6 ) ;
assign n40531 =  ( n146 ) ? ( n27421 ) : ( n40530 ) ;
assign n40532 =  ( n144 ) ? ( n27420 ) : ( n40531 ) ;
assign n40533 =  ( n142 ) ? ( n27419 ) : ( n40532 ) ;
assign n40534 =  ( n10 ) ? ( n27418 ) : ( n40533 ) ;
assign n40535 =  ( n148 ) ? ( n28456 ) : ( VREG_1_6 ) ;
assign n40536 =  ( n146 ) ? ( n28455 ) : ( n40535 ) ;
assign n40537 =  ( n144 ) ? ( n28454 ) : ( n40536 ) ;
assign n40538 =  ( n142 ) ? ( n28453 ) : ( n40537 ) ;
assign n40539 =  ( n10 ) ? ( n28452 ) : ( n40538 ) ;
assign n40540 =  ( n28463 ) ? ( VREG_1_6 ) : ( n40534 ) ;
assign n40541 =  ( n28463 ) ? ( VREG_1_6 ) : ( n40539 ) ;
assign n40542 =  ( n3034 ) ? ( n40541 ) : ( VREG_1_6 ) ;
assign n40543 =  ( n2965 ) ? ( n40540 ) : ( n40542 ) ;
assign n40544 =  ( n1930 ) ? ( n40539 ) : ( n40543 ) ;
assign n40545 =  ( n879 ) ? ( n40534 ) : ( n40544 ) ;
assign n40546 =  ( n172 ) ? ( n28474 ) : ( VREG_1_6 ) ;
assign n40547 =  ( n170 ) ? ( n28473 ) : ( n40546 ) ;
assign n40548 =  ( n168 ) ? ( n28472 ) : ( n40547 ) ;
assign n40549 =  ( n166 ) ? ( n28471 ) : ( n40548 ) ;
assign n40550 =  ( n162 ) ? ( n28470 ) : ( n40549 ) ;
assign n40551 =  ( n172 ) ? ( n28484 ) : ( VREG_1_6 ) ;
assign n40552 =  ( n170 ) ? ( n28483 ) : ( n40551 ) ;
assign n40553 =  ( n168 ) ? ( n28482 ) : ( n40552 ) ;
assign n40554 =  ( n166 ) ? ( n28481 ) : ( n40553 ) ;
assign n40555 =  ( n162 ) ? ( n28480 ) : ( n40554 ) ;
assign n40556 =  ( n28463 ) ? ( VREG_1_6 ) : ( n40555 ) ;
assign n40557 =  ( n3051 ) ? ( n40556 ) : ( VREG_1_6 ) ;
assign n40558 =  ( n3040 ) ? ( n40550 ) : ( n40557 ) ;
assign n40559 =  ( n192 ) ? ( VREG_1_6 ) : ( VREG_1_6 ) ;
assign n40560 =  ( n157 ) ? ( n40558 ) : ( n40559 ) ;
assign n40561 =  ( n6 ) ? ( n40545 ) : ( n40560 ) ;
assign n40562 =  ( n197 ) ? ( n40561 ) : ( VREG_1_6 ) ;
assign n40563 =  ( n148 ) ? ( n29541 ) : ( VREG_1_7 ) ;
assign n40564 =  ( n146 ) ? ( n29540 ) : ( n40563 ) ;
assign n40565 =  ( n144 ) ? ( n29539 ) : ( n40564 ) ;
assign n40566 =  ( n142 ) ? ( n29538 ) : ( n40565 ) ;
assign n40567 =  ( n10 ) ? ( n29537 ) : ( n40566 ) ;
assign n40568 =  ( n148 ) ? ( n30575 ) : ( VREG_1_7 ) ;
assign n40569 =  ( n146 ) ? ( n30574 ) : ( n40568 ) ;
assign n40570 =  ( n144 ) ? ( n30573 ) : ( n40569 ) ;
assign n40571 =  ( n142 ) ? ( n30572 ) : ( n40570 ) ;
assign n40572 =  ( n10 ) ? ( n30571 ) : ( n40571 ) ;
assign n40573 =  ( n30582 ) ? ( VREG_1_7 ) : ( n40567 ) ;
assign n40574 =  ( n30582 ) ? ( VREG_1_7 ) : ( n40572 ) ;
assign n40575 =  ( n3034 ) ? ( n40574 ) : ( VREG_1_7 ) ;
assign n40576 =  ( n2965 ) ? ( n40573 ) : ( n40575 ) ;
assign n40577 =  ( n1930 ) ? ( n40572 ) : ( n40576 ) ;
assign n40578 =  ( n879 ) ? ( n40567 ) : ( n40577 ) ;
assign n40579 =  ( n172 ) ? ( n30593 ) : ( VREG_1_7 ) ;
assign n40580 =  ( n170 ) ? ( n30592 ) : ( n40579 ) ;
assign n40581 =  ( n168 ) ? ( n30591 ) : ( n40580 ) ;
assign n40582 =  ( n166 ) ? ( n30590 ) : ( n40581 ) ;
assign n40583 =  ( n162 ) ? ( n30589 ) : ( n40582 ) ;
assign n40584 =  ( n172 ) ? ( n30603 ) : ( VREG_1_7 ) ;
assign n40585 =  ( n170 ) ? ( n30602 ) : ( n40584 ) ;
assign n40586 =  ( n168 ) ? ( n30601 ) : ( n40585 ) ;
assign n40587 =  ( n166 ) ? ( n30600 ) : ( n40586 ) ;
assign n40588 =  ( n162 ) ? ( n30599 ) : ( n40587 ) ;
assign n40589 =  ( n30582 ) ? ( VREG_1_7 ) : ( n40588 ) ;
assign n40590 =  ( n3051 ) ? ( n40589 ) : ( VREG_1_7 ) ;
assign n40591 =  ( n3040 ) ? ( n40583 ) : ( n40590 ) ;
assign n40592 =  ( n192 ) ? ( VREG_1_7 ) : ( VREG_1_7 ) ;
assign n40593 =  ( n157 ) ? ( n40591 ) : ( n40592 ) ;
assign n40594 =  ( n6 ) ? ( n40578 ) : ( n40593 ) ;
assign n40595 =  ( n197 ) ? ( n40594 ) : ( VREG_1_7 ) ;
assign n40596 =  ( n148 ) ? ( n31660 ) : ( VREG_1_8 ) ;
assign n40597 =  ( n146 ) ? ( n31659 ) : ( n40596 ) ;
assign n40598 =  ( n144 ) ? ( n31658 ) : ( n40597 ) ;
assign n40599 =  ( n142 ) ? ( n31657 ) : ( n40598 ) ;
assign n40600 =  ( n10 ) ? ( n31656 ) : ( n40599 ) ;
assign n40601 =  ( n148 ) ? ( n32694 ) : ( VREG_1_8 ) ;
assign n40602 =  ( n146 ) ? ( n32693 ) : ( n40601 ) ;
assign n40603 =  ( n144 ) ? ( n32692 ) : ( n40602 ) ;
assign n40604 =  ( n142 ) ? ( n32691 ) : ( n40603 ) ;
assign n40605 =  ( n10 ) ? ( n32690 ) : ( n40604 ) ;
assign n40606 =  ( n32701 ) ? ( VREG_1_8 ) : ( n40600 ) ;
assign n40607 =  ( n32701 ) ? ( VREG_1_8 ) : ( n40605 ) ;
assign n40608 =  ( n3034 ) ? ( n40607 ) : ( VREG_1_8 ) ;
assign n40609 =  ( n2965 ) ? ( n40606 ) : ( n40608 ) ;
assign n40610 =  ( n1930 ) ? ( n40605 ) : ( n40609 ) ;
assign n40611 =  ( n879 ) ? ( n40600 ) : ( n40610 ) ;
assign n40612 =  ( n172 ) ? ( n32712 ) : ( VREG_1_8 ) ;
assign n40613 =  ( n170 ) ? ( n32711 ) : ( n40612 ) ;
assign n40614 =  ( n168 ) ? ( n32710 ) : ( n40613 ) ;
assign n40615 =  ( n166 ) ? ( n32709 ) : ( n40614 ) ;
assign n40616 =  ( n162 ) ? ( n32708 ) : ( n40615 ) ;
assign n40617 =  ( n172 ) ? ( n32722 ) : ( VREG_1_8 ) ;
assign n40618 =  ( n170 ) ? ( n32721 ) : ( n40617 ) ;
assign n40619 =  ( n168 ) ? ( n32720 ) : ( n40618 ) ;
assign n40620 =  ( n166 ) ? ( n32719 ) : ( n40619 ) ;
assign n40621 =  ( n162 ) ? ( n32718 ) : ( n40620 ) ;
assign n40622 =  ( n32701 ) ? ( VREG_1_8 ) : ( n40621 ) ;
assign n40623 =  ( n3051 ) ? ( n40622 ) : ( VREG_1_8 ) ;
assign n40624 =  ( n3040 ) ? ( n40616 ) : ( n40623 ) ;
assign n40625 =  ( n192 ) ? ( VREG_1_8 ) : ( VREG_1_8 ) ;
assign n40626 =  ( n157 ) ? ( n40624 ) : ( n40625 ) ;
assign n40627 =  ( n6 ) ? ( n40611 ) : ( n40626 ) ;
assign n40628 =  ( n197 ) ? ( n40627 ) : ( VREG_1_8 ) ;
assign n40629 =  ( n148 ) ? ( n33779 ) : ( VREG_1_9 ) ;
assign n40630 =  ( n146 ) ? ( n33778 ) : ( n40629 ) ;
assign n40631 =  ( n144 ) ? ( n33777 ) : ( n40630 ) ;
assign n40632 =  ( n142 ) ? ( n33776 ) : ( n40631 ) ;
assign n40633 =  ( n10 ) ? ( n33775 ) : ( n40632 ) ;
assign n40634 =  ( n148 ) ? ( n34813 ) : ( VREG_1_9 ) ;
assign n40635 =  ( n146 ) ? ( n34812 ) : ( n40634 ) ;
assign n40636 =  ( n144 ) ? ( n34811 ) : ( n40635 ) ;
assign n40637 =  ( n142 ) ? ( n34810 ) : ( n40636 ) ;
assign n40638 =  ( n10 ) ? ( n34809 ) : ( n40637 ) ;
assign n40639 =  ( n34820 ) ? ( VREG_1_9 ) : ( n40633 ) ;
assign n40640 =  ( n34820 ) ? ( VREG_1_9 ) : ( n40638 ) ;
assign n40641 =  ( n3034 ) ? ( n40640 ) : ( VREG_1_9 ) ;
assign n40642 =  ( n2965 ) ? ( n40639 ) : ( n40641 ) ;
assign n40643 =  ( n1930 ) ? ( n40638 ) : ( n40642 ) ;
assign n40644 =  ( n879 ) ? ( n40633 ) : ( n40643 ) ;
assign n40645 =  ( n172 ) ? ( n34831 ) : ( VREG_1_9 ) ;
assign n40646 =  ( n170 ) ? ( n34830 ) : ( n40645 ) ;
assign n40647 =  ( n168 ) ? ( n34829 ) : ( n40646 ) ;
assign n40648 =  ( n166 ) ? ( n34828 ) : ( n40647 ) ;
assign n40649 =  ( n162 ) ? ( n34827 ) : ( n40648 ) ;
assign n40650 =  ( n172 ) ? ( n34841 ) : ( VREG_1_9 ) ;
assign n40651 =  ( n170 ) ? ( n34840 ) : ( n40650 ) ;
assign n40652 =  ( n168 ) ? ( n34839 ) : ( n40651 ) ;
assign n40653 =  ( n166 ) ? ( n34838 ) : ( n40652 ) ;
assign n40654 =  ( n162 ) ? ( n34837 ) : ( n40653 ) ;
assign n40655 =  ( n34820 ) ? ( VREG_1_9 ) : ( n40654 ) ;
assign n40656 =  ( n3051 ) ? ( n40655 ) : ( VREG_1_9 ) ;
assign n40657 =  ( n3040 ) ? ( n40649 ) : ( n40656 ) ;
assign n40658 =  ( n192 ) ? ( VREG_1_9 ) : ( VREG_1_9 ) ;
assign n40659 =  ( n157 ) ? ( n40657 ) : ( n40658 ) ;
assign n40660 =  ( n6 ) ? ( n40644 ) : ( n40659 ) ;
assign n40661 =  ( n197 ) ? ( n40660 ) : ( VREG_1_9 ) ;
assign n40662 =  ( n148 ) ? ( n1924 ) : ( VREG_20_0 ) ;
assign n40663 =  ( n146 ) ? ( n1923 ) : ( n40662 ) ;
assign n40664 =  ( n144 ) ? ( n1922 ) : ( n40663 ) ;
assign n40665 =  ( n142 ) ? ( n1921 ) : ( n40664 ) ;
assign n40666 =  ( n10 ) ? ( n1920 ) : ( n40665 ) ;
assign n40667 =  ( n148 ) ? ( n2959 ) : ( VREG_20_0 ) ;
assign n40668 =  ( n146 ) ? ( n2958 ) : ( n40667 ) ;
assign n40669 =  ( n144 ) ? ( n2957 ) : ( n40668 ) ;
assign n40670 =  ( n142 ) ? ( n2956 ) : ( n40669 ) ;
assign n40671 =  ( n10 ) ? ( n2955 ) : ( n40670 ) ;
assign n40672 =  ( n3032 ) ? ( VREG_20_0 ) : ( n40666 ) ;
assign n40673 =  ( n3032 ) ? ( VREG_20_0 ) : ( n40671 ) ;
assign n40674 =  ( n3034 ) ? ( n40673 ) : ( VREG_20_0 ) ;
assign n40675 =  ( n2965 ) ? ( n40672 ) : ( n40674 ) ;
assign n40676 =  ( n1930 ) ? ( n40671 ) : ( n40675 ) ;
assign n40677 =  ( n879 ) ? ( n40666 ) : ( n40676 ) ;
assign n40678 =  ( n172 ) ? ( n3045 ) : ( VREG_20_0 ) ;
assign n40679 =  ( n170 ) ? ( n3044 ) : ( n40678 ) ;
assign n40680 =  ( n168 ) ? ( n3043 ) : ( n40679 ) ;
assign n40681 =  ( n166 ) ? ( n3042 ) : ( n40680 ) ;
assign n40682 =  ( n162 ) ? ( n3041 ) : ( n40681 ) ;
assign n40683 =  ( n172 ) ? ( n3056 ) : ( VREG_20_0 ) ;
assign n40684 =  ( n170 ) ? ( n3055 ) : ( n40683 ) ;
assign n40685 =  ( n168 ) ? ( n3054 ) : ( n40684 ) ;
assign n40686 =  ( n166 ) ? ( n3053 ) : ( n40685 ) ;
assign n40687 =  ( n162 ) ? ( n3052 ) : ( n40686 ) ;
assign n40688 =  ( n3032 ) ? ( VREG_20_0 ) : ( n40687 ) ;
assign n40689 =  ( n3051 ) ? ( n40688 ) : ( VREG_20_0 ) ;
assign n40690 =  ( n3040 ) ? ( n40682 ) : ( n40689 ) ;
assign n40691 =  ( n192 ) ? ( VREG_20_0 ) : ( VREG_20_0 ) ;
assign n40692 =  ( n157 ) ? ( n40690 ) : ( n40691 ) ;
assign n40693 =  ( n6 ) ? ( n40677 ) : ( n40692 ) ;
assign n40694 =  ( n461 ) ? ( n40693 ) : ( VREG_20_0 ) ;
assign n40695 =  ( n148 ) ? ( n4113 ) : ( VREG_20_1 ) ;
assign n40696 =  ( n146 ) ? ( n4112 ) : ( n40695 ) ;
assign n40697 =  ( n144 ) ? ( n4111 ) : ( n40696 ) ;
assign n40698 =  ( n142 ) ? ( n4110 ) : ( n40697 ) ;
assign n40699 =  ( n10 ) ? ( n4109 ) : ( n40698 ) ;
assign n40700 =  ( n148 ) ? ( n5147 ) : ( VREG_20_1 ) ;
assign n40701 =  ( n146 ) ? ( n5146 ) : ( n40700 ) ;
assign n40702 =  ( n144 ) ? ( n5145 ) : ( n40701 ) ;
assign n40703 =  ( n142 ) ? ( n5144 ) : ( n40702 ) ;
assign n40704 =  ( n10 ) ? ( n5143 ) : ( n40703 ) ;
assign n40705 =  ( n5154 ) ? ( VREG_20_1 ) : ( n40699 ) ;
assign n40706 =  ( n5154 ) ? ( VREG_20_1 ) : ( n40704 ) ;
assign n40707 =  ( n3034 ) ? ( n40706 ) : ( VREG_20_1 ) ;
assign n40708 =  ( n2965 ) ? ( n40705 ) : ( n40707 ) ;
assign n40709 =  ( n1930 ) ? ( n40704 ) : ( n40708 ) ;
assign n40710 =  ( n879 ) ? ( n40699 ) : ( n40709 ) ;
assign n40711 =  ( n172 ) ? ( n5165 ) : ( VREG_20_1 ) ;
assign n40712 =  ( n170 ) ? ( n5164 ) : ( n40711 ) ;
assign n40713 =  ( n168 ) ? ( n5163 ) : ( n40712 ) ;
assign n40714 =  ( n166 ) ? ( n5162 ) : ( n40713 ) ;
assign n40715 =  ( n162 ) ? ( n5161 ) : ( n40714 ) ;
assign n40716 =  ( n172 ) ? ( n5175 ) : ( VREG_20_1 ) ;
assign n40717 =  ( n170 ) ? ( n5174 ) : ( n40716 ) ;
assign n40718 =  ( n168 ) ? ( n5173 ) : ( n40717 ) ;
assign n40719 =  ( n166 ) ? ( n5172 ) : ( n40718 ) ;
assign n40720 =  ( n162 ) ? ( n5171 ) : ( n40719 ) ;
assign n40721 =  ( n5154 ) ? ( VREG_20_1 ) : ( n40720 ) ;
assign n40722 =  ( n3051 ) ? ( n40721 ) : ( VREG_20_1 ) ;
assign n40723 =  ( n3040 ) ? ( n40715 ) : ( n40722 ) ;
assign n40724 =  ( n192 ) ? ( VREG_20_1 ) : ( VREG_20_1 ) ;
assign n40725 =  ( n157 ) ? ( n40723 ) : ( n40724 ) ;
assign n40726 =  ( n6 ) ? ( n40710 ) : ( n40725 ) ;
assign n40727 =  ( n461 ) ? ( n40726 ) : ( VREG_20_1 ) ;
assign n40728 =  ( n148 ) ? ( n6232 ) : ( VREG_20_10 ) ;
assign n40729 =  ( n146 ) ? ( n6231 ) : ( n40728 ) ;
assign n40730 =  ( n144 ) ? ( n6230 ) : ( n40729 ) ;
assign n40731 =  ( n142 ) ? ( n6229 ) : ( n40730 ) ;
assign n40732 =  ( n10 ) ? ( n6228 ) : ( n40731 ) ;
assign n40733 =  ( n148 ) ? ( n7266 ) : ( VREG_20_10 ) ;
assign n40734 =  ( n146 ) ? ( n7265 ) : ( n40733 ) ;
assign n40735 =  ( n144 ) ? ( n7264 ) : ( n40734 ) ;
assign n40736 =  ( n142 ) ? ( n7263 ) : ( n40735 ) ;
assign n40737 =  ( n10 ) ? ( n7262 ) : ( n40736 ) ;
assign n40738 =  ( n7273 ) ? ( VREG_20_10 ) : ( n40732 ) ;
assign n40739 =  ( n7273 ) ? ( VREG_20_10 ) : ( n40737 ) ;
assign n40740 =  ( n3034 ) ? ( n40739 ) : ( VREG_20_10 ) ;
assign n40741 =  ( n2965 ) ? ( n40738 ) : ( n40740 ) ;
assign n40742 =  ( n1930 ) ? ( n40737 ) : ( n40741 ) ;
assign n40743 =  ( n879 ) ? ( n40732 ) : ( n40742 ) ;
assign n40744 =  ( n172 ) ? ( n7284 ) : ( VREG_20_10 ) ;
assign n40745 =  ( n170 ) ? ( n7283 ) : ( n40744 ) ;
assign n40746 =  ( n168 ) ? ( n7282 ) : ( n40745 ) ;
assign n40747 =  ( n166 ) ? ( n7281 ) : ( n40746 ) ;
assign n40748 =  ( n162 ) ? ( n7280 ) : ( n40747 ) ;
assign n40749 =  ( n172 ) ? ( n7294 ) : ( VREG_20_10 ) ;
assign n40750 =  ( n170 ) ? ( n7293 ) : ( n40749 ) ;
assign n40751 =  ( n168 ) ? ( n7292 ) : ( n40750 ) ;
assign n40752 =  ( n166 ) ? ( n7291 ) : ( n40751 ) ;
assign n40753 =  ( n162 ) ? ( n7290 ) : ( n40752 ) ;
assign n40754 =  ( n7273 ) ? ( VREG_20_10 ) : ( n40753 ) ;
assign n40755 =  ( n3051 ) ? ( n40754 ) : ( VREG_20_10 ) ;
assign n40756 =  ( n3040 ) ? ( n40748 ) : ( n40755 ) ;
assign n40757 =  ( n192 ) ? ( VREG_20_10 ) : ( VREG_20_10 ) ;
assign n40758 =  ( n157 ) ? ( n40756 ) : ( n40757 ) ;
assign n40759 =  ( n6 ) ? ( n40743 ) : ( n40758 ) ;
assign n40760 =  ( n461 ) ? ( n40759 ) : ( VREG_20_10 ) ;
assign n40761 =  ( n148 ) ? ( n8351 ) : ( VREG_20_11 ) ;
assign n40762 =  ( n146 ) ? ( n8350 ) : ( n40761 ) ;
assign n40763 =  ( n144 ) ? ( n8349 ) : ( n40762 ) ;
assign n40764 =  ( n142 ) ? ( n8348 ) : ( n40763 ) ;
assign n40765 =  ( n10 ) ? ( n8347 ) : ( n40764 ) ;
assign n40766 =  ( n148 ) ? ( n9385 ) : ( VREG_20_11 ) ;
assign n40767 =  ( n146 ) ? ( n9384 ) : ( n40766 ) ;
assign n40768 =  ( n144 ) ? ( n9383 ) : ( n40767 ) ;
assign n40769 =  ( n142 ) ? ( n9382 ) : ( n40768 ) ;
assign n40770 =  ( n10 ) ? ( n9381 ) : ( n40769 ) ;
assign n40771 =  ( n9392 ) ? ( VREG_20_11 ) : ( n40765 ) ;
assign n40772 =  ( n9392 ) ? ( VREG_20_11 ) : ( n40770 ) ;
assign n40773 =  ( n3034 ) ? ( n40772 ) : ( VREG_20_11 ) ;
assign n40774 =  ( n2965 ) ? ( n40771 ) : ( n40773 ) ;
assign n40775 =  ( n1930 ) ? ( n40770 ) : ( n40774 ) ;
assign n40776 =  ( n879 ) ? ( n40765 ) : ( n40775 ) ;
assign n40777 =  ( n172 ) ? ( n9403 ) : ( VREG_20_11 ) ;
assign n40778 =  ( n170 ) ? ( n9402 ) : ( n40777 ) ;
assign n40779 =  ( n168 ) ? ( n9401 ) : ( n40778 ) ;
assign n40780 =  ( n166 ) ? ( n9400 ) : ( n40779 ) ;
assign n40781 =  ( n162 ) ? ( n9399 ) : ( n40780 ) ;
assign n40782 =  ( n172 ) ? ( n9413 ) : ( VREG_20_11 ) ;
assign n40783 =  ( n170 ) ? ( n9412 ) : ( n40782 ) ;
assign n40784 =  ( n168 ) ? ( n9411 ) : ( n40783 ) ;
assign n40785 =  ( n166 ) ? ( n9410 ) : ( n40784 ) ;
assign n40786 =  ( n162 ) ? ( n9409 ) : ( n40785 ) ;
assign n40787 =  ( n9392 ) ? ( VREG_20_11 ) : ( n40786 ) ;
assign n40788 =  ( n3051 ) ? ( n40787 ) : ( VREG_20_11 ) ;
assign n40789 =  ( n3040 ) ? ( n40781 ) : ( n40788 ) ;
assign n40790 =  ( n192 ) ? ( VREG_20_11 ) : ( VREG_20_11 ) ;
assign n40791 =  ( n157 ) ? ( n40789 ) : ( n40790 ) ;
assign n40792 =  ( n6 ) ? ( n40776 ) : ( n40791 ) ;
assign n40793 =  ( n461 ) ? ( n40792 ) : ( VREG_20_11 ) ;
assign n40794 =  ( n148 ) ? ( n10470 ) : ( VREG_20_12 ) ;
assign n40795 =  ( n146 ) ? ( n10469 ) : ( n40794 ) ;
assign n40796 =  ( n144 ) ? ( n10468 ) : ( n40795 ) ;
assign n40797 =  ( n142 ) ? ( n10467 ) : ( n40796 ) ;
assign n40798 =  ( n10 ) ? ( n10466 ) : ( n40797 ) ;
assign n40799 =  ( n148 ) ? ( n11504 ) : ( VREG_20_12 ) ;
assign n40800 =  ( n146 ) ? ( n11503 ) : ( n40799 ) ;
assign n40801 =  ( n144 ) ? ( n11502 ) : ( n40800 ) ;
assign n40802 =  ( n142 ) ? ( n11501 ) : ( n40801 ) ;
assign n40803 =  ( n10 ) ? ( n11500 ) : ( n40802 ) ;
assign n40804 =  ( n11511 ) ? ( VREG_20_12 ) : ( n40798 ) ;
assign n40805 =  ( n11511 ) ? ( VREG_20_12 ) : ( n40803 ) ;
assign n40806 =  ( n3034 ) ? ( n40805 ) : ( VREG_20_12 ) ;
assign n40807 =  ( n2965 ) ? ( n40804 ) : ( n40806 ) ;
assign n40808 =  ( n1930 ) ? ( n40803 ) : ( n40807 ) ;
assign n40809 =  ( n879 ) ? ( n40798 ) : ( n40808 ) ;
assign n40810 =  ( n172 ) ? ( n11522 ) : ( VREG_20_12 ) ;
assign n40811 =  ( n170 ) ? ( n11521 ) : ( n40810 ) ;
assign n40812 =  ( n168 ) ? ( n11520 ) : ( n40811 ) ;
assign n40813 =  ( n166 ) ? ( n11519 ) : ( n40812 ) ;
assign n40814 =  ( n162 ) ? ( n11518 ) : ( n40813 ) ;
assign n40815 =  ( n172 ) ? ( n11532 ) : ( VREG_20_12 ) ;
assign n40816 =  ( n170 ) ? ( n11531 ) : ( n40815 ) ;
assign n40817 =  ( n168 ) ? ( n11530 ) : ( n40816 ) ;
assign n40818 =  ( n166 ) ? ( n11529 ) : ( n40817 ) ;
assign n40819 =  ( n162 ) ? ( n11528 ) : ( n40818 ) ;
assign n40820 =  ( n11511 ) ? ( VREG_20_12 ) : ( n40819 ) ;
assign n40821 =  ( n3051 ) ? ( n40820 ) : ( VREG_20_12 ) ;
assign n40822 =  ( n3040 ) ? ( n40814 ) : ( n40821 ) ;
assign n40823 =  ( n192 ) ? ( VREG_20_12 ) : ( VREG_20_12 ) ;
assign n40824 =  ( n157 ) ? ( n40822 ) : ( n40823 ) ;
assign n40825 =  ( n6 ) ? ( n40809 ) : ( n40824 ) ;
assign n40826 =  ( n461 ) ? ( n40825 ) : ( VREG_20_12 ) ;
assign n40827 =  ( n148 ) ? ( n12589 ) : ( VREG_20_13 ) ;
assign n40828 =  ( n146 ) ? ( n12588 ) : ( n40827 ) ;
assign n40829 =  ( n144 ) ? ( n12587 ) : ( n40828 ) ;
assign n40830 =  ( n142 ) ? ( n12586 ) : ( n40829 ) ;
assign n40831 =  ( n10 ) ? ( n12585 ) : ( n40830 ) ;
assign n40832 =  ( n148 ) ? ( n13623 ) : ( VREG_20_13 ) ;
assign n40833 =  ( n146 ) ? ( n13622 ) : ( n40832 ) ;
assign n40834 =  ( n144 ) ? ( n13621 ) : ( n40833 ) ;
assign n40835 =  ( n142 ) ? ( n13620 ) : ( n40834 ) ;
assign n40836 =  ( n10 ) ? ( n13619 ) : ( n40835 ) ;
assign n40837 =  ( n13630 ) ? ( VREG_20_13 ) : ( n40831 ) ;
assign n40838 =  ( n13630 ) ? ( VREG_20_13 ) : ( n40836 ) ;
assign n40839 =  ( n3034 ) ? ( n40838 ) : ( VREG_20_13 ) ;
assign n40840 =  ( n2965 ) ? ( n40837 ) : ( n40839 ) ;
assign n40841 =  ( n1930 ) ? ( n40836 ) : ( n40840 ) ;
assign n40842 =  ( n879 ) ? ( n40831 ) : ( n40841 ) ;
assign n40843 =  ( n172 ) ? ( n13641 ) : ( VREG_20_13 ) ;
assign n40844 =  ( n170 ) ? ( n13640 ) : ( n40843 ) ;
assign n40845 =  ( n168 ) ? ( n13639 ) : ( n40844 ) ;
assign n40846 =  ( n166 ) ? ( n13638 ) : ( n40845 ) ;
assign n40847 =  ( n162 ) ? ( n13637 ) : ( n40846 ) ;
assign n40848 =  ( n172 ) ? ( n13651 ) : ( VREG_20_13 ) ;
assign n40849 =  ( n170 ) ? ( n13650 ) : ( n40848 ) ;
assign n40850 =  ( n168 ) ? ( n13649 ) : ( n40849 ) ;
assign n40851 =  ( n166 ) ? ( n13648 ) : ( n40850 ) ;
assign n40852 =  ( n162 ) ? ( n13647 ) : ( n40851 ) ;
assign n40853 =  ( n13630 ) ? ( VREG_20_13 ) : ( n40852 ) ;
assign n40854 =  ( n3051 ) ? ( n40853 ) : ( VREG_20_13 ) ;
assign n40855 =  ( n3040 ) ? ( n40847 ) : ( n40854 ) ;
assign n40856 =  ( n192 ) ? ( VREG_20_13 ) : ( VREG_20_13 ) ;
assign n40857 =  ( n157 ) ? ( n40855 ) : ( n40856 ) ;
assign n40858 =  ( n6 ) ? ( n40842 ) : ( n40857 ) ;
assign n40859 =  ( n461 ) ? ( n40858 ) : ( VREG_20_13 ) ;
assign n40860 =  ( n148 ) ? ( n14708 ) : ( VREG_20_14 ) ;
assign n40861 =  ( n146 ) ? ( n14707 ) : ( n40860 ) ;
assign n40862 =  ( n144 ) ? ( n14706 ) : ( n40861 ) ;
assign n40863 =  ( n142 ) ? ( n14705 ) : ( n40862 ) ;
assign n40864 =  ( n10 ) ? ( n14704 ) : ( n40863 ) ;
assign n40865 =  ( n148 ) ? ( n15742 ) : ( VREG_20_14 ) ;
assign n40866 =  ( n146 ) ? ( n15741 ) : ( n40865 ) ;
assign n40867 =  ( n144 ) ? ( n15740 ) : ( n40866 ) ;
assign n40868 =  ( n142 ) ? ( n15739 ) : ( n40867 ) ;
assign n40869 =  ( n10 ) ? ( n15738 ) : ( n40868 ) ;
assign n40870 =  ( n15749 ) ? ( VREG_20_14 ) : ( n40864 ) ;
assign n40871 =  ( n15749 ) ? ( VREG_20_14 ) : ( n40869 ) ;
assign n40872 =  ( n3034 ) ? ( n40871 ) : ( VREG_20_14 ) ;
assign n40873 =  ( n2965 ) ? ( n40870 ) : ( n40872 ) ;
assign n40874 =  ( n1930 ) ? ( n40869 ) : ( n40873 ) ;
assign n40875 =  ( n879 ) ? ( n40864 ) : ( n40874 ) ;
assign n40876 =  ( n172 ) ? ( n15760 ) : ( VREG_20_14 ) ;
assign n40877 =  ( n170 ) ? ( n15759 ) : ( n40876 ) ;
assign n40878 =  ( n168 ) ? ( n15758 ) : ( n40877 ) ;
assign n40879 =  ( n166 ) ? ( n15757 ) : ( n40878 ) ;
assign n40880 =  ( n162 ) ? ( n15756 ) : ( n40879 ) ;
assign n40881 =  ( n172 ) ? ( n15770 ) : ( VREG_20_14 ) ;
assign n40882 =  ( n170 ) ? ( n15769 ) : ( n40881 ) ;
assign n40883 =  ( n168 ) ? ( n15768 ) : ( n40882 ) ;
assign n40884 =  ( n166 ) ? ( n15767 ) : ( n40883 ) ;
assign n40885 =  ( n162 ) ? ( n15766 ) : ( n40884 ) ;
assign n40886 =  ( n15749 ) ? ( VREG_20_14 ) : ( n40885 ) ;
assign n40887 =  ( n3051 ) ? ( n40886 ) : ( VREG_20_14 ) ;
assign n40888 =  ( n3040 ) ? ( n40880 ) : ( n40887 ) ;
assign n40889 =  ( n192 ) ? ( VREG_20_14 ) : ( VREG_20_14 ) ;
assign n40890 =  ( n157 ) ? ( n40888 ) : ( n40889 ) ;
assign n40891 =  ( n6 ) ? ( n40875 ) : ( n40890 ) ;
assign n40892 =  ( n461 ) ? ( n40891 ) : ( VREG_20_14 ) ;
assign n40893 =  ( n148 ) ? ( n16827 ) : ( VREG_20_15 ) ;
assign n40894 =  ( n146 ) ? ( n16826 ) : ( n40893 ) ;
assign n40895 =  ( n144 ) ? ( n16825 ) : ( n40894 ) ;
assign n40896 =  ( n142 ) ? ( n16824 ) : ( n40895 ) ;
assign n40897 =  ( n10 ) ? ( n16823 ) : ( n40896 ) ;
assign n40898 =  ( n148 ) ? ( n17861 ) : ( VREG_20_15 ) ;
assign n40899 =  ( n146 ) ? ( n17860 ) : ( n40898 ) ;
assign n40900 =  ( n144 ) ? ( n17859 ) : ( n40899 ) ;
assign n40901 =  ( n142 ) ? ( n17858 ) : ( n40900 ) ;
assign n40902 =  ( n10 ) ? ( n17857 ) : ( n40901 ) ;
assign n40903 =  ( n17868 ) ? ( VREG_20_15 ) : ( n40897 ) ;
assign n40904 =  ( n17868 ) ? ( VREG_20_15 ) : ( n40902 ) ;
assign n40905 =  ( n3034 ) ? ( n40904 ) : ( VREG_20_15 ) ;
assign n40906 =  ( n2965 ) ? ( n40903 ) : ( n40905 ) ;
assign n40907 =  ( n1930 ) ? ( n40902 ) : ( n40906 ) ;
assign n40908 =  ( n879 ) ? ( n40897 ) : ( n40907 ) ;
assign n40909 =  ( n172 ) ? ( n17879 ) : ( VREG_20_15 ) ;
assign n40910 =  ( n170 ) ? ( n17878 ) : ( n40909 ) ;
assign n40911 =  ( n168 ) ? ( n17877 ) : ( n40910 ) ;
assign n40912 =  ( n166 ) ? ( n17876 ) : ( n40911 ) ;
assign n40913 =  ( n162 ) ? ( n17875 ) : ( n40912 ) ;
assign n40914 =  ( n172 ) ? ( n17889 ) : ( VREG_20_15 ) ;
assign n40915 =  ( n170 ) ? ( n17888 ) : ( n40914 ) ;
assign n40916 =  ( n168 ) ? ( n17887 ) : ( n40915 ) ;
assign n40917 =  ( n166 ) ? ( n17886 ) : ( n40916 ) ;
assign n40918 =  ( n162 ) ? ( n17885 ) : ( n40917 ) ;
assign n40919 =  ( n17868 ) ? ( VREG_20_15 ) : ( n40918 ) ;
assign n40920 =  ( n3051 ) ? ( n40919 ) : ( VREG_20_15 ) ;
assign n40921 =  ( n3040 ) ? ( n40913 ) : ( n40920 ) ;
assign n40922 =  ( n192 ) ? ( VREG_20_15 ) : ( VREG_20_15 ) ;
assign n40923 =  ( n157 ) ? ( n40921 ) : ( n40922 ) ;
assign n40924 =  ( n6 ) ? ( n40908 ) : ( n40923 ) ;
assign n40925 =  ( n461 ) ? ( n40924 ) : ( VREG_20_15 ) ;
assign n40926 =  ( n148 ) ? ( n18946 ) : ( VREG_20_2 ) ;
assign n40927 =  ( n146 ) ? ( n18945 ) : ( n40926 ) ;
assign n40928 =  ( n144 ) ? ( n18944 ) : ( n40927 ) ;
assign n40929 =  ( n142 ) ? ( n18943 ) : ( n40928 ) ;
assign n40930 =  ( n10 ) ? ( n18942 ) : ( n40929 ) ;
assign n40931 =  ( n148 ) ? ( n19980 ) : ( VREG_20_2 ) ;
assign n40932 =  ( n146 ) ? ( n19979 ) : ( n40931 ) ;
assign n40933 =  ( n144 ) ? ( n19978 ) : ( n40932 ) ;
assign n40934 =  ( n142 ) ? ( n19977 ) : ( n40933 ) ;
assign n40935 =  ( n10 ) ? ( n19976 ) : ( n40934 ) ;
assign n40936 =  ( n19987 ) ? ( VREG_20_2 ) : ( n40930 ) ;
assign n40937 =  ( n19987 ) ? ( VREG_20_2 ) : ( n40935 ) ;
assign n40938 =  ( n3034 ) ? ( n40937 ) : ( VREG_20_2 ) ;
assign n40939 =  ( n2965 ) ? ( n40936 ) : ( n40938 ) ;
assign n40940 =  ( n1930 ) ? ( n40935 ) : ( n40939 ) ;
assign n40941 =  ( n879 ) ? ( n40930 ) : ( n40940 ) ;
assign n40942 =  ( n172 ) ? ( n19998 ) : ( VREG_20_2 ) ;
assign n40943 =  ( n170 ) ? ( n19997 ) : ( n40942 ) ;
assign n40944 =  ( n168 ) ? ( n19996 ) : ( n40943 ) ;
assign n40945 =  ( n166 ) ? ( n19995 ) : ( n40944 ) ;
assign n40946 =  ( n162 ) ? ( n19994 ) : ( n40945 ) ;
assign n40947 =  ( n172 ) ? ( n20008 ) : ( VREG_20_2 ) ;
assign n40948 =  ( n170 ) ? ( n20007 ) : ( n40947 ) ;
assign n40949 =  ( n168 ) ? ( n20006 ) : ( n40948 ) ;
assign n40950 =  ( n166 ) ? ( n20005 ) : ( n40949 ) ;
assign n40951 =  ( n162 ) ? ( n20004 ) : ( n40950 ) ;
assign n40952 =  ( n19987 ) ? ( VREG_20_2 ) : ( n40951 ) ;
assign n40953 =  ( n3051 ) ? ( n40952 ) : ( VREG_20_2 ) ;
assign n40954 =  ( n3040 ) ? ( n40946 ) : ( n40953 ) ;
assign n40955 =  ( n192 ) ? ( VREG_20_2 ) : ( VREG_20_2 ) ;
assign n40956 =  ( n157 ) ? ( n40954 ) : ( n40955 ) ;
assign n40957 =  ( n6 ) ? ( n40941 ) : ( n40956 ) ;
assign n40958 =  ( n461 ) ? ( n40957 ) : ( VREG_20_2 ) ;
assign n40959 =  ( n148 ) ? ( n21065 ) : ( VREG_20_3 ) ;
assign n40960 =  ( n146 ) ? ( n21064 ) : ( n40959 ) ;
assign n40961 =  ( n144 ) ? ( n21063 ) : ( n40960 ) ;
assign n40962 =  ( n142 ) ? ( n21062 ) : ( n40961 ) ;
assign n40963 =  ( n10 ) ? ( n21061 ) : ( n40962 ) ;
assign n40964 =  ( n148 ) ? ( n22099 ) : ( VREG_20_3 ) ;
assign n40965 =  ( n146 ) ? ( n22098 ) : ( n40964 ) ;
assign n40966 =  ( n144 ) ? ( n22097 ) : ( n40965 ) ;
assign n40967 =  ( n142 ) ? ( n22096 ) : ( n40966 ) ;
assign n40968 =  ( n10 ) ? ( n22095 ) : ( n40967 ) ;
assign n40969 =  ( n22106 ) ? ( VREG_20_3 ) : ( n40963 ) ;
assign n40970 =  ( n22106 ) ? ( VREG_20_3 ) : ( n40968 ) ;
assign n40971 =  ( n3034 ) ? ( n40970 ) : ( VREG_20_3 ) ;
assign n40972 =  ( n2965 ) ? ( n40969 ) : ( n40971 ) ;
assign n40973 =  ( n1930 ) ? ( n40968 ) : ( n40972 ) ;
assign n40974 =  ( n879 ) ? ( n40963 ) : ( n40973 ) ;
assign n40975 =  ( n172 ) ? ( n22117 ) : ( VREG_20_3 ) ;
assign n40976 =  ( n170 ) ? ( n22116 ) : ( n40975 ) ;
assign n40977 =  ( n168 ) ? ( n22115 ) : ( n40976 ) ;
assign n40978 =  ( n166 ) ? ( n22114 ) : ( n40977 ) ;
assign n40979 =  ( n162 ) ? ( n22113 ) : ( n40978 ) ;
assign n40980 =  ( n172 ) ? ( n22127 ) : ( VREG_20_3 ) ;
assign n40981 =  ( n170 ) ? ( n22126 ) : ( n40980 ) ;
assign n40982 =  ( n168 ) ? ( n22125 ) : ( n40981 ) ;
assign n40983 =  ( n166 ) ? ( n22124 ) : ( n40982 ) ;
assign n40984 =  ( n162 ) ? ( n22123 ) : ( n40983 ) ;
assign n40985 =  ( n22106 ) ? ( VREG_20_3 ) : ( n40984 ) ;
assign n40986 =  ( n3051 ) ? ( n40985 ) : ( VREG_20_3 ) ;
assign n40987 =  ( n3040 ) ? ( n40979 ) : ( n40986 ) ;
assign n40988 =  ( n192 ) ? ( VREG_20_3 ) : ( VREG_20_3 ) ;
assign n40989 =  ( n157 ) ? ( n40987 ) : ( n40988 ) ;
assign n40990 =  ( n6 ) ? ( n40974 ) : ( n40989 ) ;
assign n40991 =  ( n461 ) ? ( n40990 ) : ( VREG_20_3 ) ;
assign n40992 =  ( n148 ) ? ( n23184 ) : ( VREG_20_4 ) ;
assign n40993 =  ( n146 ) ? ( n23183 ) : ( n40992 ) ;
assign n40994 =  ( n144 ) ? ( n23182 ) : ( n40993 ) ;
assign n40995 =  ( n142 ) ? ( n23181 ) : ( n40994 ) ;
assign n40996 =  ( n10 ) ? ( n23180 ) : ( n40995 ) ;
assign n40997 =  ( n148 ) ? ( n24218 ) : ( VREG_20_4 ) ;
assign n40998 =  ( n146 ) ? ( n24217 ) : ( n40997 ) ;
assign n40999 =  ( n144 ) ? ( n24216 ) : ( n40998 ) ;
assign n41000 =  ( n142 ) ? ( n24215 ) : ( n40999 ) ;
assign n41001 =  ( n10 ) ? ( n24214 ) : ( n41000 ) ;
assign n41002 =  ( n24225 ) ? ( VREG_20_4 ) : ( n40996 ) ;
assign n41003 =  ( n24225 ) ? ( VREG_20_4 ) : ( n41001 ) ;
assign n41004 =  ( n3034 ) ? ( n41003 ) : ( VREG_20_4 ) ;
assign n41005 =  ( n2965 ) ? ( n41002 ) : ( n41004 ) ;
assign n41006 =  ( n1930 ) ? ( n41001 ) : ( n41005 ) ;
assign n41007 =  ( n879 ) ? ( n40996 ) : ( n41006 ) ;
assign n41008 =  ( n172 ) ? ( n24236 ) : ( VREG_20_4 ) ;
assign n41009 =  ( n170 ) ? ( n24235 ) : ( n41008 ) ;
assign n41010 =  ( n168 ) ? ( n24234 ) : ( n41009 ) ;
assign n41011 =  ( n166 ) ? ( n24233 ) : ( n41010 ) ;
assign n41012 =  ( n162 ) ? ( n24232 ) : ( n41011 ) ;
assign n41013 =  ( n172 ) ? ( n24246 ) : ( VREG_20_4 ) ;
assign n41014 =  ( n170 ) ? ( n24245 ) : ( n41013 ) ;
assign n41015 =  ( n168 ) ? ( n24244 ) : ( n41014 ) ;
assign n41016 =  ( n166 ) ? ( n24243 ) : ( n41015 ) ;
assign n41017 =  ( n162 ) ? ( n24242 ) : ( n41016 ) ;
assign n41018 =  ( n24225 ) ? ( VREG_20_4 ) : ( n41017 ) ;
assign n41019 =  ( n3051 ) ? ( n41018 ) : ( VREG_20_4 ) ;
assign n41020 =  ( n3040 ) ? ( n41012 ) : ( n41019 ) ;
assign n41021 =  ( n192 ) ? ( VREG_20_4 ) : ( VREG_20_4 ) ;
assign n41022 =  ( n157 ) ? ( n41020 ) : ( n41021 ) ;
assign n41023 =  ( n6 ) ? ( n41007 ) : ( n41022 ) ;
assign n41024 =  ( n461 ) ? ( n41023 ) : ( VREG_20_4 ) ;
assign n41025 =  ( n148 ) ? ( n25303 ) : ( VREG_20_5 ) ;
assign n41026 =  ( n146 ) ? ( n25302 ) : ( n41025 ) ;
assign n41027 =  ( n144 ) ? ( n25301 ) : ( n41026 ) ;
assign n41028 =  ( n142 ) ? ( n25300 ) : ( n41027 ) ;
assign n41029 =  ( n10 ) ? ( n25299 ) : ( n41028 ) ;
assign n41030 =  ( n148 ) ? ( n26337 ) : ( VREG_20_5 ) ;
assign n41031 =  ( n146 ) ? ( n26336 ) : ( n41030 ) ;
assign n41032 =  ( n144 ) ? ( n26335 ) : ( n41031 ) ;
assign n41033 =  ( n142 ) ? ( n26334 ) : ( n41032 ) ;
assign n41034 =  ( n10 ) ? ( n26333 ) : ( n41033 ) ;
assign n41035 =  ( n26344 ) ? ( VREG_20_5 ) : ( n41029 ) ;
assign n41036 =  ( n26344 ) ? ( VREG_20_5 ) : ( n41034 ) ;
assign n41037 =  ( n3034 ) ? ( n41036 ) : ( VREG_20_5 ) ;
assign n41038 =  ( n2965 ) ? ( n41035 ) : ( n41037 ) ;
assign n41039 =  ( n1930 ) ? ( n41034 ) : ( n41038 ) ;
assign n41040 =  ( n879 ) ? ( n41029 ) : ( n41039 ) ;
assign n41041 =  ( n172 ) ? ( n26355 ) : ( VREG_20_5 ) ;
assign n41042 =  ( n170 ) ? ( n26354 ) : ( n41041 ) ;
assign n41043 =  ( n168 ) ? ( n26353 ) : ( n41042 ) ;
assign n41044 =  ( n166 ) ? ( n26352 ) : ( n41043 ) ;
assign n41045 =  ( n162 ) ? ( n26351 ) : ( n41044 ) ;
assign n41046 =  ( n172 ) ? ( n26365 ) : ( VREG_20_5 ) ;
assign n41047 =  ( n170 ) ? ( n26364 ) : ( n41046 ) ;
assign n41048 =  ( n168 ) ? ( n26363 ) : ( n41047 ) ;
assign n41049 =  ( n166 ) ? ( n26362 ) : ( n41048 ) ;
assign n41050 =  ( n162 ) ? ( n26361 ) : ( n41049 ) ;
assign n41051 =  ( n26344 ) ? ( VREG_20_5 ) : ( n41050 ) ;
assign n41052 =  ( n3051 ) ? ( n41051 ) : ( VREG_20_5 ) ;
assign n41053 =  ( n3040 ) ? ( n41045 ) : ( n41052 ) ;
assign n41054 =  ( n192 ) ? ( VREG_20_5 ) : ( VREG_20_5 ) ;
assign n41055 =  ( n157 ) ? ( n41053 ) : ( n41054 ) ;
assign n41056 =  ( n6 ) ? ( n41040 ) : ( n41055 ) ;
assign n41057 =  ( n461 ) ? ( n41056 ) : ( VREG_20_5 ) ;
assign n41058 =  ( n148 ) ? ( n27422 ) : ( VREG_20_6 ) ;
assign n41059 =  ( n146 ) ? ( n27421 ) : ( n41058 ) ;
assign n41060 =  ( n144 ) ? ( n27420 ) : ( n41059 ) ;
assign n41061 =  ( n142 ) ? ( n27419 ) : ( n41060 ) ;
assign n41062 =  ( n10 ) ? ( n27418 ) : ( n41061 ) ;
assign n41063 =  ( n148 ) ? ( n28456 ) : ( VREG_20_6 ) ;
assign n41064 =  ( n146 ) ? ( n28455 ) : ( n41063 ) ;
assign n41065 =  ( n144 ) ? ( n28454 ) : ( n41064 ) ;
assign n41066 =  ( n142 ) ? ( n28453 ) : ( n41065 ) ;
assign n41067 =  ( n10 ) ? ( n28452 ) : ( n41066 ) ;
assign n41068 =  ( n28463 ) ? ( VREG_20_6 ) : ( n41062 ) ;
assign n41069 =  ( n28463 ) ? ( VREG_20_6 ) : ( n41067 ) ;
assign n41070 =  ( n3034 ) ? ( n41069 ) : ( VREG_20_6 ) ;
assign n41071 =  ( n2965 ) ? ( n41068 ) : ( n41070 ) ;
assign n41072 =  ( n1930 ) ? ( n41067 ) : ( n41071 ) ;
assign n41073 =  ( n879 ) ? ( n41062 ) : ( n41072 ) ;
assign n41074 =  ( n172 ) ? ( n28474 ) : ( VREG_20_6 ) ;
assign n41075 =  ( n170 ) ? ( n28473 ) : ( n41074 ) ;
assign n41076 =  ( n168 ) ? ( n28472 ) : ( n41075 ) ;
assign n41077 =  ( n166 ) ? ( n28471 ) : ( n41076 ) ;
assign n41078 =  ( n162 ) ? ( n28470 ) : ( n41077 ) ;
assign n41079 =  ( n172 ) ? ( n28484 ) : ( VREG_20_6 ) ;
assign n41080 =  ( n170 ) ? ( n28483 ) : ( n41079 ) ;
assign n41081 =  ( n168 ) ? ( n28482 ) : ( n41080 ) ;
assign n41082 =  ( n166 ) ? ( n28481 ) : ( n41081 ) ;
assign n41083 =  ( n162 ) ? ( n28480 ) : ( n41082 ) ;
assign n41084 =  ( n28463 ) ? ( VREG_20_6 ) : ( n41083 ) ;
assign n41085 =  ( n3051 ) ? ( n41084 ) : ( VREG_20_6 ) ;
assign n41086 =  ( n3040 ) ? ( n41078 ) : ( n41085 ) ;
assign n41087 =  ( n192 ) ? ( VREG_20_6 ) : ( VREG_20_6 ) ;
assign n41088 =  ( n157 ) ? ( n41086 ) : ( n41087 ) ;
assign n41089 =  ( n6 ) ? ( n41073 ) : ( n41088 ) ;
assign n41090 =  ( n461 ) ? ( n41089 ) : ( VREG_20_6 ) ;
assign n41091 =  ( n148 ) ? ( n29541 ) : ( VREG_20_7 ) ;
assign n41092 =  ( n146 ) ? ( n29540 ) : ( n41091 ) ;
assign n41093 =  ( n144 ) ? ( n29539 ) : ( n41092 ) ;
assign n41094 =  ( n142 ) ? ( n29538 ) : ( n41093 ) ;
assign n41095 =  ( n10 ) ? ( n29537 ) : ( n41094 ) ;
assign n41096 =  ( n148 ) ? ( n30575 ) : ( VREG_20_7 ) ;
assign n41097 =  ( n146 ) ? ( n30574 ) : ( n41096 ) ;
assign n41098 =  ( n144 ) ? ( n30573 ) : ( n41097 ) ;
assign n41099 =  ( n142 ) ? ( n30572 ) : ( n41098 ) ;
assign n41100 =  ( n10 ) ? ( n30571 ) : ( n41099 ) ;
assign n41101 =  ( n30582 ) ? ( VREG_20_7 ) : ( n41095 ) ;
assign n41102 =  ( n30582 ) ? ( VREG_20_7 ) : ( n41100 ) ;
assign n41103 =  ( n3034 ) ? ( n41102 ) : ( VREG_20_7 ) ;
assign n41104 =  ( n2965 ) ? ( n41101 ) : ( n41103 ) ;
assign n41105 =  ( n1930 ) ? ( n41100 ) : ( n41104 ) ;
assign n41106 =  ( n879 ) ? ( n41095 ) : ( n41105 ) ;
assign n41107 =  ( n172 ) ? ( n30593 ) : ( VREG_20_7 ) ;
assign n41108 =  ( n170 ) ? ( n30592 ) : ( n41107 ) ;
assign n41109 =  ( n168 ) ? ( n30591 ) : ( n41108 ) ;
assign n41110 =  ( n166 ) ? ( n30590 ) : ( n41109 ) ;
assign n41111 =  ( n162 ) ? ( n30589 ) : ( n41110 ) ;
assign n41112 =  ( n172 ) ? ( n30603 ) : ( VREG_20_7 ) ;
assign n41113 =  ( n170 ) ? ( n30602 ) : ( n41112 ) ;
assign n41114 =  ( n168 ) ? ( n30601 ) : ( n41113 ) ;
assign n41115 =  ( n166 ) ? ( n30600 ) : ( n41114 ) ;
assign n41116 =  ( n162 ) ? ( n30599 ) : ( n41115 ) ;
assign n41117 =  ( n30582 ) ? ( VREG_20_7 ) : ( n41116 ) ;
assign n41118 =  ( n3051 ) ? ( n41117 ) : ( VREG_20_7 ) ;
assign n41119 =  ( n3040 ) ? ( n41111 ) : ( n41118 ) ;
assign n41120 =  ( n192 ) ? ( VREG_20_7 ) : ( VREG_20_7 ) ;
assign n41121 =  ( n157 ) ? ( n41119 ) : ( n41120 ) ;
assign n41122 =  ( n6 ) ? ( n41106 ) : ( n41121 ) ;
assign n41123 =  ( n461 ) ? ( n41122 ) : ( VREG_20_7 ) ;
assign n41124 =  ( n148 ) ? ( n31660 ) : ( VREG_20_8 ) ;
assign n41125 =  ( n146 ) ? ( n31659 ) : ( n41124 ) ;
assign n41126 =  ( n144 ) ? ( n31658 ) : ( n41125 ) ;
assign n41127 =  ( n142 ) ? ( n31657 ) : ( n41126 ) ;
assign n41128 =  ( n10 ) ? ( n31656 ) : ( n41127 ) ;
assign n41129 =  ( n148 ) ? ( n32694 ) : ( VREG_20_8 ) ;
assign n41130 =  ( n146 ) ? ( n32693 ) : ( n41129 ) ;
assign n41131 =  ( n144 ) ? ( n32692 ) : ( n41130 ) ;
assign n41132 =  ( n142 ) ? ( n32691 ) : ( n41131 ) ;
assign n41133 =  ( n10 ) ? ( n32690 ) : ( n41132 ) ;
assign n41134 =  ( n32701 ) ? ( VREG_20_8 ) : ( n41128 ) ;
assign n41135 =  ( n32701 ) ? ( VREG_20_8 ) : ( n41133 ) ;
assign n41136 =  ( n3034 ) ? ( n41135 ) : ( VREG_20_8 ) ;
assign n41137 =  ( n2965 ) ? ( n41134 ) : ( n41136 ) ;
assign n41138 =  ( n1930 ) ? ( n41133 ) : ( n41137 ) ;
assign n41139 =  ( n879 ) ? ( n41128 ) : ( n41138 ) ;
assign n41140 =  ( n172 ) ? ( n32712 ) : ( VREG_20_8 ) ;
assign n41141 =  ( n170 ) ? ( n32711 ) : ( n41140 ) ;
assign n41142 =  ( n168 ) ? ( n32710 ) : ( n41141 ) ;
assign n41143 =  ( n166 ) ? ( n32709 ) : ( n41142 ) ;
assign n41144 =  ( n162 ) ? ( n32708 ) : ( n41143 ) ;
assign n41145 =  ( n172 ) ? ( n32722 ) : ( VREG_20_8 ) ;
assign n41146 =  ( n170 ) ? ( n32721 ) : ( n41145 ) ;
assign n41147 =  ( n168 ) ? ( n32720 ) : ( n41146 ) ;
assign n41148 =  ( n166 ) ? ( n32719 ) : ( n41147 ) ;
assign n41149 =  ( n162 ) ? ( n32718 ) : ( n41148 ) ;
assign n41150 =  ( n32701 ) ? ( VREG_20_8 ) : ( n41149 ) ;
assign n41151 =  ( n3051 ) ? ( n41150 ) : ( VREG_20_8 ) ;
assign n41152 =  ( n3040 ) ? ( n41144 ) : ( n41151 ) ;
assign n41153 =  ( n192 ) ? ( VREG_20_8 ) : ( VREG_20_8 ) ;
assign n41154 =  ( n157 ) ? ( n41152 ) : ( n41153 ) ;
assign n41155 =  ( n6 ) ? ( n41139 ) : ( n41154 ) ;
assign n41156 =  ( n461 ) ? ( n41155 ) : ( VREG_20_8 ) ;
assign n41157 =  ( n148 ) ? ( n33779 ) : ( VREG_20_9 ) ;
assign n41158 =  ( n146 ) ? ( n33778 ) : ( n41157 ) ;
assign n41159 =  ( n144 ) ? ( n33777 ) : ( n41158 ) ;
assign n41160 =  ( n142 ) ? ( n33776 ) : ( n41159 ) ;
assign n41161 =  ( n10 ) ? ( n33775 ) : ( n41160 ) ;
assign n41162 =  ( n148 ) ? ( n34813 ) : ( VREG_20_9 ) ;
assign n41163 =  ( n146 ) ? ( n34812 ) : ( n41162 ) ;
assign n41164 =  ( n144 ) ? ( n34811 ) : ( n41163 ) ;
assign n41165 =  ( n142 ) ? ( n34810 ) : ( n41164 ) ;
assign n41166 =  ( n10 ) ? ( n34809 ) : ( n41165 ) ;
assign n41167 =  ( n34820 ) ? ( VREG_20_9 ) : ( n41161 ) ;
assign n41168 =  ( n34820 ) ? ( VREG_20_9 ) : ( n41166 ) ;
assign n41169 =  ( n3034 ) ? ( n41168 ) : ( VREG_20_9 ) ;
assign n41170 =  ( n2965 ) ? ( n41167 ) : ( n41169 ) ;
assign n41171 =  ( n1930 ) ? ( n41166 ) : ( n41170 ) ;
assign n41172 =  ( n879 ) ? ( n41161 ) : ( n41171 ) ;
assign n41173 =  ( n172 ) ? ( n34831 ) : ( VREG_20_9 ) ;
assign n41174 =  ( n170 ) ? ( n34830 ) : ( n41173 ) ;
assign n41175 =  ( n168 ) ? ( n34829 ) : ( n41174 ) ;
assign n41176 =  ( n166 ) ? ( n34828 ) : ( n41175 ) ;
assign n41177 =  ( n162 ) ? ( n34827 ) : ( n41176 ) ;
assign n41178 =  ( n172 ) ? ( n34841 ) : ( VREG_20_9 ) ;
assign n41179 =  ( n170 ) ? ( n34840 ) : ( n41178 ) ;
assign n41180 =  ( n168 ) ? ( n34839 ) : ( n41179 ) ;
assign n41181 =  ( n166 ) ? ( n34838 ) : ( n41180 ) ;
assign n41182 =  ( n162 ) ? ( n34837 ) : ( n41181 ) ;
assign n41183 =  ( n34820 ) ? ( VREG_20_9 ) : ( n41182 ) ;
assign n41184 =  ( n3051 ) ? ( n41183 ) : ( VREG_20_9 ) ;
assign n41185 =  ( n3040 ) ? ( n41177 ) : ( n41184 ) ;
assign n41186 =  ( n192 ) ? ( VREG_20_9 ) : ( VREG_20_9 ) ;
assign n41187 =  ( n157 ) ? ( n41185 ) : ( n41186 ) ;
assign n41188 =  ( n6 ) ? ( n41172 ) : ( n41187 ) ;
assign n41189 =  ( n461 ) ? ( n41188 ) : ( VREG_20_9 ) ;
assign n41190 =  ( n148 ) ? ( n1924 ) : ( VREG_21_0 ) ;
assign n41191 =  ( n146 ) ? ( n1923 ) : ( n41190 ) ;
assign n41192 =  ( n144 ) ? ( n1922 ) : ( n41191 ) ;
assign n41193 =  ( n142 ) ? ( n1921 ) : ( n41192 ) ;
assign n41194 =  ( n10 ) ? ( n1920 ) : ( n41193 ) ;
assign n41195 =  ( n148 ) ? ( n2959 ) : ( VREG_21_0 ) ;
assign n41196 =  ( n146 ) ? ( n2958 ) : ( n41195 ) ;
assign n41197 =  ( n144 ) ? ( n2957 ) : ( n41196 ) ;
assign n41198 =  ( n142 ) ? ( n2956 ) : ( n41197 ) ;
assign n41199 =  ( n10 ) ? ( n2955 ) : ( n41198 ) ;
assign n41200 =  ( n3032 ) ? ( VREG_21_0 ) : ( n41194 ) ;
assign n41201 =  ( n3032 ) ? ( VREG_21_0 ) : ( n41199 ) ;
assign n41202 =  ( n3034 ) ? ( n41201 ) : ( VREG_21_0 ) ;
assign n41203 =  ( n2965 ) ? ( n41200 ) : ( n41202 ) ;
assign n41204 =  ( n1930 ) ? ( n41199 ) : ( n41203 ) ;
assign n41205 =  ( n879 ) ? ( n41194 ) : ( n41204 ) ;
assign n41206 =  ( n172 ) ? ( n3045 ) : ( VREG_21_0 ) ;
assign n41207 =  ( n170 ) ? ( n3044 ) : ( n41206 ) ;
assign n41208 =  ( n168 ) ? ( n3043 ) : ( n41207 ) ;
assign n41209 =  ( n166 ) ? ( n3042 ) : ( n41208 ) ;
assign n41210 =  ( n162 ) ? ( n3041 ) : ( n41209 ) ;
assign n41211 =  ( n172 ) ? ( n3056 ) : ( VREG_21_0 ) ;
assign n41212 =  ( n170 ) ? ( n3055 ) : ( n41211 ) ;
assign n41213 =  ( n168 ) ? ( n3054 ) : ( n41212 ) ;
assign n41214 =  ( n166 ) ? ( n3053 ) : ( n41213 ) ;
assign n41215 =  ( n162 ) ? ( n3052 ) : ( n41214 ) ;
assign n41216 =  ( n3032 ) ? ( VREG_21_0 ) : ( n41215 ) ;
assign n41217 =  ( n3051 ) ? ( n41216 ) : ( VREG_21_0 ) ;
assign n41218 =  ( n3040 ) ? ( n41210 ) : ( n41217 ) ;
assign n41219 =  ( n192 ) ? ( VREG_21_0 ) : ( VREG_21_0 ) ;
assign n41220 =  ( n157 ) ? ( n41218 ) : ( n41219 ) ;
assign n41221 =  ( n6 ) ? ( n41205 ) : ( n41220 ) ;
assign n41222 =  ( n483 ) ? ( n41221 ) : ( VREG_21_0 ) ;
assign n41223 =  ( n148 ) ? ( n4113 ) : ( VREG_21_1 ) ;
assign n41224 =  ( n146 ) ? ( n4112 ) : ( n41223 ) ;
assign n41225 =  ( n144 ) ? ( n4111 ) : ( n41224 ) ;
assign n41226 =  ( n142 ) ? ( n4110 ) : ( n41225 ) ;
assign n41227 =  ( n10 ) ? ( n4109 ) : ( n41226 ) ;
assign n41228 =  ( n148 ) ? ( n5147 ) : ( VREG_21_1 ) ;
assign n41229 =  ( n146 ) ? ( n5146 ) : ( n41228 ) ;
assign n41230 =  ( n144 ) ? ( n5145 ) : ( n41229 ) ;
assign n41231 =  ( n142 ) ? ( n5144 ) : ( n41230 ) ;
assign n41232 =  ( n10 ) ? ( n5143 ) : ( n41231 ) ;
assign n41233 =  ( n5154 ) ? ( VREG_21_1 ) : ( n41227 ) ;
assign n41234 =  ( n5154 ) ? ( VREG_21_1 ) : ( n41232 ) ;
assign n41235 =  ( n3034 ) ? ( n41234 ) : ( VREG_21_1 ) ;
assign n41236 =  ( n2965 ) ? ( n41233 ) : ( n41235 ) ;
assign n41237 =  ( n1930 ) ? ( n41232 ) : ( n41236 ) ;
assign n41238 =  ( n879 ) ? ( n41227 ) : ( n41237 ) ;
assign n41239 =  ( n172 ) ? ( n5165 ) : ( VREG_21_1 ) ;
assign n41240 =  ( n170 ) ? ( n5164 ) : ( n41239 ) ;
assign n41241 =  ( n168 ) ? ( n5163 ) : ( n41240 ) ;
assign n41242 =  ( n166 ) ? ( n5162 ) : ( n41241 ) ;
assign n41243 =  ( n162 ) ? ( n5161 ) : ( n41242 ) ;
assign n41244 =  ( n172 ) ? ( n5175 ) : ( VREG_21_1 ) ;
assign n41245 =  ( n170 ) ? ( n5174 ) : ( n41244 ) ;
assign n41246 =  ( n168 ) ? ( n5173 ) : ( n41245 ) ;
assign n41247 =  ( n166 ) ? ( n5172 ) : ( n41246 ) ;
assign n41248 =  ( n162 ) ? ( n5171 ) : ( n41247 ) ;
assign n41249 =  ( n5154 ) ? ( VREG_21_1 ) : ( n41248 ) ;
assign n41250 =  ( n3051 ) ? ( n41249 ) : ( VREG_21_1 ) ;
assign n41251 =  ( n3040 ) ? ( n41243 ) : ( n41250 ) ;
assign n41252 =  ( n192 ) ? ( VREG_21_1 ) : ( VREG_21_1 ) ;
assign n41253 =  ( n157 ) ? ( n41251 ) : ( n41252 ) ;
assign n41254 =  ( n6 ) ? ( n41238 ) : ( n41253 ) ;
assign n41255 =  ( n483 ) ? ( n41254 ) : ( VREG_21_1 ) ;
assign n41256 =  ( n148 ) ? ( n6232 ) : ( VREG_21_10 ) ;
assign n41257 =  ( n146 ) ? ( n6231 ) : ( n41256 ) ;
assign n41258 =  ( n144 ) ? ( n6230 ) : ( n41257 ) ;
assign n41259 =  ( n142 ) ? ( n6229 ) : ( n41258 ) ;
assign n41260 =  ( n10 ) ? ( n6228 ) : ( n41259 ) ;
assign n41261 =  ( n148 ) ? ( n7266 ) : ( VREG_21_10 ) ;
assign n41262 =  ( n146 ) ? ( n7265 ) : ( n41261 ) ;
assign n41263 =  ( n144 ) ? ( n7264 ) : ( n41262 ) ;
assign n41264 =  ( n142 ) ? ( n7263 ) : ( n41263 ) ;
assign n41265 =  ( n10 ) ? ( n7262 ) : ( n41264 ) ;
assign n41266 =  ( n7273 ) ? ( VREG_21_10 ) : ( n41260 ) ;
assign n41267 =  ( n7273 ) ? ( VREG_21_10 ) : ( n41265 ) ;
assign n41268 =  ( n3034 ) ? ( n41267 ) : ( VREG_21_10 ) ;
assign n41269 =  ( n2965 ) ? ( n41266 ) : ( n41268 ) ;
assign n41270 =  ( n1930 ) ? ( n41265 ) : ( n41269 ) ;
assign n41271 =  ( n879 ) ? ( n41260 ) : ( n41270 ) ;
assign n41272 =  ( n172 ) ? ( n7284 ) : ( VREG_21_10 ) ;
assign n41273 =  ( n170 ) ? ( n7283 ) : ( n41272 ) ;
assign n41274 =  ( n168 ) ? ( n7282 ) : ( n41273 ) ;
assign n41275 =  ( n166 ) ? ( n7281 ) : ( n41274 ) ;
assign n41276 =  ( n162 ) ? ( n7280 ) : ( n41275 ) ;
assign n41277 =  ( n172 ) ? ( n7294 ) : ( VREG_21_10 ) ;
assign n41278 =  ( n170 ) ? ( n7293 ) : ( n41277 ) ;
assign n41279 =  ( n168 ) ? ( n7292 ) : ( n41278 ) ;
assign n41280 =  ( n166 ) ? ( n7291 ) : ( n41279 ) ;
assign n41281 =  ( n162 ) ? ( n7290 ) : ( n41280 ) ;
assign n41282 =  ( n7273 ) ? ( VREG_21_10 ) : ( n41281 ) ;
assign n41283 =  ( n3051 ) ? ( n41282 ) : ( VREG_21_10 ) ;
assign n41284 =  ( n3040 ) ? ( n41276 ) : ( n41283 ) ;
assign n41285 =  ( n192 ) ? ( VREG_21_10 ) : ( VREG_21_10 ) ;
assign n41286 =  ( n157 ) ? ( n41284 ) : ( n41285 ) ;
assign n41287 =  ( n6 ) ? ( n41271 ) : ( n41286 ) ;
assign n41288 =  ( n483 ) ? ( n41287 ) : ( VREG_21_10 ) ;
assign n41289 =  ( n148 ) ? ( n8351 ) : ( VREG_21_11 ) ;
assign n41290 =  ( n146 ) ? ( n8350 ) : ( n41289 ) ;
assign n41291 =  ( n144 ) ? ( n8349 ) : ( n41290 ) ;
assign n41292 =  ( n142 ) ? ( n8348 ) : ( n41291 ) ;
assign n41293 =  ( n10 ) ? ( n8347 ) : ( n41292 ) ;
assign n41294 =  ( n148 ) ? ( n9385 ) : ( VREG_21_11 ) ;
assign n41295 =  ( n146 ) ? ( n9384 ) : ( n41294 ) ;
assign n41296 =  ( n144 ) ? ( n9383 ) : ( n41295 ) ;
assign n41297 =  ( n142 ) ? ( n9382 ) : ( n41296 ) ;
assign n41298 =  ( n10 ) ? ( n9381 ) : ( n41297 ) ;
assign n41299 =  ( n9392 ) ? ( VREG_21_11 ) : ( n41293 ) ;
assign n41300 =  ( n9392 ) ? ( VREG_21_11 ) : ( n41298 ) ;
assign n41301 =  ( n3034 ) ? ( n41300 ) : ( VREG_21_11 ) ;
assign n41302 =  ( n2965 ) ? ( n41299 ) : ( n41301 ) ;
assign n41303 =  ( n1930 ) ? ( n41298 ) : ( n41302 ) ;
assign n41304 =  ( n879 ) ? ( n41293 ) : ( n41303 ) ;
assign n41305 =  ( n172 ) ? ( n9403 ) : ( VREG_21_11 ) ;
assign n41306 =  ( n170 ) ? ( n9402 ) : ( n41305 ) ;
assign n41307 =  ( n168 ) ? ( n9401 ) : ( n41306 ) ;
assign n41308 =  ( n166 ) ? ( n9400 ) : ( n41307 ) ;
assign n41309 =  ( n162 ) ? ( n9399 ) : ( n41308 ) ;
assign n41310 =  ( n172 ) ? ( n9413 ) : ( VREG_21_11 ) ;
assign n41311 =  ( n170 ) ? ( n9412 ) : ( n41310 ) ;
assign n41312 =  ( n168 ) ? ( n9411 ) : ( n41311 ) ;
assign n41313 =  ( n166 ) ? ( n9410 ) : ( n41312 ) ;
assign n41314 =  ( n162 ) ? ( n9409 ) : ( n41313 ) ;
assign n41315 =  ( n9392 ) ? ( VREG_21_11 ) : ( n41314 ) ;
assign n41316 =  ( n3051 ) ? ( n41315 ) : ( VREG_21_11 ) ;
assign n41317 =  ( n3040 ) ? ( n41309 ) : ( n41316 ) ;
assign n41318 =  ( n192 ) ? ( VREG_21_11 ) : ( VREG_21_11 ) ;
assign n41319 =  ( n157 ) ? ( n41317 ) : ( n41318 ) ;
assign n41320 =  ( n6 ) ? ( n41304 ) : ( n41319 ) ;
assign n41321 =  ( n483 ) ? ( n41320 ) : ( VREG_21_11 ) ;
assign n41322 =  ( n148 ) ? ( n10470 ) : ( VREG_21_12 ) ;
assign n41323 =  ( n146 ) ? ( n10469 ) : ( n41322 ) ;
assign n41324 =  ( n144 ) ? ( n10468 ) : ( n41323 ) ;
assign n41325 =  ( n142 ) ? ( n10467 ) : ( n41324 ) ;
assign n41326 =  ( n10 ) ? ( n10466 ) : ( n41325 ) ;
assign n41327 =  ( n148 ) ? ( n11504 ) : ( VREG_21_12 ) ;
assign n41328 =  ( n146 ) ? ( n11503 ) : ( n41327 ) ;
assign n41329 =  ( n144 ) ? ( n11502 ) : ( n41328 ) ;
assign n41330 =  ( n142 ) ? ( n11501 ) : ( n41329 ) ;
assign n41331 =  ( n10 ) ? ( n11500 ) : ( n41330 ) ;
assign n41332 =  ( n11511 ) ? ( VREG_21_12 ) : ( n41326 ) ;
assign n41333 =  ( n11511 ) ? ( VREG_21_12 ) : ( n41331 ) ;
assign n41334 =  ( n3034 ) ? ( n41333 ) : ( VREG_21_12 ) ;
assign n41335 =  ( n2965 ) ? ( n41332 ) : ( n41334 ) ;
assign n41336 =  ( n1930 ) ? ( n41331 ) : ( n41335 ) ;
assign n41337 =  ( n879 ) ? ( n41326 ) : ( n41336 ) ;
assign n41338 =  ( n172 ) ? ( n11522 ) : ( VREG_21_12 ) ;
assign n41339 =  ( n170 ) ? ( n11521 ) : ( n41338 ) ;
assign n41340 =  ( n168 ) ? ( n11520 ) : ( n41339 ) ;
assign n41341 =  ( n166 ) ? ( n11519 ) : ( n41340 ) ;
assign n41342 =  ( n162 ) ? ( n11518 ) : ( n41341 ) ;
assign n41343 =  ( n172 ) ? ( n11532 ) : ( VREG_21_12 ) ;
assign n41344 =  ( n170 ) ? ( n11531 ) : ( n41343 ) ;
assign n41345 =  ( n168 ) ? ( n11530 ) : ( n41344 ) ;
assign n41346 =  ( n166 ) ? ( n11529 ) : ( n41345 ) ;
assign n41347 =  ( n162 ) ? ( n11528 ) : ( n41346 ) ;
assign n41348 =  ( n11511 ) ? ( VREG_21_12 ) : ( n41347 ) ;
assign n41349 =  ( n3051 ) ? ( n41348 ) : ( VREG_21_12 ) ;
assign n41350 =  ( n3040 ) ? ( n41342 ) : ( n41349 ) ;
assign n41351 =  ( n192 ) ? ( VREG_21_12 ) : ( VREG_21_12 ) ;
assign n41352 =  ( n157 ) ? ( n41350 ) : ( n41351 ) ;
assign n41353 =  ( n6 ) ? ( n41337 ) : ( n41352 ) ;
assign n41354 =  ( n483 ) ? ( n41353 ) : ( VREG_21_12 ) ;
assign n41355 =  ( n148 ) ? ( n12589 ) : ( VREG_21_13 ) ;
assign n41356 =  ( n146 ) ? ( n12588 ) : ( n41355 ) ;
assign n41357 =  ( n144 ) ? ( n12587 ) : ( n41356 ) ;
assign n41358 =  ( n142 ) ? ( n12586 ) : ( n41357 ) ;
assign n41359 =  ( n10 ) ? ( n12585 ) : ( n41358 ) ;
assign n41360 =  ( n148 ) ? ( n13623 ) : ( VREG_21_13 ) ;
assign n41361 =  ( n146 ) ? ( n13622 ) : ( n41360 ) ;
assign n41362 =  ( n144 ) ? ( n13621 ) : ( n41361 ) ;
assign n41363 =  ( n142 ) ? ( n13620 ) : ( n41362 ) ;
assign n41364 =  ( n10 ) ? ( n13619 ) : ( n41363 ) ;
assign n41365 =  ( n13630 ) ? ( VREG_21_13 ) : ( n41359 ) ;
assign n41366 =  ( n13630 ) ? ( VREG_21_13 ) : ( n41364 ) ;
assign n41367 =  ( n3034 ) ? ( n41366 ) : ( VREG_21_13 ) ;
assign n41368 =  ( n2965 ) ? ( n41365 ) : ( n41367 ) ;
assign n41369 =  ( n1930 ) ? ( n41364 ) : ( n41368 ) ;
assign n41370 =  ( n879 ) ? ( n41359 ) : ( n41369 ) ;
assign n41371 =  ( n172 ) ? ( n13641 ) : ( VREG_21_13 ) ;
assign n41372 =  ( n170 ) ? ( n13640 ) : ( n41371 ) ;
assign n41373 =  ( n168 ) ? ( n13639 ) : ( n41372 ) ;
assign n41374 =  ( n166 ) ? ( n13638 ) : ( n41373 ) ;
assign n41375 =  ( n162 ) ? ( n13637 ) : ( n41374 ) ;
assign n41376 =  ( n172 ) ? ( n13651 ) : ( VREG_21_13 ) ;
assign n41377 =  ( n170 ) ? ( n13650 ) : ( n41376 ) ;
assign n41378 =  ( n168 ) ? ( n13649 ) : ( n41377 ) ;
assign n41379 =  ( n166 ) ? ( n13648 ) : ( n41378 ) ;
assign n41380 =  ( n162 ) ? ( n13647 ) : ( n41379 ) ;
assign n41381 =  ( n13630 ) ? ( VREG_21_13 ) : ( n41380 ) ;
assign n41382 =  ( n3051 ) ? ( n41381 ) : ( VREG_21_13 ) ;
assign n41383 =  ( n3040 ) ? ( n41375 ) : ( n41382 ) ;
assign n41384 =  ( n192 ) ? ( VREG_21_13 ) : ( VREG_21_13 ) ;
assign n41385 =  ( n157 ) ? ( n41383 ) : ( n41384 ) ;
assign n41386 =  ( n6 ) ? ( n41370 ) : ( n41385 ) ;
assign n41387 =  ( n483 ) ? ( n41386 ) : ( VREG_21_13 ) ;
assign n41388 =  ( n148 ) ? ( n14708 ) : ( VREG_21_14 ) ;
assign n41389 =  ( n146 ) ? ( n14707 ) : ( n41388 ) ;
assign n41390 =  ( n144 ) ? ( n14706 ) : ( n41389 ) ;
assign n41391 =  ( n142 ) ? ( n14705 ) : ( n41390 ) ;
assign n41392 =  ( n10 ) ? ( n14704 ) : ( n41391 ) ;
assign n41393 =  ( n148 ) ? ( n15742 ) : ( VREG_21_14 ) ;
assign n41394 =  ( n146 ) ? ( n15741 ) : ( n41393 ) ;
assign n41395 =  ( n144 ) ? ( n15740 ) : ( n41394 ) ;
assign n41396 =  ( n142 ) ? ( n15739 ) : ( n41395 ) ;
assign n41397 =  ( n10 ) ? ( n15738 ) : ( n41396 ) ;
assign n41398 =  ( n15749 ) ? ( VREG_21_14 ) : ( n41392 ) ;
assign n41399 =  ( n15749 ) ? ( VREG_21_14 ) : ( n41397 ) ;
assign n41400 =  ( n3034 ) ? ( n41399 ) : ( VREG_21_14 ) ;
assign n41401 =  ( n2965 ) ? ( n41398 ) : ( n41400 ) ;
assign n41402 =  ( n1930 ) ? ( n41397 ) : ( n41401 ) ;
assign n41403 =  ( n879 ) ? ( n41392 ) : ( n41402 ) ;
assign n41404 =  ( n172 ) ? ( n15760 ) : ( VREG_21_14 ) ;
assign n41405 =  ( n170 ) ? ( n15759 ) : ( n41404 ) ;
assign n41406 =  ( n168 ) ? ( n15758 ) : ( n41405 ) ;
assign n41407 =  ( n166 ) ? ( n15757 ) : ( n41406 ) ;
assign n41408 =  ( n162 ) ? ( n15756 ) : ( n41407 ) ;
assign n41409 =  ( n172 ) ? ( n15770 ) : ( VREG_21_14 ) ;
assign n41410 =  ( n170 ) ? ( n15769 ) : ( n41409 ) ;
assign n41411 =  ( n168 ) ? ( n15768 ) : ( n41410 ) ;
assign n41412 =  ( n166 ) ? ( n15767 ) : ( n41411 ) ;
assign n41413 =  ( n162 ) ? ( n15766 ) : ( n41412 ) ;
assign n41414 =  ( n15749 ) ? ( VREG_21_14 ) : ( n41413 ) ;
assign n41415 =  ( n3051 ) ? ( n41414 ) : ( VREG_21_14 ) ;
assign n41416 =  ( n3040 ) ? ( n41408 ) : ( n41415 ) ;
assign n41417 =  ( n192 ) ? ( VREG_21_14 ) : ( VREG_21_14 ) ;
assign n41418 =  ( n157 ) ? ( n41416 ) : ( n41417 ) ;
assign n41419 =  ( n6 ) ? ( n41403 ) : ( n41418 ) ;
assign n41420 =  ( n483 ) ? ( n41419 ) : ( VREG_21_14 ) ;
assign n41421 =  ( n148 ) ? ( n16827 ) : ( VREG_21_15 ) ;
assign n41422 =  ( n146 ) ? ( n16826 ) : ( n41421 ) ;
assign n41423 =  ( n144 ) ? ( n16825 ) : ( n41422 ) ;
assign n41424 =  ( n142 ) ? ( n16824 ) : ( n41423 ) ;
assign n41425 =  ( n10 ) ? ( n16823 ) : ( n41424 ) ;
assign n41426 =  ( n148 ) ? ( n17861 ) : ( VREG_21_15 ) ;
assign n41427 =  ( n146 ) ? ( n17860 ) : ( n41426 ) ;
assign n41428 =  ( n144 ) ? ( n17859 ) : ( n41427 ) ;
assign n41429 =  ( n142 ) ? ( n17858 ) : ( n41428 ) ;
assign n41430 =  ( n10 ) ? ( n17857 ) : ( n41429 ) ;
assign n41431 =  ( n17868 ) ? ( VREG_21_15 ) : ( n41425 ) ;
assign n41432 =  ( n17868 ) ? ( VREG_21_15 ) : ( n41430 ) ;
assign n41433 =  ( n3034 ) ? ( n41432 ) : ( VREG_21_15 ) ;
assign n41434 =  ( n2965 ) ? ( n41431 ) : ( n41433 ) ;
assign n41435 =  ( n1930 ) ? ( n41430 ) : ( n41434 ) ;
assign n41436 =  ( n879 ) ? ( n41425 ) : ( n41435 ) ;
assign n41437 =  ( n172 ) ? ( n17879 ) : ( VREG_21_15 ) ;
assign n41438 =  ( n170 ) ? ( n17878 ) : ( n41437 ) ;
assign n41439 =  ( n168 ) ? ( n17877 ) : ( n41438 ) ;
assign n41440 =  ( n166 ) ? ( n17876 ) : ( n41439 ) ;
assign n41441 =  ( n162 ) ? ( n17875 ) : ( n41440 ) ;
assign n41442 =  ( n172 ) ? ( n17889 ) : ( VREG_21_15 ) ;
assign n41443 =  ( n170 ) ? ( n17888 ) : ( n41442 ) ;
assign n41444 =  ( n168 ) ? ( n17887 ) : ( n41443 ) ;
assign n41445 =  ( n166 ) ? ( n17886 ) : ( n41444 ) ;
assign n41446 =  ( n162 ) ? ( n17885 ) : ( n41445 ) ;
assign n41447 =  ( n17868 ) ? ( VREG_21_15 ) : ( n41446 ) ;
assign n41448 =  ( n3051 ) ? ( n41447 ) : ( VREG_21_15 ) ;
assign n41449 =  ( n3040 ) ? ( n41441 ) : ( n41448 ) ;
assign n41450 =  ( n192 ) ? ( VREG_21_15 ) : ( VREG_21_15 ) ;
assign n41451 =  ( n157 ) ? ( n41449 ) : ( n41450 ) ;
assign n41452 =  ( n6 ) ? ( n41436 ) : ( n41451 ) ;
assign n41453 =  ( n483 ) ? ( n41452 ) : ( VREG_21_15 ) ;
assign n41454 =  ( n148 ) ? ( n18946 ) : ( VREG_21_2 ) ;
assign n41455 =  ( n146 ) ? ( n18945 ) : ( n41454 ) ;
assign n41456 =  ( n144 ) ? ( n18944 ) : ( n41455 ) ;
assign n41457 =  ( n142 ) ? ( n18943 ) : ( n41456 ) ;
assign n41458 =  ( n10 ) ? ( n18942 ) : ( n41457 ) ;
assign n41459 =  ( n148 ) ? ( n19980 ) : ( VREG_21_2 ) ;
assign n41460 =  ( n146 ) ? ( n19979 ) : ( n41459 ) ;
assign n41461 =  ( n144 ) ? ( n19978 ) : ( n41460 ) ;
assign n41462 =  ( n142 ) ? ( n19977 ) : ( n41461 ) ;
assign n41463 =  ( n10 ) ? ( n19976 ) : ( n41462 ) ;
assign n41464 =  ( n19987 ) ? ( VREG_21_2 ) : ( n41458 ) ;
assign n41465 =  ( n19987 ) ? ( VREG_21_2 ) : ( n41463 ) ;
assign n41466 =  ( n3034 ) ? ( n41465 ) : ( VREG_21_2 ) ;
assign n41467 =  ( n2965 ) ? ( n41464 ) : ( n41466 ) ;
assign n41468 =  ( n1930 ) ? ( n41463 ) : ( n41467 ) ;
assign n41469 =  ( n879 ) ? ( n41458 ) : ( n41468 ) ;
assign n41470 =  ( n172 ) ? ( n19998 ) : ( VREG_21_2 ) ;
assign n41471 =  ( n170 ) ? ( n19997 ) : ( n41470 ) ;
assign n41472 =  ( n168 ) ? ( n19996 ) : ( n41471 ) ;
assign n41473 =  ( n166 ) ? ( n19995 ) : ( n41472 ) ;
assign n41474 =  ( n162 ) ? ( n19994 ) : ( n41473 ) ;
assign n41475 =  ( n172 ) ? ( n20008 ) : ( VREG_21_2 ) ;
assign n41476 =  ( n170 ) ? ( n20007 ) : ( n41475 ) ;
assign n41477 =  ( n168 ) ? ( n20006 ) : ( n41476 ) ;
assign n41478 =  ( n166 ) ? ( n20005 ) : ( n41477 ) ;
assign n41479 =  ( n162 ) ? ( n20004 ) : ( n41478 ) ;
assign n41480 =  ( n19987 ) ? ( VREG_21_2 ) : ( n41479 ) ;
assign n41481 =  ( n3051 ) ? ( n41480 ) : ( VREG_21_2 ) ;
assign n41482 =  ( n3040 ) ? ( n41474 ) : ( n41481 ) ;
assign n41483 =  ( n192 ) ? ( VREG_21_2 ) : ( VREG_21_2 ) ;
assign n41484 =  ( n157 ) ? ( n41482 ) : ( n41483 ) ;
assign n41485 =  ( n6 ) ? ( n41469 ) : ( n41484 ) ;
assign n41486 =  ( n483 ) ? ( n41485 ) : ( VREG_21_2 ) ;
assign n41487 =  ( n148 ) ? ( n21065 ) : ( VREG_21_3 ) ;
assign n41488 =  ( n146 ) ? ( n21064 ) : ( n41487 ) ;
assign n41489 =  ( n144 ) ? ( n21063 ) : ( n41488 ) ;
assign n41490 =  ( n142 ) ? ( n21062 ) : ( n41489 ) ;
assign n41491 =  ( n10 ) ? ( n21061 ) : ( n41490 ) ;
assign n41492 =  ( n148 ) ? ( n22099 ) : ( VREG_21_3 ) ;
assign n41493 =  ( n146 ) ? ( n22098 ) : ( n41492 ) ;
assign n41494 =  ( n144 ) ? ( n22097 ) : ( n41493 ) ;
assign n41495 =  ( n142 ) ? ( n22096 ) : ( n41494 ) ;
assign n41496 =  ( n10 ) ? ( n22095 ) : ( n41495 ) ;
assign n41497 =  ( n22106 ) ? ( VREG_21_3 ) : ( n41491 ) ;
assign n41498 =  ( n22106 ) ? ( VREG_21_3 ) : ( n41496 ) ;
assign n41499 =  ( n3034 ) ? ( n41498 ) : ( VREG_21_3 ) ;
assign n41500 =  ( n2965 ) ? ( n41497 ) : ( n41499 ) ;
assign n41501 =  ( n1930 ) ? ( n41496 ) : ( n41500 ) ;
assign n41502 =  ( n879 ) ? ( n41491 ) : ( n41501 ) ;
assign n41503 =  ( n172 ) ? ( n22117 ) : ( VREG_21_3 ) ;
assign n41504 =  ( n170 ) ? ( n22116 ) : ( n41503 ) ;
assign n41505 =  ( n168 ) ? ( n22115 ) : ( n41504 ) ;
assign n41506 =  ( n166 ) ? ( n22114 ) : ( n41505 ) ;
assign n41507 =  ( n162 ) ? ( n22113 ) : ( n41506 ) ;
assign n41508 =  ( n172 ) ? ( n22127 ) : ( VREG_21_3 ) ;
assign n41509 =  ( n170 ) ? ( n22126 ) : ( n41508 ) ;
assign n41510 =  ( n168 ) ? ( n22125 ) : ( n41509 ) ;
assign n41511 =  ( n166 ) ? ( n22124 ) : ( n41510 ) ;
assign n41512 =  ( n162 ) ? ( n22123 ) : ( n41511 ) ;
assign n41513 =  ( n22106 ) ? ( VREG_21_3 ) : ( n41512 ) ;
assign n41514 =  ( n3051 ) ? ( n41513 ) : ( VREG_21_3 ) ;
assign n41515 =  ( n3040 ) ? ( n41507 ) : ( n41514 ) ;
assign n41516 =  ( n192 ) ? ( VREG_21_3 ) : ( VREG_21_3 ) ;
assign n41517 =  ( n157 ) ? ( n41515 ) : ( n41516 ) ;
assign n41518 =  ( n6 ) ? ( n41502 ) : ( n41517 ) ;
assign n41519 =  ( n483 ) ? ( n41518 ) : ( VREG_21_3 ) ;
assign n41520 =  ( n148 ) ? ( n23184 ) : ( VREG_21_4 ) ;
assign n41521 =  ( n146 ) ? ( n23183 ) : ( n41520 ) ;
assign n41522 =  ( n144 ) ? ( n23182 ) : ( n41521 ) ;
assign n41523 =  ( n142 ) ? ( n23181 ) : ( n41522 ) ;
assign n41524 =  ( n10 ) ? ( n23180 ) : ( n41523 ) ;
assign n41525 =  ( n148 ) ? ( n24218 ) : ( VREG_21_4 ) ;
assign n41526 =  ( n146 ) ? ( n24217 ) : ( n41525 ) ;
assign n41527 =  ( n144 ) ? ( n24216 ) : ( n41526 ) ;
assign n41528 =  ( n142 ) ? ( n24215 ) : ( n41527 ) ;
assign n41529 =  ( n10 ) ? ( n24214 ) : ( n41528 ) ;
assign n41530 =  ( n24225 ) ? ( VREG_21_4 ) : ( n41524 ) ;
assign n41531 =  ( n24225 ) ? ( VREG_21_4 ) : ( n41529 ) ;
assign n41532 =  ( n3034 ) ? ( n41531 ) : ( VREG_21_4 ) ;
assign n41533 =  ( n2965 ) ? ( n41530 ) : ( n41532 ) ;
assign n41534 =  ( n1930 ) ? ( n41529 ) : ( n41533 ) ;
assign n41535 =  ( n879 ) ? ( n41524 ) : ( n41534 ) ;
assign n41536 =  ( n172 ) ? ( n24236 ) : ( VREG_21_4 ) ;
assign n41537 =  ( n170 ) ? ( n24235 ) : ( n41536 ) ;
assign n41538 =  ( n168 ) ? ( n24234 ) : ( n41537 ) ;
assign n41539 =  ( n166 ) ? ( n24233 ) : ( n41538 ) ;
assign n41540 =  ( n162 ) ? ( n24232 ) : ( n41539 ) ;
assign n41541 =  ( n172 ) ? ( n24246 ) : ( VREG_21_4 ) ;
assign n41542 =  ( n170 ) ? ( n24245 ) : ( n41541 ) ;
assign n41543 =  ( n168 ) ? ( n24244 ) : ( n41542 ) ;
assign n41544 =  ( n166 ) ? ( n24243 ) : ( n41543 ) ;
assign n41545 =  ( n162 ) ? ( n24242 ) : ( n41544 ) ;
assign n41546 =  ( n24225 ) ? ( VREG_21_4 ) : ( n41545 ) ;
assign n41547 =  ( n3051 ) ? ( n41546 ) : ( VREG_21_4 ) ;
assign n41548 =  ( n3040 ) ? ( n41540 ) : ( n41547 ) ;
assign n41549 =  ( n192 ) ? ( VREG_21_4 ) : ( VREG_21_4 ) ;
assign n41550 =  ( n157 ) ? ( n41548 ) : ( n41549 ) ;
assign n41551 =  ( n6 ) ? ( n41535 ) : ( n41550 ) ;
assign n41552 =  ( n483 ) ? ( n41551 ) : ( VREG_21_4 ) ;
assign n41553 =  ( n148 ) ? ( n25303 ) : ( VREG_21_5 ) ;
assign n41554 =  ( n146 ) ? ( n25302 ) : ( n41553 ) ;
assign n41555 =  ( n144 ) ? ( n25301 ) : ( n41554 ) ;
assign n41556 =  ( n142 ) ? ( n25300 ) : ( n41555 ) ;
assign n41557 =  ( n10 ) ? ( n25299 ) : ( n41556 ) ;
assign n41558 =  ( n148 ) ? ( n26337 ) : ( VREG_21_5 ) ;
assign n41559 =  ( n146 ) ? ( n26336 ) : ( n41558 ) ;
assign n41560 =  ( n144 ) ? ( n26335 ) : ( n41559 ) ;
assign n41561 =  ( n142 ) ? ( n26334 ) : ( n41560 ) ;
assign n41562 =  ( n10 ) ? ( n26333 ) : ( n41561 ) ;
assign n41563 =  ( n26344 ) ? ( VREG_21_5 ) : ( n41557 ) ;
assign n41564 =  ( n26344 ) ? ( VREG_21_5 ) : ( n41562 ) ;
assign n41565 =  ( n3034 ) ? ( n41564 ) : ( VREG_21_5 ) ;
assign n41566 =  ( n2965 ) ? ( n41563 ) : ( n41565 ) ;
assign n41567 =  ( n1930 ) ? ( n41562 ) : ( n41566 ) ;
assign n41568 =  ( n879 ) ? ( n41557 ) : ( n41567 ) ;
assign n41569 =  ( n172 ) ? ( n26355 ) : ( VREG_21_5 ) ;
assign n41570 =  ( n170 ) ? ( n26354 ) : ( n41569 ) ;
assign n41571 =  ( n168 ) ? ( n26353 ) : ( n41570 ) ;
assign n41572 =  ( n166 ) ? ( n26352 ) : ( n41571 ) ;
assign n41573 =  ( n162 ) ? ( n26351 ) : ( n41572 ) ;
assign n41574 =  ( n172 ) ? ( n26365 ) : ( VREG_21_5 ) ;
assign n41575 =  ( n170 ) ? ( n26364 ) : ( n41574 ) ;
assign n41576 =  ( n168 ) ? ( n26363 ) : ( n41575 ) ;
assign n41577 =  ( n166 ) ? ( n26362 ) : ( n41576 ) ;
assign n41578 =  ( n162 ) ? ( n26361 ) : ( n41577 ) ;
assign n41579 =  ( n26344 ) ? ( VREG_21_5 ) : ( n41578 ) ;
assign n41580 =  ( n3051 ) ? ( n41579 ) : ( VREG_21_5 ) ;
assign n41581 =  ( n3040 ) ? ( n41573 ) : ( n41580 ) ;
assign n41582 =  ( n192 ) ? ( VREG_21_5 ) : ( VREG_21_5 ) ;
assign n41583 =  ( n157 ) ? ( n41581 ) : ( n41582 ) ;
assign n41584 =  ( n6 ) ? ( n41568 ) : ( n41583 ) ;
assign n41585 =  ( n483 ) ? ( n41584 ) : ( VREG_21_5 ) ;
assign n41586 =  ( n148 ) ? ( n27422 ) : ( VREG_21_6 ) ;
assign n41587 =  ( n146 ) ? ( n27421 ) : ( n41586 ) ;
assign n41588 =  ( n144 ) ? ( n27420 ) : ( n41587 ) ;
assign n41589 =  ( n142 ) ? ( n27419 ) : ( n41588 ) ;
assign n41590 =  ( n10 ) ? ( n27418 ) : ( n41589 ) ;
assign n41591 =  ( n148 ) ? ( n28456 ) : ( VREG_21_6 ) ;
assign n41592 =  ( n146 ) ? ( n28455 ) : ( n41591 ) ;
assign n41593 =  ( n144 ) ? ( n28454 ) : ( n41592 ) ;
assign n41594 =  ( n142 ) ? ( n28453 ) : ( n41593 ) ;
assign n41595 =  ( n10 ) ? ( n28452 ) : ( n41594 ) ;
assign n41596 =  ( n28463 ) ? ( VREG_21_6 ) : ( n41590 ) ;
assign n41597 =  ( n28463 ) ? ( VREG_21_6 ) : ( n41595 ) ;
assign n41598 =  ( n3034 ) ? ( n41597 ) : ( VREG_21_6 ) ;
assign n41599 =  ( n2965 ) ? ( n41596 ) : ( n41598 ) ;
assign n41600 =  ( n1930 ) ? ( n41595 ) : ( n41599 ) ;
assign n41601 =  ( n879 ) ? ( n41590 ) : ( n41600 ) ;
assign n41602 =  ( n172 ) ? ( n28474 ) : ( VREG_21_6 ) ;
assign n41603 =  ( n170 ) ? ( n28473 ) : ( n41602 ) ;
assign n41604 =  ( n168 ) ? ( n28472 ) : ( n41603 ) ;
assign n41605 =  ( n166 ) ? ( n28471 ) : ( n41604 ) ;
assign n41606 =  ( n162 ) ? ( n28470 ) : ( n41605 ) ;
assign n41607 =  ( n172 ) ? ( n28484 ) : ( VREG_21_6 ) ;
assign n41608 =  ( n170 ) ? ( n28483 ) : ( n41607 ) ;
assign n41609 =  ( n168 ) ? ( n28482 ) : ( n41608 ) ;
assign n41610 =  ( n166 ) ? ( n28481 ) : ( n41609 ) ;
assign n41611 =  ( n162 ) ? ( n28480 ) : ( n41610 ) ;
assign n41612 =  ( n28463 ) ? ( VREG_21_6 ) : ( n41611 ) ;
assign n41613 =  ( n3051 ) ? ( n41612 ) : ( VREG_21_6 ) ;
assign n41614 =  ( n3040 ) ? ( n41606 ) : ( n41613 ) ;
assign n41615 =  ( n192 ) ? ( VREG_21_6 ) : ( VREG_21_6 ) ;
assign n41616 =  ( n157 ) ? ( n41614 ) : ( n41615 ) ;
assign n41617 =  ( n6 ) ? ( n41601 ) : ( n41616 ) ;
assign n41618 =  ( n483 ) ? ( n41617 ) : ( VREG_21_6 ) ;
assign n41619 =  ( n148 ) ? ( n29541 ) : ( VREG_21_7 ) ;
assign n41620 =  ( n146 ) ? ( n29540 ) : ( n41619 ) ;
assign n41621 =  ( n144 ) ? ( n29539 ) : ( n41620 ) ;
assign n41622 =  ( n142 ) ? ( n29538 ) : ( n41621 ) ;
assign n41623 =  ( n10 ) ? ( n29537 ) : ( n41622 ) ;
assign n41624 =  ( n148 ) ? ( n30575 ) : ( VREG_21_7 ) ;
assign n41625 =  ( n146 ) ? ( n30574 ) : ( n41624 ) ;
assign n41626 =  ( n144 ) ? ( n30573 ) : ( n41625 ) ;
assign n41627 =  ( n142 ) ? ( n30572 ) : ( n41626 ) ;
assign n41628 =  ( n10 ) ? ( n30571 ) : ( n41627 ) ;
assign n41629 =  ( n30582 ) ? ( VREG_21_7 ) : ( n41623 ) ;
assign n41630 =  ( n30582 ) ? ( VREG_21_7 ) : ( n41628 ) ;
assign n41631 =  ( n3034 ) ? ( n41630 ) : ( VREG_21_7 ) ;
assign n41632 =  ( n2965 ) ? ( n41629 ) : ( n41631 ) ;
assign n41633 =  ( n1930 ) ? ( n41628 ) : ( n41632 ) ;
assign n41634 =  ( n879 ) ? ( n41623 ) : ( n41633 ) ;
assign n41635 =  ( n172 ) ? ( n30593 ) : ( VREG_21_7 ) ;
assign n41636 =  ( n170 ) ? ( n30592 ) : ( n41635 ) ;
assign n41637 =  ( n168 ) ? ( n30591 ) : ( n41636 ) ;
assign n41638 =  ( n166 ) ? ( n30590 ) : ( n41637 ) ;
assign n41639 =  ( n162 ) ? ( n30589 ) : ( n41638 ) ;
assign n41640 =  ( n172 ) ? ( n30603 ) : ( VREG_21_7 ) ;
assign n41641 =  ( n170 ) ? ( n30602 ) : ( n41640 ) ;
assign n41642 =  ( n168 ) ? ( n30601 ) : ( n41641 ) ;
assign n41643 =  ( n166 ) ? ( n30600 ) : ( n41642 ) ;
assign n41644 =  ( n162 ) ? ( n30599 ) : ( n41643 ) ;
assign n41645 =  ( n30582 ) ? ( VREG_21_7 ) : ( n41644 ) ;
assign n41646 =  ( n3051 ) ? ( n41645 ) : ( VREG_21_7 ) ;
assign n41647 =  ( n3040 ) ? ( n41639 ) : ( n41646 ) ;
assign n41648 =  ( n192 ) ? ( VREG_21_7 ) : ( VREG_21_7 ) ;
assign n41649 =  ( n157 ) ? ( n41647 ) : ( n41648 ) ;
assign n41650 =  ( n6 ) ? ( n41634 ) : ( n41649 ) ;
assign n41651 =  ( n483 ) ? ( n41650 ) : ( VREG_21_7 ) ;
assign n41652 =  ( n148 ) ? ( n31660 ) : ( VREG_21_8 ) ;
assign n41653 =  ( n146 ) ? ( n31659 ) : ( n41652 ) ;
assign n41654 =  ( n144 ) ? ( n31658 ) : ( n41653 ) ;
assign n41655 =  ( n142 ) ? ( n31657 ) : ( n41654 ) ;
assign n41656 =  ( n10 ) ? ( n31656 ) : ( n41655 ) ;
assign n41657 =  ( n148 ) ? ( n32694 ) : ( VREG_21_8 ) ;
assign n41658 =  ( n146 ) ? ( n32693 ) : ( n41657 ) ;
assign n41659 =  ( n144 ) ? ( n32692 ) : ( n41658 ) ;
assign n41660 =  ( n142 ) ? ( n32691 ) : ( n41659 ) ;
assign n41661 =  ( n10 ) ? ( n32690 ) : ( n41660 ) ;
assign n41662 =  ( n32701 ) ? ( VREG_21_8 ) : ( n41656 ) ;
assign n41663 =  ( n32701 ) ? ( VREG_21_8 ) : ( n41661 ) ;
assign n41664 =  ( n3034 ) ? ( n41663 ) : ( VREG_21_8 ) ;
assign n41665 =  ( n2965 ) ? ( n41662 ) : ( n41664 ) ;
assign n41666 =  ( n1930 ) ? ( n41661 ) : ( n41665 ) ;
assign n41667 =  ( n879 ) ? ( n41656 ) : ( n41666 ) ;
assign n41668 =  ( n172 ) ? ( n32712 ) : ( VREG_21_8 ) ;
assign n41669 =  ( n170 ) ? ( n32711 ) : ( n41668 ) ;
assign n41670 =  ( n168 ) ? ( n32710 ) : ( n41669 ) ;
assign n41671 =  ( n166 ) ? ( n32709 ) : ( n41670 ) ;
assign n41672 =  ( n162 ) ? ( n32708 ) : ( n41671 ) ;
assign n41673 =  ( n172 ) ? ( n32722 ) : ( VREG_21_8 ) ;
assign n41674 =  ( n170 ) ? ( n32721 ) : ( n41673 ) ;
assign n41675 =  ( n168 ) ? ( n32720 ) : ( n41674 ) ;
assign n41676 =  ( n166 ) ? ( n32719 ) : ( n41675 ) ;
assign n41677 =  ( n162 ) ? ( n32718 ) : ( n41676 ) ;
assign n41678 =  ( n32701 ) ? ( VREG_21_8 ) : ( n41677 ) ;
assign n41679 =  ( n3051 ) ? ( n41678 ) : ( VREG_21_8 ) ;
assign n41680 =  ( n3040 ) ? ( n41672 ) : ( n41679 ) ;
assign n41681 =  ( n192 ) ? ( VREG_21_8 ) : ( VREG_21_8 ) ;
assign n41682 =  ( n157 ) ? ( n41680 ) : ( n41681 ) ;
assign n41683 =  ( n6 ) ? ( n41667 ) : ( n41682 ) ;
assign n41684 =  ( n483 ) ? ( n41683 ) : ( VREG_21_8 ) ;
assign n41685 =  ( n148 ) ? ( n33779 ) : ( VREG_21_9 ) ;
assign n41686 =  ( n146 ) ? ( n33778 ) : ( n41685 ) ;
assign n41687 =  ( n144 ) ? ( n33777 ) : ( n41686 ) ;
assign n41688 =  ( n142 ) ? ( n33776 ) : ( n41687 ) ;
assign n41689 =  ( n10 ) ? ( n33775 ) : ( n41688 ) ;
assign n41690 =  ( n148 ) ? ( n34813 ) : ( VREG_21_9 ) ;
assign n41691 =  ( n146 ) ? ( n34812 ) : ( n41690 ) ;
assign n41692 =  ( n144 ) ? ( n34811 ) : ( n41691 ) ;
assign n41693 =  ( n142 ) ? ( n34810 ) : ( n41692 ) ;
assign n41694 =  ( n10 ) ? ( n34809 ) : ( n41693 ) ;
assign n41695 =  ( n34820 ) ? ( VREG_21_9 ) : ( n41689 ) ;
assign n41696 =  ( n34820 ) ? ( VREG_21_9 ) : ( n41694 ) ;
assign n41697 =  ( n3034 ) ? ( n41696 ) : ( VREG_21_9 ) ;
assign n41698 =  ( n2965 ) ? ( n41695 ) : ( n41697 ) ;
assign n41699 =  ( n1930 ) ? ( n41694 ) : ( n41698 ) ;
assign n41700 =  ( n879 ) ? ( n41689 ) : ( n41699 ) ;
assign n41701 =  ( n172 ) ? ( n34831 ) : ( VREG_21_9 ) ;
assign n41702 =  ( n170 ) ? ( n34830 ) : ( n41701 ) ;
assign n41703 =  ( n168 ) ? ( n34829 ) : ( n41702 ) ;
assign n41704 =  ( n166 ) ? ( n34828 ) : ( n41703 ) ;
assign n41705 =  ( n162 ) ? ( n34827 ) : ( n41704 ) ;
assign n41706 =  ( n172 ) ? ( n34841 ) : ( VREG_21_9 ) ;
assign n41707 =  ( n170 ) ? ( n34840 ) : ( n41706 ) ;
assign n41708 =  ( n168 ) ? ( n34839 ) : ( n41707 ) ;
assign n41709 =  ( n166 ) ? ( n34838 ) : ( n41708 ) ;
assign n41710 =  ( n162 ) ? ( n34837 ) : ( n41709 ) ;
assign n41711 =  ( n34820 ) ? ( VREG_21_9 ) : ( n41710 ) ;
assign n41712 =  ( n3051 ) ? ( n41711 ) : ( VREG_21_9 ) ;
assign n41713 =  ( n3040 ) ? ( n41705 ) : ( n41712 ) ;
assign n41714 =  ( n192 ) ? ( VREG_21_9 ) : ( VREG_21_9 ) ;
assign n41715 =  ( n157 ) ? ( n41713 ) : ( n41714 ) ;
assign n41716 =  ( n6 ) ? ( n41700 ) : ( n41715 ) ;
assign n41717 =  ( n483 ) ? ( n41716 ) : ( VREG_21_9 ) ;
assign n41718 =  ( n148 ) ? ( n1924 ) : ( VREG_22_0 ) ;
assign n41719 =  ( n146 ) ? ( n1923 ) : ( n41718 ) ;
assign n41720 =  ( n144 ) ? ( n1922 ) : ( n41719 ) ;
assign n41721 =  ( n142 ) ? ( n1921 ) : ( n41720 ) ;
assign n41722 =  ( n10 ) ? ( n1920 ) : ( n41721 ) ;
assign n41723 =  ( n148 ) ? ( n2959 ) : ( VREG_22_0 ) ;
assign n41724 =  ( n146 ) ? ( n2958 ) : ( n41723 ) ;
assign n41725 =  ( n144 ) ? ( n2957 ) : ( n41724 ) ;
assign n41726 =  ( n142 ) ? ( n2956 ) : ( n41725 ) ;
assign n41727 =  ( n10 ) ? ( n2955 ) : ( n41726 ) ;
assign n41728 =  ( n3032 ) ? ( VREG_22_0 ) : ( n41722 ) ;
assign n41729 =  ( n3032 ) ? ( VREG_22_0 ) : ( n41727 ) ;
assign n41730 =  ( n3034 ) ? ( n41729 ) : ( VREG_22_0 ) ;
assign n41731 =  ( n2965 ) ? ( n41728 ) : ( n41730 ) ;
assign n41732 =  ( n1930 ) ? ( n41727 ) : ( n41731 ) ;
assign n41733 =  ( n879 ) ? ( n41722 ) : ( n41732 ) ;
assign n41734 =  ( n172 ) ? ( n3045 ) : ( VREG_22_0 ) ;
assign n41735 =  ( n170 ) ? ( n3044 ) : ( n41734 ) ;
assign n41736 =  ( n168 ) ? ( n3043 ) : ( n41735 ) ;
assign n41737 =  ( n166 ) ? ( n3042 ) : ( n41736 ) ;
assign n41738 =  ( n162 ) ? ( n3041 ) : ( n41737 ) ;
assign n41739 =  ( n172 ) ? ( n3056 ) : ( VREG_22_0 ) ;
assign n41740 =  ( n170 ) ? ( n3055 ) : ( n41739 ) ;
assign n41741 =  ( n168 ) ? ( n3054 ) : ( n41740 ) ;
assign n41742 =  ( n166 ) ? ( n3053 ) : ( n41741 ) ;
assign n41743 =  ( n162 ) ? ( n3052 ) : ( n41742 ) ;
assign n41744 =  ( n3032 ) ? ( VREG_22_0 ) : ( n41743 ) ;
assign n41745 =  ( n3051 ) ? ( n41744 ) : ( VREG_22_0 ) ;
assign n41746 =  ( n3040 ) ? ( n41738 ) : ( n41745 ) ;
assign n41747 =  ( n192 ) ? ( VREG_22_0 ) : ( VREG_22_0 ) ;
assign n41748 =  ( n157 ) ? ( n41746 ) : ( n41747 ) ;
assign n41749 =  ( n6 ) ? ( n41733 ) : ( n41748 ) ;
assign n41750 =  ( n505 ) ? ( n41749 ) : ( VREG_22_0 ) ;
assign n41751 =  ( n148 ) ? ( n4113 ) : ( VREG_22_1 ) ;
assign n41752 =  ( n146 ) ? ( n4112 ) : ( n41751 ) ;
assign n41753 =  ( n144 ) ? ( n4111 ) : ( n41752 ) ;
assign n41754 =  ( n142 ) ? ( n4110 ) : ( n41753 ) ;
assign n41755 =  ( n10 ) ? ( n4109 ) : ( n41754 ) ;
assign n41756 =  ( n148 ) ? ( n5147 ) : ( VREG_22_1 ) ;
assign n41757 =  ( n146 ) ? ( n5146 ) : ( n41756 ) ;
assign n41758 =  ( n144 ) ? ( n5145 ) : ( n41757 ) ;
assign n41759 =  ( n142 ) ? ( n5144 ) : ( n41758 ) ;
assign n41760 =  ( n10 ) ? ( n5143 ) : ( n41759 ) ;
assign n41761 =  ( n5154 ) ? ( VREG_22_1 ) : ( n41755 ) ;
assign n41762 =  ( n5154 ) ? ( VREG_22_1 ) : ( n41760 ) ;
assign n41763 =  ( n3034 ) ? ( n41762 ) : ( VREG_22_1 ) ;
assign n41764 =  ( n2965 ) ? ( n41761 ) : ( n41763 ) ;
assign n41765 =  ( n1930 ) ? ( n41760 ) : ( n41764 ) ;
assign n41766 =  ( n879 ) ? ( n41755 ) : ( n41765 ) ;
assign n41767 =  ( n172 ) ? ( n5165 ) : ( VREG_22_1 ) ;
assign n41768 =  ( n170 ) ? ( n5164 ) : ( n41767 ) ;
assign n41769 =  ( n168 ) ? ( n5163 ) : ( n41768 ) ;
assign n41770 =  ( n166 ) ? ( n5162 ) : ( n41769 ) ;
assign n41771 =  ( n162 ) ? ( n5161 ) : ( n41770 ) ;
assign n41772 =  ( n172 ) ? ( n5175 ) : ( VREG_22_1 ) ;
assign n41773 =  ( n170 ) ? ( n5174 ) : ( n41772 ) ;
assign n41774 =  ( n168 ) ? ( n5173 ) : ( n41773 ) ;
assign n41775 =  ( n166 ) ? ( n5172 ) : ( n41774 ) ;
assign n41776 =  ( n162 ) ? ( n5171 ) : ( n41775 ) ;
assign n41777 =  ( n5154 ) ? ( VREG_22_1 ) : ( n41776 ) ;
assign n41778 =  ( n3051 ) ? ( n41777 ) : ( VREG_22_1 ) ;
assign n41779 =  ( n3040 ) ? ( n41771 ) : ( n41778 ) ;
assign n41780 =  ( n192 ) ? ( VREG_22_1 ) : ( VREG_22_1 ) ;
assign n41781 =  ( n157 ) ? ( n41779 ) : ( n41780 ) ;
assign n41782 =  ( n6 ) ? ( n41766 ) : ( n41781 ) ;
assign n41783 =  ( n505 ) ? ( n41782 ) : ( VREG_22_1 ) ;
assign n41784 =  ( n148 ) ? ( n6232 ) : ( VREG_22_10 ) ;
assign n41785 =  ( n146 ) ? ( n6231 ) : ( n41784 ) ;
assign n41786 =  ( n144 ) ? ( n6230 ) : ( n41785 ) ;
assign n41787 =  ( n142 ) ? ( n6229 ) : ( n41786 ) ;
assign n41788 =  ( n10 ) ? ( n6228 ) : ( n41787 ) ;
assign n41789 =  ( n148 ) ? ( n7266 ) : ( VREG_22_10 ) ;
assign n41790 =  ( n146 ) ? ( n7265 ) : ( n41789 ) ;
assign n41791 =  ( n144 ) ? ( n7264 ) : ( n41790 ) ;
assign n41792 =  ( n142 ) ? ( n7263 ) : ( n41791 ) ;
assign n41793 =  ( n10 ) ? ( n7262 ) : ( n41792 ) ;
assign n41794 =  ( n7273 ) ? ( VREG_22_10 ) : ( n41788 ) ;
assign n41795 =  ( n7273 ) ? ( VREG_22_10 ) : ( n41793 ) ;
assign n41796 =  ( n3034 ) ? ( n41795 ) : ( VREG_22_10 ) ;
assign n41797 =  ( n2965 ) ? ( n41794 ) : ( n41796 ) ;
assign n41798 =  ( n1930 ) ? ( n41793 ) : ( n41797 ) ;
assign n41799 =  ( n879 ) ? ( n41788 ) : ( n41798 ) ;
assign n41800 =  ( n172 ) ? ( n7284 ) : ( VREG_22_10 ) ;
assign n41801 =  ( n170 ) ? ( n7283 ) : ( n41800 ) ;
assign n41802 =  ( n168 ) ? ( n7282 ) : ( n41801 ) ;
assign n41803 =  ( n166 ) ? ( n7281 ) : ( n41802 ) ;
assign n41804 =  ( n162 ) ? ( n7280 ) : ( n41803 ) ;
assign n41805 =  ( n172 ) ? ( n7294 ) : ( VREG_22_10 ) ;
assign n41806 =  ( n170 ) ? ( n7293 ) : ( n41805 ) ;
assign n41807 =  ( n168 ) ? ( n7292 ) : ( n41806 ) ;
assign n41808 =  ( n166 ) ? ( n7291 ) : ( n41807 ) ;
assign n41809 =  ( n162 ) ? ( n7290 ) : ( n41808 ) ;
assign n41810 =  ( n7273 ) ? ( VREG_22_10 ) : ( n41809 ) ;
assign n41811 =  ( n3051 ) ? ( n41810 ) : ( VREG_22_10 ) ;
assign n41812 =  ( n3040 ) ? ( n41804 ) : ( n41811 ) ;
assign n41813 =  ( n192 ) ? ( VREG_22_10 ) : ( VREG_22_10 ) ;
assign n41814 =  ( n157 ) ? ( n41812 ) : ( n41813 ) ;
assign n41815 =  ( n6 ) ? ( n41799 ) : ( n41814 ) ;
assign n41816 =  ( n505 ) ? ( n41815 ) : ( VREG_22_10 ) ;
assign n41817 =  ( n148 ) ? ( n8351 ) : ( VREG_22_11 ) ;
assign n41818 =  ( n146 ) ? ( n8350 ) : ( n41817 ) ;
assign n41819 =  ( n144 ) ? ( n8349 ) : ( n41818 ) ;
assign n41820 =  ( n142 ) ? ( n8348 ) : ( n41819 ) ;
assign n41821 =  ( n10 ) ? ( n8347 ) : ( n41820 ) ;
assign n41822 =  ( n148 ) ? ( n9385 ) : ( VREG_22_11 ) ;
assign n41823 =  ( n146 ) ? ( n9384 ) : ( n41822 ) ;
assign n41824 =  ( n144 ) ? ( n9383 ) : ( n41823 ) ;
assign n41825 =  ( n142 ) ? ( n9382 ) : ( n41824 ) ;
assign n41826 =  ( n10 ) ? ( n9381 ) : ( n41825 ) ;
assign n41827 =  ( n9392 ) ? ( VREG_22_11 ) : ( n41821 ) ;
assign n41828 =  ( n9392 ) ? ( VREG_22_11 ) : ( n41826 ) ;
assign n41829 =  ( n3034 ) ? ( n41828 ) : ( VREG_22_11 ) ;
assign n41830 =  ( n2965 ) ? ( n41827 ) : ( n41829 ) ;
assign n41831 =  ( n1930 ) ? ( n41826 ) : ( n41830 ) ;
assign n41832 =  ( n879 ) ? ( n41821 ) : ( n41831 ) ;
assign n41833 =  ( n172 ) ? ( n9403 ) : ( VREG_22_11 ) ;
assign n41834 =  ( n170 ) ? ( n9402 ) : ( n41833 ) ;
assign n41835 =  ( n168 ) ? ( n9401 ) : ( n41834 ) ;
assign n41836 =  ( n166 ) ? ( n9400 ) : ( n41835 ) ;
assign n41837 =  ( n162 ) ? ( n9399 ) : ( n41836 ) ;
assign n41838 =  ( n172 ) ? ( n9413 ) : ( VREG_22_11 ) ;
assign n41839 =  ( n170 ) ? ( n9412 ) : ( n41838 ) ;
assign n41840 =  ( n168 ) ? ( n9411 ) : ( n41839 ) ;
assign n41841 =  ( n166 ) ? ( n9410 ) : ( n41840 ) ;
assign n41842 =  ( n162 ) ? ( n9409 ) : ( n41841 ) ;
assign n41843 =  ( n9392 ) ? ( VREG_22_11 ) : ( n41842 ) ;
assign n41844 =  ( n3051 ) ? ( n41843 ) : ( VREG_22_11 ) ;
assign n41845 =  ( n3040 ) ? ( n41837 ) : ( n41844 ) ;
assign n41846 =  ( n192 ) ? ( VREG_22_11 ) : ( VREG_22_11 ) ;
assign n41847 =  ( n157 ) ? ( n41845 ) : ( n41846 ) ;
assign n41848 =  ( n6 ) ? ( n41832 ) : ( n41847 ) ;
assign n41849 =  ( n505 ) ? ( n41848 ) : ( VREG_22_11 ) ;
assign n41850 =  ( n148 ) ? ( n10470 ) : ( VREG_22_12 ) ;
assign n41851 =  ( n146 ) ? ( n10469 ) : ( n41850 ) ;
assign n41852 =  ( n144 ) ? ( n10468 ) : ( n41851 ) ;
assign n41853 =  ( n142 ) ? ( n10467 ) : ( n41852 ) ;
assign n41854 =  ( n10 ) ? ( n10466 ) : ( n41853 ) ;
assign n41855 =  ( n148 ) ? ( n11504 ) : ( VREG_22_12 ) ;
assign n41856 =  ( n146 ) ? ( n11503 ) : ( n41855 ) ;
assign n41857 =  ( n144 ) ? ( n11502 ) : ( n41856 ) ;
assign n41858 =  ( n142 ) ? ( n11501 ) : ( n41857 ) ;
assign n41859 =  ( n10 ) ? ( n11500 ) : ( n41858 ) ;
assign n41860 =  ( n11511 ) ? ( VREG_22_12 ) : ( n41854 ) ;
assign n41861 =  ( n11511 ) ? ( VREG_22_12 ) : ( n41859 ) ;
assign n41862 =  ( n3034 ) ? ( n41861 ) : ( VREG_22_12 ) ;
assign n41863 =  ( n2965 ) ? ( n41860 ) : ( n41862 ) ;
assign n41864 =  ( n1930 ) ? ( n41859 ) : ( n41863 ) ;
assign n41865 =  ( n879 ) ? ( n41854 ) : ( n41864 ) ;
assign n41866 =  ( n172 ) ? ( n11522 ) : ( VREG_22_12 ) ;
assign n41867 =  ( n170 ) ? ( n11521 ) : ( n41866 ) ;
assign n41868 =  ( n168 ) ? ( n11520 ) : ( n41867 ) ;
assign n41869 =  ( n166 ) ? ( n11519 ) : ( n41868 ) ;
assign n41870 =  ( n162 ) ? ( n11518 ) : ( n41869 ) ;
assign n41871 =  ( n172 ) ? ( n11532 ) : ( VREG_22_12 ) ;
assign n41872 =  ( n170 ) ? ( n11531 ) : ( n41871 ) ;
assign n41873 =  ( n168 ) ? ( n11530 ) : ( n41872 ) ;
assign n41874 =  ( n166 ) ? ( n11529 ) : ( n41873 ) ;
assign n41875 =  ( n162 ) ? ( n11528 ) : ( n41874 ) ;
assign n41876 =  ( n11511 ) ? ( VREG_22_12 ) : ( n41875 ) ;
assign n41877 =  ( n3051 ) ? ( n41876 ) : ( VREG_22_12 ) ;
assign n41878 =  ( n3040 ) ? ( n41870 ) : ( n41877 ) ;
assign n41879 =  ( n192 ) ? ( VREG_22_12 ) : ( VREG_22_12 ) ;
assign n41880 =  ( n157 ) ? ( n41878 ) : ( n41879 ) ;
assign n41881 =  ( n6 ) ? ( n41865 ) : ( n41880 ) ;
assign n41882 =  ( n505 ) ? ( n41881 ) : ( VREG_22_12 ) ;
assign n41883 =  ( n148 ) ? ( n12589 ) : ( VREG_22_13 ) ;
assign n41884 =  ( n146 ) ? ( n12588 ) : ( n41883 ) ;
assign n41885 =  ( n144 ) ? ( n12587 ) : ( n41884 ) ;
assign n41886 =  ( n142 ) ? ( n12586 ) : ( n41885 ) ;
assign n41887 =  ( n10 ) ? ( n12585 ) : ( n41886 ) ;
assign n41888 =  ( n148 ) ? ( n13623 ) : ( VREG_22_13 ) ;
assign n41889 =  ( n146 ) ? ( n13622 ) : ( n41888 ) ;
assign n41890 =  ( n144 ) ? ( n13621 ) : ( n41889 ) ;
assign n41891 =  ( n142 ) ? ( n13620 ) : ( n41890 ) ;
assign n41892 =  ( n10 ) ? ( n13619 ) : ( n41891 ) ;
assign n41893 =  ( n13630 ) ? ( VREG_22_13 ) : ( n41887 ) ;
assign n41894 =  ( n13630 ) ? ( VREG_22_13 ) : ( n41892 ) ;
assign n41895 =  ( n3034 ) ? ( n41894 ) : ( VREG_22_13 ) ;
assign n41896 =  ( n2965 ) ? ( n41893 ) : ( n41895 ) ;
assign n41897 =  ( n1930 ) ? ( n41892 ) : ( n41896 ) ;
assign n41898 =  ( n879 ) ? ( n41887 ) : ( n41897 ) ;
assign n41899 =  ( n172 ) ? ( n13641 ) : ( VREG_22_13 ) ;
assign n41900 =  ( n170 ) ? ( n13640 ) : ( n41899 ) ;
assign n41901 =  ( n168 ) ? ( n13639 ) : ( n41900 ) ;
assign n41902 =  ( n166 ) ? ( n13638 ) : ( n41901 ) ;
assign n41903 =  ( n162 ) ? ( n13637 ) : ( n41902 ) ;
assign n41904 =  ( n172 ) ? ( n13651 ) : ( VREG_22_13 ) ;
assign n41905 =  ( n170 ) ? ( n13650 ) : ( n41904 ) ;
assign n41906 =  ( n168 ) ? ( n13649 ) : ( n41905 ) ;
assign n41907 =  ( n166 ) ? ( n13648 ) : ( n41906 ) ;
assign n41908 =  ( n162 ) ? ( n13647 ) : ( n41907 ) ;
assign n41909 =  ( n13630 ) ? ( VREG_22_13 ) : ( n41908 ) ;
assign n41910 =  ( n3051 ) ? ( n41909 ) : ( VREG_22_13 ) ;
assign n41911 =  ( n3040 ) ? ( n41903 ) : ( n41910 ) ;
assign n41912 =  ( n192 ) ? ( VREG_22_13 ) : ( VREG_22_13 ) ;
assign n41913 =  ( n157 ) ? ( n41911 ) : ( n41912 ) ;
assign n41914 =  ( n6 ) ? ( n41898 ) : ( n41913 ) ;
assign n41915 =  ( n505 ) ? ( n41914 ) : ( VREG_22_13 ) ;
assign n41916 =  ( n148 ) ? ( n14708 ) : ( VREG_22_14 ) ;
assign n41917 =  ( n146 ) ? ( n14707 ) : ( n41916 ) ;
assign n41918 =  ( n144 ) ? ( n14706 ) : ( n41917 ) ;
assign n41919 =  ( n142 ) ? ( n14705 ) : ( n41918 ) ;
assign n41920 =  ( n10 ) ? ( n14704 ) : ( n41919 ) ;
assign n41921 =  ( n148 ) ? ( n15742 ) : ( VREG_22_14 ) ;
assign n41922 =  ( n146 ) ? ( n15741 ) : ( n41921 ) ;
assign n41923 =  ( n144 ) ? ( n15740 ) : ( n41922 ) ;
assign n41924 =  ( n142 ) ? ( n15739 ) : ( n41923 ) ;
assign n41925 =  ( n10 ) ? ( n15738 ) : ( n41924 ) ;
assign n41926 =  ( n15749 ) ? ( VREG_22_14 ) : ( n41920 ) ;
assign n41927 =  ( n15749 ) ? ( VREG_22_14 ) : ( n41925 ) ;
assign n41928 =  ( n3034 ) ? ( n41927 ) : ( VREG_22_14 ) ;
assign n41929 =  ( n2965 ) ? ( n41926 ) : ( n41928 ) ;
assign n41930 =  ( n1930 ) ? ( n41925 ) : ( n41929 ) ;
assign n41931 =  ( n879 ) ? ( n41920 ) : ( n41930 ) ;
assign n41932 =  ( n172 ) ? ( n15760 ) : ( VREG_22_14 ) ;
assign n41933 =  ( n170 ) ? ( n15759 ) : ( n41932 ) ;
assign n41934 =  ( n168 ) ? ( n15758 ) : ( n41933 ) ;
assign n41935 =  ( n166 ) ? ( n15757 ) : ( n41934 ) ;
assign n41936 =  ( n162 ) ? ( n15756 ) : ( n41935 ) ;
assign n41937 =  ( n172 ) ? ( n15770 ) : ( VREG_22_14 ) ;
assign n41938 =  ( n170 ) ? ( n15769 ) : ( n41937 ) ;
assign n41939 =  ( n168 ) ? ( n15768 ) : ( n41938 ) ;
assign n41940 =  ( n166 ) ? ( n15767 ) : ( n41939 ) ;
assign n41941 =  ( n162 ) ? ( n15766 ) : ( n41940 ) ;
assign n41942 =  ( n15749 ) ? ( VREG_22_14 ) : ( n41941 ) ;
assign n41943 =  ( n3051 ) ? ( n41942 ) : ( VREG_22_14 ) ;
assign n41944 =  ( n3040 ) ? ( n41936 ) : ( n41943 ) ;
assign n41945 =  ( n192 ) ? ( VREG_22_14 ) : ( VREG_22_14 ) ;
assign n41946 =  ( n157 ) ? ( n41944 ) : ( n41945 ) ;
assign n41947 =  ( n6 ) ? ( n41931 ) : ( n41946 ) ;
assign n41948 =  ( n505 ) ? ( n41947 ) : ( VREG_22_14 ) ;
assign n41949 =  ( n148 ) ? ( n16827 ) : ( VREG_22_15 ) ;
assign n41950 =  ( n146 ) ? ( n16826 ) : ( n41949 ) ;
assign n41951 =  ( n144 ) ? ( n16825 ) : ( n41950 ) ;
assign n41952 =  ( n142 ) ? ( n16824 ) : ( n41951 ) ;
assign n41953 =  ( n10 ) ? ( n16823 ) : ( n41952 ) ;
assign n41954 =  ( n148 ) ? ( n17861 ) : ( VREG_22_15 ) ;
assign n41955 =  ( n146 ) ? ( n17860 ) : ( n41954 ) ;
assign n41956 =  ( n144 ) ? ( n17859 ) : ( n41955 ) ;
assign n41957 =  ( n142 ) ? ( n17858 ) : ( n41956 ) ;
assign n41958 =  ( n10 ) ? ( n17857 ) : ( n41957 ) ;
assign n41959 =  ( n17868 ) ? ( VREG_22_15 ) : ( n41953 ) ;
assign n41960 =  ( n17868 ) ? ( VREG_22_15 ) : ( n41958 ) ;
assign n41961 =  ( n3034 ) ? ( n41960 ) : ( VREG_22_15 ) ;
assign n41962 =  ( n2965 ) ? ( n41959 ) : ( n41961 ) ;
assign n41963 =  ( n1930 ) ? ( n41958 ) : ( n41962 ) ;
assign n41964 =  ( n879 ) ? ( n41953 ) : ( n41963 ) ;
assign n41965 =  ( n172 ) ? ( n17879 ) : ( VREG_22_15 ) ;
assign n41966 =  ( n170 ) ? ( n17878 ) : ( n41965 ) ;
assign n41967 =  ( n168 ) ? ( n17877 ) : ( n41966 ) ;
assign n41968 =  ( n166 ) ? ( n17876 ) : ( n41967 ) ;
assign n41969 =  ( n162 ) ? ( n17875 ) : ( n41968 ) ;
assign n41970 =  ( n172 ) ? ( n17889 ) : ( VREG_22_15 ) ;
assign n41971 =  ( n170 ) ? ( n17888 ) : ( n41970 ) ;
assign n41972 =  ( n168 ) ? ( n17887 ) : ( n41971 ) ;
assign n41973 =  ( n166 ) ? ( n17886 ) : ( n41972 ) ;
assign n41974 =  ( n162 ) ? ( n17885 ) : ( n41973 ) ;
assign n41975 =  ( n17868 ) ? ( VREG_22_15 ) : ( n41974 ) ;
assign n41976 =  ( n3051 ) ? ( n41975 ) : ( VREG_22_15 ) ;
assign n41977 =  ( n3040 ) ? ( n41969 ) : ( n41976 ) ;
assign n41978 =  ( n192 ) ? ( VREG_22_15 ) : ( VREG_22_15 ) ;
assign n41979 =  ( n157 ) ? ( n41977 ) : ( n41978 ) ;
assign n41980 =  ( n6 ) ? ( n41964 ) : ( n41979 ) ;
assign n41981 =  ( n505 ) ? ( n41980 ) : ( VREG_22_15 ) ;
assign n41982 =  ( n148 ) ? ( n18946 ) : ( VREG_22_2 ) ;
assign n41983 =  ( n146 ) ? ( n18945 ) : ( n41982 ) ;
assign n41984 =  ( n144 ) ? ( n18944 ) : ( n41983 ) ;
assign n41985 =  ( n142 ) ? ( n18943 ) : ( n41984 ) ;
assign n41986 =  ( n10 ) ? ( n18942 ) : ( n41985 ) ;
assign n41987 =  ( n148 ) ? ( n19980 ) : ( VREG_22_2 ) ;
assign n41988 =  ( n146 ) ? ( n19979 ) : ( n41987 ) ;
assign n41989 =  ( n144 ) ? ( n19978 ) : ( n41988 ) ;
assign n41990 =  ( n142 ) ? ( n19977 ) : ( n41989 ) ;
assign n41991 =  ( n10 ) ? ( n19976 ) : ( n41990 ) ;
assign n41992 =  ( n19987 ) ? ( VREG_22_2 ) : ( n41986 ) ;
assign n41993 =  ( n19987 ) ? ( VREG_22_2 ) : ( n41991 ) ;
assign n41994 =  ( n3034 ) ? ( n41993 ) : ( VREG_22_2 ) ;
assign n41995 =  ( n2965 ) ? ( n41992 ) : ( n41994 ) ;
assign n41996 =  ( n1930 ) ? ( n41991 ) : ( n41995 ) ;
assign n41997 =  ( n879 ) ? ( n41986 ) : ( n41996 ) ;
assign n41998 =  ( n172 ) ? ( n19998 ) : ( VREG_22_2 ) ;
assign n41999 =  ( n170 ) ? ( n19997 ) : ( n41998 ) ;
assign n42000 =  ( n168 ) ? ( n19996 ) : ( n41999 ) ;
assign n42001 =  ( n166 ) ? ( n19995 ) : ( n42000 ) ;
assign n42002 =  ( n162 ) ? ( n19994 ) : ( n42001 ) ;
assign n42003 =  ( n172 ) ? ( n20008 ) : ( VREG_22_2 ) ;
assign n42004 =  ( n170 ) ? ( n20007 ) : ( n42003 ) ;
assign n42005 =  ( n168 ) ? ( n20006 ) : ( n42004 ) ;
assign n42006 =  ( n166 ) ? ( n20005 ) : ( n42005 ) ;
assign n42007 =  ( n162 ) ? ( n20004 ) : ( n42006 ) ;
assign n42008 =  ( n19987 ) ? ( VREG_22_2 ) : ( n42007 ) ;
assign n42009 =  ( n3051 ) ? ( n42008 ) : ( VREG_22_2 ) ;
assign n42010 =  ( n3040 ) ? ( n42002 ) : ( n42009 ) ;
assign n42011 =  ( n192 ) ? ( VREG_22_2 ) : ( VREG_22_2 ) ;
assign n42012 =  ( n157 ) ? ( n42010 ) : ( n42011 ) ;
assign n42013 =  ( n6 ) ? ( n41997 ) : ( n42012 ) ;
assign n42014 =  ( n505 ) ? ( n42013 ) : ( VREG_22_2 ) ;
assign n42015 =  ( n148 ) ? ( n21065 ) : ( VREG_22_3 ) ;
assign n42016 =  ( n146 ) ? ( n21064 ) : ( n42015 ) ;
assign n42017 =  ( n144 ) ? ( n21063 ) : ( n42016 ) ;
assign n42018 =  ( n142 ) ? ( n21062 ) : ( n42017 ) ;
assign n42019 =  ( n10 ) ? ( n21061 ) : ( n42018 ) ;
assign n42020 =  ( n148 ) ? ( n22099 ) : ( VREG_22_3 ) ;
assign n42021 =  ( n146 ) ? ( n22098 ) : ( n42020 ) ;
assign n42022 =  ( n144 ) ? ( n22097 ) : ( n42021 ) ;
assign n42023 =  ( n142 ) ? ( n22096 ) : ( n42022 ) ;
assign n42024 =  ( n10 ) ? ( n22095 ) : ( n42023 ) ;
assign n42025 =  ( n22106 ) ? ( VREG_22_3 ) : ( n42019 ) ;
assign n42026 =  ( n22106 ) ? ( VREG_22_3 ) : ( n42024 ) ;
assign n42027 =  ( n3034 ) ? ( n42026 ) : ( VREG_22_3 ) ;
assign n42028 =  ( n2965 ) ? ( n42025 ) : ( n42027 ) ;
assign n42029 =  ( n1930 ) ? ( n42024 ) : ( n42028 ) ;
assign n42030 =  ( n879 ) ? ( n42019 ) : ( n42029 ) ;
assign n42031 =  ( n172 ) ? ( n22117 ) : ( VREG_22_3 ) ;
assign n42032 =  ( n170 ) ? ( n22116 ) : ( n42031 ) ;
assign n42033 =  ( n168 ) ? ( n22115 ) : ( n42032 ) ;
assign n42034 =  ( n166 ) ? ( n22114 ) : ( n42033 ) ;
assign n42035 =  ( n162 ) ? ( n22113 ) : ( n42034 ) ;
assign n42036 =  ( n172 ) ? ( n22127 ) : ( VREG_22_3 ) ;
assign n42037 =  ( n170 ) ? ( n22126 ) : ( n42036 ) ;
assign n42038 =  ( n168 ) ? ( n22125 ) : ( n42037 ) ;
assign n42039 =  ( n166 ) ? ( n22124 ) : ( n42038 ) ;
assign n42040 =  ( n162 ) ? ( n22123 ) : ( n42039 ) ;
assign n42041 =  ( n22106 ) ? ( VREG_22_3 ) : ( n42040 ) ;
assign n42042 =  ( n3051 ) ? ( n42041 ) : ( VREG_22_3 ) ;
assign n42043 =  ( n3040 ) ? ( n42035 ) : ( n42042 ) ;
assign n42044 =  ( n192 ) ? ( VREG_22_3 ) : ( VREG_22_3 ) ;
assign n42045 =  ( n157 ) ? ( n42043 ) : ( n42044 ) ;
assign n42046 =  ( n6 ) ? ( n42030 ) : ( n42045 ) ;
assign n42047 =  ( n505 ) ? ( n42046 ) : ( VREG_22_3 ) ;
assign n42048 =  ( n148 ) ? ( n23184 ) : ( VREG_22_4 ) ;
assign n42049 =  ( n146 ) ? ( n23183 ) : ( n42048 ) ;
assign n42050 =  ( n144 ) ? ( n23182 ) : ( n42049 ) ;
assign n42051 =  ( n142 ) ? ( n23181 ) : ( n42050 ) ;
assign n42052 =  ( n10 ) ? ( n23180 ) : ( n42051 ) ;
assign n42053 =  ( n148 ) ? ( n24218 ) : ( VREG_22_4 ) ;
assign n42054 =  ( n146 ) ? ( n24217 ) : ( n42053 ) ;
assign n42055 =  ( n144 ) ? ( n24216 ) : ( n42054 ) ;
assign n42056 =  ( n142 ) ? ( n24215 ) : ( n42055 ) ;
assign n42057 =  ( n10 ) ? ( n24214 ) : ( n42056 ) ;
assign n42058 =  ( n24225 ) ? ( VREG_22_4 ) : ( n42052 ) ;
assign n42059 =  ( n24225 ) ? ( VREG_22_4 ) : ( n42057 ) ;
assign n42060 =  ( n3034 ) ? ( n42059 ) : ( VREG_22_4 ) ;
assign n42061 =  ( n2965 ) ? ( n42058 ) : ( n42060 ) ;
assign n42062 =  ( n1930 ) ? ( n42057 ) : ( n42061 ) ;
assign n42063 =  ( n879 ) ? ( n42052 ) : ( n42062 ) ;
assign n42064 =  ( n172 ) ? ( n24236 ) : ( VREG_22_4 ) ;
assign n42065 =  ( n170 ) ? ( n24235 ) : ( n42064 ) ;
assign n42066 =  ( n168 ) ? ( n24234 ) : ( n42065 ) ;
assign n42067 =  ( n166 ) ? ( n24233 ) : ( n42066 ) ;
assign n42068 =  ( n162 ) ? ( n24232 ) : ( n42067 ) ;
assign n42069 =  ( n172 ) ? ( n24246 ) : ( VREG_22_4 ) ;
assign n42070 =  ( n170 ) ? ( n24245 ) : ( n42069 ) ;
assign n42071 =  ( n168 ) ? ( n24244 ) : ( n42070 ) ;
assign n42072 =  ( n166 ) ? ( n24243 ) : ( n42071 ) ;
assign n42073 =  ( n162 ) ? ( n24242 ) : ( n42072 ) ;
assign n42074 =  ( n24225 ) ? ( VREG_22_4 ) : ( n42073 ) ;
assign n42075 =  ( n3051 ) ? ( n42074 ) : ( VREG_22_4 ) ;
assign n42076 =  ( n3040 ) ? ( n42068 ) : ( n42075 ) ;
assign n42077 =  ( n192 ) ? ( VREG_22_4 ) : ( VREG_22_4 ) ;
assign n42078 =  ( n157 ) ? ( n42076 ) : ( n42077 ) ;
assign n42079 =  ( n6 ) ? ( n42063 ) : ( n42078 ) ;
assign n42080 =  ( n505 ) ? ( n42079 ) : ( VREG_22_4 ) ;
assign n42081 =  ( n148 ) ? ( n25303 ) : ( VREG_22_5 ) ;
assign n42082 =  ( n146 ) ? ( n25302 ) : ( n42081 ) ;
assign n42083 =  ( n144 ) ? ( n25301 ) : ( n42082 ) ;
assign n42084 =  ( n142 ) ? ( n25300 ) : ( n42083 ) ;
assign n42085 =  ( n10 ) ? ( n25299 ) : ( n42084 ) ;
assign n42086 =  ( n148 ) ? ( n26337 ) : ( VREG_22_5 ) ;
assign n42087 =  ( n146 ) ? ( n26336 ) : ( n42086 ) ;
assign n42088 =  ( n144 ) ? ( n26335 ) : ( n42087 ) ;
assign n42089 =  ( n142 ) ? ( n26334 ) : ( n42088 ) ;
assign n42090 =  ( n10 ) ? ( n26333 ) : ( n42089 ) ;
assign n42091 =  ( n26344 ) ? ( VREG_22_5 ) : ( n42085 ) ;
assign n42092 =  ( n26344 ) ? ( VREG_22_5 ) : ( n42090 ) ;
assign n42093 =  ( n3034 ) ? ( n42092 ) : ( VREG_22_5 ) ;
assign n42094 =  ( n2965 ) ? ( n42091 ) : ( n42093 ) ;
assign n42095 =  ( n1930 ) ? ( n42090 ) : ( n42094 ) ;
assign n42096 =  ( n879 ) ? ( n42085 ) : ( n42095 ) ;
assign n42097 =  ( n172 ) ? ( n26355 ) : ( VREG_22_5 ) ;
assign n42098 =  ( n170 ) ? ( n26354 ) : ( n42097 ) ;
assign n42099 =  ( n168 ) ? ( n26353 ) : ( n42098 ) ;
assign n42100 =  ( n166 ) ? ( n26352 ) : ( n42099 ) ;
assign n42101 =  ( n162 ) ? ( n26351 ) : ( n42100 ) ;
assign n42102 =  ( n172 ) ? ( n26365 ) : ( VREG_22_5 ) ;
assign n42103 =  ( n170 ) ? ( n26364 ) : ( n42102 ) ;
assign n42104 =  ( n168 ) ? ( n26363 ) : ( n42103 ) ;
assign n42105 =  ( n166 ) ? ( n26362 ) : ( n42104 ) ;
assign n42106 =  ( n162 ) ? ( n26361 ) : ( n42105 ) ;
assign n42107 =  ( n26344 ) ? ( VREG_22_5 ) : ( n42106 ) ;
assign n42108 =  ( n3051 ) ? ( n42107 ) : ( VREG_22_5 ) ;
assign n42109 =  ( n3040 ) ? ( n42101 ) : ( n42108 ) ;
assign n42110 =  ( n192 ) ? ( VREG_22_5 ) : ( VREG_22_5 ) ;
assign n42111 =  ( n157 ) ? ( n42109 ) : ( n42110 ) ;
assign n42112 =  ( n6 ) ? ( n42096 ) : ( n42111 ) ;
assign n42113 =  ( n505 ) ? ( n42112 ) : ( VREG_22_5 ) ;
assign n42114 =  ( n148 ) ? ( n27422 ) : ( VREG_22_6 ) ;
assign n42115 =  ( n146 ) ? ( n27421 ) : ( n42114 ) ;
assign n42116 =  ( n144 ) ? ( n27420 ) : ( n42115 ) ;
assign n42117 =  ( n142 ) ? ( n27419 ) : ( n42116 ) ;
assign n42118 =  ( n10 ) ? ( n27418 ) : ( n42117 ) ;
assign n42119 =  ( n148 ) ? ( n28456 ) : ( VREG_22_6 ) ;
assign n42120 =  ( n146 ) ? ( n28455 ) : ( n42119 ) ;
assign n42121 =  ( n144 ) ? ( n28454 ) : ( n42120 ) ;
assign n42122 =  ( n142 ) ? ( n28453 ) : ( n42121 ) ;
assign n42123 =  ( n10 ) ? ( n28452 ) : ( n42122 ) ;
assign n42124 =  ( n28463 ) ? ( VREG_22_6 ) : ( n42118 ) ;
assign n42125 =  ( n28463 ) ? ( VREG_22_6 ) : ( n42123 ) ;
assign n42126 =  ( n3034 ) ? ( n42125 ) : ( VREG_22_6 ) ;
assign n42127 =  ( n2965 ) ? ( n42124 ) : ( n42126 ) ;
assign n42128 =  ( n1930 ) ? ( n42123 ) : ( n42127 ) ;
assign n42129 =  ( n879 ) ? ( n42118 ) : ( n42128 ) ;
assign n42130 =  ( n172 ) ? ( n28474 ) : ( VREG_22_6 ) ;
assign n42131 =  ( n170 ) ? ( n28473 ) : ( n42130 ) ;
assign n42132 =  ( n168 ) ? ( n28472 ) : ( n42131 ) ;
assign n42133 =  ( n166 ) ? ( n28471 ) : ( n42132 ) ;
assign n42134 =  ( n162 ) ? ( n28470 ) : ( n42133 ) ;
assign n42135 =  ( n172 ) ? ( n28484 ) : ( VREG_22_6 ) ;
assign n42136 =  ( n170 ) ? ( n28483 ) : ( n42135 ) ;
assign n42137 =  ( n168 ) ? ( n28482 ) : ( n42136 ) ;
assign n42138 =  ( n166 ) ? ( n28481 ) : ( n42137 ) ;
assign n42139 =  ( n162 ) ? ( n28480 ) : ( n42138 ) ;
assign n42140 =  ( n28463 ) ? ( VREG_22_6 ) : ( n42139 ) ;
assign n42141 =  ( n3051 ) ? ( n42140 ) : ( VREG_22_6 ) ;
assign n42142 =  ( n3040 ) ? ( n42134 ) : ( n42141 ) ;
assign n42143 =  ( n192 ) ? ( VREG_22_6 ) : ( VREG_22_6 ) ;
assign n42144 =  ( n157 ) ? ( n42142 ) : ( n42143 ) ;
assign n42145 =  ( n6 ) ? ( n42129 ) : ( n42144 ) ;
assign n42146 =  ( n505 ) ? ( n42145 ) : ( VREG_22_6 ) ;
assign n42147 =  ( n148 ) ? ( n29541 ) : ( VREG_22_7 ) ;
assign n42148 =  ( n146 ) ? ( n29540 ) : ( n42147 ) ;
assign n42149 =  ( n144 ) ? ( n29539 ) : ( n42148 ) ;
assign n42150 =  ( n142 ) ? ( n29538 ) : ( n42149 ) ;
assign n42151 =  ( n10 ) ? ( n29537 ) : ( n42150 ) ;
assign n42152 =  ( n148 ) ? ( n30575 ) : ( VREG_22_7 ) ;
assign n42153 =  ( n146 ) ? ( n30574 ) : ( n42152 ) ;
assign n42154 =  ( n144 ) ? ( n30573 ) : ( n42153 ) ;
assign n42155 =  ( n142 ) ? ( n30572 ) : ( n42154 ) ;
assign n42156 =  ( n10 ) ? ( n30571 ) : ( n42155 ) ;
assign n42157 =  ( n30582 ) ? ( VREG_22_7 ) : ( n42151 ) ;
assign n42158 =  ( n30582 ) ? ( VREG_22_7 ) : ( n42156 ) ;
assign n42159 =  ( n3034 ) ? ( n42158 ) : ( VREG_22_7 ) ;
assign n42160 =  ( n2965 ) ? ( n42157 ) : ( n42159 ) ;
assign n42161 =  ( n1930 ) ? ( n42156 ) : ( n42160 ) ;
assign n42162 =  ( n879 ) ? ( n42151 ) : ( n42161 ) ;
assign n42163 =  ( n172 ) ? ( n30593 ) : ( VREG_22_7 ) ;
assign n42164 =  ( n170 ) ? ( n30592 ) : ( n42163 ) ;
assign n42165 =  ( n168 ) ? ( n30591 ) : ( n42164 ) ;
assign n42166 =  ( n166 ) ? ( n30590 ) : ( n42165 ) ;
assign n42167 =  ( n162 ) ? ( n30589 ) : ( n42166 ) ;
assign n42168 =  ( n172 ) ? ( n30603 ) : ( VREG_22_7 ) ;
assign n42169 =  ( n170 ) ? ( n30602 ) : ( n42168 ) ;
assign n42170 =  ( n168 ) ? ( n30601 ) : ( n42169 ) ;
assign n42171 =  ( n166 ) ? ( n30600 ) : ( n42170 ) ;
assign n42172 =  ( n162 ) ? ( n30599 ) : ( n42171 ) ;
assign n42173 =  ( n30582 ) ? ( VREG_22_7 ) : ( n42172 ) ;
assign n42174 =  ( n3051 ) ? ( n42173 ) : ( VREG_22_7 ) ;
assign n42175 =  ( n3040 ) ? ( n42167 ) : ( n42174 ) ;
assign n42176 =  ( n192 ) ? ( VREG_22_7 ) : ( VREG_22_7 ) ;
assign n42177 =  ( n157 ) ? ( n42175 ) : ( n42176 ) ;
assign n42178 =  ( n6 ) ? ( n42162 ) : ( n42177 ) ;
assign n42179 =  ( n505 ) ? ( n42178 ) : ( VREG_22_7 ) ;
assign n42180 =  ( n148 ) ? ( n31660 ) : ( VREG_22_8 ) ;
assign n42181 =  ( n146 ) ? ( n31659 ) : ( n42180 ) ;
assign n42182 =  ( n144 ) ? ( n31658 ) : ( n42181 ) ;
assign n42183 =  ( n142 ) ? ( n31657 ) : ( n42182 ) ;
assign n42184 =  ( n10 ) ? ( n31656 ) : ( n42183 ) ;
assign n42185 =  ( n148 ) ? ( n32694 ) : ( VREG_22_8 ) ;
assign n42186 =  ( n146 ) ? ( n32693 ) : ( n42185 ) ;
assign n42187 =  ( n144 ) ? ( n32692 ) : ( n42186 ) ;
assign n42188 =  ( n142 ) ? ( n32691 ) : ( n42187 ) ;
assign n42189 =  ( n10 ) ? ( n32690 ) : ( n42188 ) ;
assign n42190 =  ( n32701 ) ? ( VREG_22_8 ) : ( n42184 ) ;
assign n42191 =  ( n32701 ) ? ( VREG_22_8 ) : ( n42189 ) ;
assign n42192 =  ( n3034 ) ? ( n42191 ) : ( VREG_22_8 ) ;
assign n42193 =  ( n2965 ) ? ( n42190 ) : ( n42192 ) ;
assign n42194 =  ( n1930 ) ? ( n42189 ) : ( n42193 ) ;
assign n42195 =  ( n879 ) ? ( n42184 ) : ( n42194 ) ;
assign n42196 =  ( n172 ) ? ( n32712 ) : ( VREG_22_8 ) ;
assign n42197 =  ( n170 ) ? ( n32711 ) : ( n42196 ) ;
assign n42198 =  ( n168 ) ? ( n32710 ) : ( n42197 ) ;
assign n42199 =  ( n166 ) ? ( n32709 ) : ( n42198 ) ;
assign n42200 =  ( n162 ) ? ( n32708 ) : ( n42199 ) ;
assign n42201 =  ( n172 ) ? ( n32722 ) : ( VREG_22_8 ) ;
assign n42202 =  ( n170 ) ? ( n32721 ) : ( n42201 ) ;
assign n42203 =  ( n168 ) ? ( n32720 ) : ( n42202 ) ;
assign n42204 =  ( n166 ) ? ( n32719 ) : ( n42203 ) ;
assign n42205 =  ( n162 ) ? ( n32718 ) : ( n42204 ) ;
assign n42206 =  ( n32701 ) ? ( VREG_22_8 ) : ( n42205 ) ;
assign n42207 =  ( n3051 ) ? ( n42206 ) : ( VREG_22_8 ) ;
assign n42208 =  ( n3040 ) ? ( n42200 ) : ( n42207 ) ;
assign n42209 =  ( n192 ) ? ( VREG_22_8 ) : ( VREG_22_8 ) ;
assign n42210 =  ( n157 ) ? ( n42208 ) : ( n42209 ) ;
assign n42211 =  ( n6 ) ? ( n42195 ) : ( n42210 ) ;
assign n42212 =  ( n505 ) ? ( n42211 ) : ( VREG_22_8 ) ;
assign n42213 =  ( n148 ) ? ( n33779 ) : ( VREG_22_9 ) ;
assign n42214 =  ( n146 ) ? ( n33778 ) : ( n42213 ) ;
assign n42215 =  ( n144 ) ? ( n33777 ) : ( n42214 ) ;
assign n42216 =  ( n142 ) ? ( n33776 ) : ( n42215 ) ;
assign n42217 =  ( n10 ) ? ( n33775 ) : ( n42216 ) ;
assign n42218 =  ( n148 ) ? ( n34813 ) : ( VREG_22_9 ) ;
assign n42219 =  ( n146 ) ? ( n34812 ) : ( n42218 ) ;
assign n42220 =  ( n144 ) ? ( n34811 ) : ( n42219 ) ;
assign n42221 =  ( n142 ) ? ( n34810 ) : ( n42220 ) ;
assign n42222 =  ( n10 ) ? ( n34809 ) : ( n42221 ) ;
assign n42223 =  ( n34820 ) ? ( VREG_22_9 ) : ( n42217 ) ;
assign n42224 =  ( n34820 ) ? ( VREG_22_9 ) : ( n42222 ) ;
assign n42225 =  ( n3034 ) ? ( n42224 ) : ( VREG_22_9 ) ;
assign n42226 =  ( n2965 ) ? ( n42223 ) : ( n42225 ) ;
assign n42227 =  ( n1930 ) ? ( n42222 ) : ( n42226 ) ;
assign n42228 =  ( n879 ) ? ( n42217 ) : ( n42227 ) ;
assign n42229 =  ( n172 ) ? ( n34831 ) : ( VREG_22_9 ) ;
assign n42230 =  ( n170 ) ? ( n34830 ) : ( n42229 ) ;
assign n42231 =  ( n168 ) ? ( n34829 ) : ( n42230 ) ;
assign n42232 =  ( n166 ) ? ( n34828 ) : ( n42231 ) ;
assign n42233 =  ( n162 ) ? ( n34827 ) : ( n42232 ) ;
assign n42234 =  ( n172 ) ? ( n34841 ) : ( VREG_22_9 ) ;
assign n42235 =  ( n170 ) ? ( n34840 ) : ( n42234 ) ;
assign n42236 =  ( n168 ) ? ( n34839 ) : ( n42235 ) ;
assign n42237 =  ( n166 ) ? ( n34838 ) : ( n42236 ) ;
assign n42238 =  ( n162 ) ? ( n34837 ) : ( n42237 ) ;
assign n42239 =  ( n34820 ) ? ( VREG_22_9 ) : ( n42238 ) ;
assign n42240 =  ( n3051 ) ? ( n42239 ) : ( VREG_22_9 ) ;
assign n42241 =  ( n3040 ) ? ( n42233 ) : ( n42240 ) ;
assign n42242 =  ( n192 ) ? ( VREG_22_9 ) : ( VREG_22_9 ) ;
assign n42243 =  ( n157 ) ? ( n42241 ) : ( n42242 ) ;
assign n42244 =  ( n6 ) ? ( n42228 ) : ( n42243 ) ;
assign n42245 =  ( n505 ) ? ( n42244 ) : ( VREG_22_9 ) ;
assign n42246 =  ( n148 ) ? ( n1924 ) : ( VREG_23_0 ) ;
assign n42247 =  ( n146 ) ? ( n1923 ) : ( n42246 ) ;
assign n42248 =  ( n144 ) ? ( n1922 ) : ( n42247 ) ;
assign n42249 =  ( n142 ) ? ( n1921 ) : ( n42248 ) ;
assign n42250 =  ( n10 ) ? ( n1920 ) : ( n42249 ) ;
assign n42251 =  ( n148 ) ? ( n2959 ) : ( VREG_23_0 ) ;
assign n42252 =  ( n146 ) ? ( n2958 ) : ( n42251 ) ;
assign n42253 =  ( n144 ) ? ( n2957 ) : ( n42252 ) ;
assign n42254 =  ( n142 ) ? ( n2956 ) : ( n42253 ) ;
assign n42255 =  ( n10 ) ? ( n2955 ) : ( n42254 ) ;
assign n42256 =  ( n3032 ) ? ( VREG_23_0 ) : ( n42250 ) ;
assign n42257 =  ( n3032 ) ? ( VREG_23_0 ) : ( n42255 ) ;
assign n42258 =  ( n3034 ) ? ( n42257 ) : ( VREG_23_0 ) ;
assign n42259 =  ( n2965 ) ? ( n42256 ) : ( n42258 ) ;
assign n42260 =  ( n1930 ) ? ( n42255 ) : ( n42259 ) ;
assign n42261 =  ( n879 ) ? ( n42250 ) : ( n42260 ) ;
assign n42262 =  ( n172 ) ? ( n3045 ) : ( VREG_23_0 ) ;
assign n42263 =  ( n170 ) ? ( n3044 ) : ( n42262 ) ;
assign n42264 =  ( n168 ) ? ( n3043 ) : ( n42263 ) ;
assign n42265 =  ( n166 ) ? ( n3042 ) : ( n42264 ) ;
assign n42266 =  ( n162 ) ? ( n3041 ) : ( n42265 ) ;
assign n42267 =  ( n172 ) ? ( n3056 ) : ( VREG_23_0 ) ;
assign n42268 =  ( n170 ) ? ( n3055 ) : ( n42267 ) ;
assign n42269 =  ( n168 ) ? ( n3054 ) : ( n42268 ) ;
assign n42270 =  ( n166 ) ? ( n3053 ) : ( n42269 ) ;
assign n42271 =  ( n162 ) ? ( n3052 ) : ( n42270 ) ;
assign n42272 =  ( n3032 ) ? ( VREG_23_0 ) : ( n42271 ) ;
assign n42273 =  ( n3051 ) ? ( n42272 ) : ( VREG_23_0 ) ;
assign n42274 =  ( n3040 ) ? ( n42266 ) : ( n42273 ) ;
assign n42275 =  ( n192 ) ? ( VREG_23_0 ) : ( VREG_23_0 ) ;
assign n42276 =  ( n157 ) ? ( n42274 ) : ( n42275 ) ;
assign n42277 =  ( n6 ) ? ( n42261 ) : ( n42276 ) ;
assign n42278 =  ( n527 ) ? ( n42277 ) : ( VREG_23_0 ) ;
assign n42279 =  ( n148 ) ? ( n4113 ) : ( VREG_23_1 ) ;
assign n42280 =  ( n146 ) ? ( n4112 ) : ( n42279 ) ;
assign n42281 =  ( n144 ) ? ( n4111 ) : ( n42280 ) ;
assign n42282 =  ( n142 ) ? ( n4110 ) : ( n42281 ) ;
assign n42283 =  ( n10 ) ? ( n4109 ) : ( n42282 ) ;
assign n42284 =  ( n148 ) ? ( n5147 ) : ( VREG_23_1 ) ;
assign n42285 =  ( n146 ) ? ( n5146 ) : ( n42284 ) ;
assign n42286 =  ( n144 ) ? ( n5145 ) : ( n42285 ) ;
assign n42287 =  ( n142 ) ? ( n5144 ) : ( n42286 ) ;
assign n42288 =  ( n10 ) ? ( n5143 ) : ( n42287 ) ;
assign n42289 =  ( n5154 ) ? ( VREG_23_1 ) : ( n42283 ) ;
assign n42290 =  ( n5154 ) ? ( VREG_23_1 ) : ( n42288 ) ;
assign n42291 =  ( n3034 ) ? ( n42290 ) : ( VREG_23_1 ) ;
assign n42292 =  ( n2965 ) ? ( n42289 ) : ( n42291 ) ;
assign n42293 =  ( n1930 ) ? ( n42288 ) : ( n42292 ) ;
assign n42294 =  ( n879 ) ? ( n42283 ) : ( n42293 ) ;
assign n42295 =  ( n172 ) ? ( n5165 ) : ( VREG_23_1 ) ;
assign n42296 =  ( n170 ) ? ( n5164 ) : ( n42295 ) ;
assign n42297 =  ( n168 ) ? ( n5163 ) : ( n42296 ) ;
assign n42298 =  ( n166 ) ? ( n5162 ) : ( n42297 ) ;
assign n42299 =  ( n162 ) ? ( n5161 ) : ( n42298 ) ;
assign n42300 =  ( n172 ) ? ( n5175 ) : ( VREG_23_1 ) ;
assign n42301 =  ( n170 ) ? ( n5174 ) : ( n42300 ) ;
assign n42302 =  ( n168 ) ? ( n5173 ) : ( n42301 ) ;
assign n42303 =  ( n166 ) ? ( n5172 ) : ( n42302 ) ;
assign n42304 =  ( n162 ) ? ( n5171 ) : ( n42303 ) ;
assign n42305 =  ( n5154 ) ? ( VREG_23_1 ) : ( n42304 ) ;
assign n42306 =  ( n3051 ) ? ( n42305 ) : ( VREG_23_1 ) ;
assign n42307 =  ( n3040 ) ? ( n42299 ) : ( n42306 ) ;
assign n42308 =  ( n192 ) ? ( VREG_23_1 ) : ( VREG_23_1 ) ;
assign n42309 =  ( n157 ) ? ( n42307 ) : ( n42308 ) ;
assign n42310 =  ( n6 ) ? ( n42294 ) : ( n42309 ) ;
assign n42311 =  ( n527 ) ? ( n42310 ) : ( VREG_23_1 ) ;
assign n42312 =  ( n148 ) ? ( n6232 ) : ( VREG_23_10 ) ;
assign n42313 =  ( n146 ) ? ( n6231 ) : ( n42312 ) ;
assign n42314 =  ( n144 ) ? ( n6230 ) : ( n42313 ) ;
assign n42315 =  ( n142 ) ? ( n6229 ) : ( n42314 ) ;
assign n42316 =  ( n10 ) ? ( n6228 ) : ( n42315 ) ;
assign n42317 =  ( n148 ) ? ( n7266 ) : ( VREG_23_10 ) ;
assign n42318 =  ( n146 ) ? ( n7265 ) : ( n42317 ) ;
assign n42319 =  ( n144 ) ? ( n7264 ) : ( n42318 ) ;
assign n42320 =  ( n142 ) ? ( n7263 ) : ( n42319 ) ;
assign n42321 =  ( n10 ) ? ( n7262 ) : ( n42320 ) ;
assign n42322 =  ( n7273 ) ? ( VREG_23_10 ) : ( n42316 ) ;
assign n42323 =  ( n7273 ) ? ( VREG_23_10 ) : ( n42321 ) ;
assign n42324 =  ( n3034 ) ? ( n42323 ) : ( VREG_23_10 ) ;
assign n42325 =  ( n2965 ) ? ( n42322 ) : ( n42324 ) ;
assign n42326 =  ( n1930 ) ? ( n42321 ) : ( n42325 ) ;
assign n42327 =  ( n879 ) ? ( n42316 ) : ( n42326 ) ;
assign n42328 =  ( n172 ) ? ( n7284 ) : ( VREG_23_10 ) ;
assign n42329 =  ( n170 ) ? ( n7283 ) : ( n42328 ) ;
assign n42330 =  ( n168 ) ? ( n7282 ) : ( n42329 ) ;
assign n42331 =  ( n166 ) ? ( n7281 ) : ( n42330 ) ;
assign n42332 =  ( n162 ) ? ( n7280 ) : ( n42331 ) ;
assign n42333 =  ( n172 ) ? ( n7294 ) : ( VREG_23_10 ) ;
assign n42334 =  ( n170 ) ? ( n7293 ) : ( n42333 ) ;
assign n42335 =  ( n168 ) ? ( n7292 ) : ( n42334 ) ;
assign n42336 =  ( n166 ) ? ( n7291 ) : ( n42335 ) ;
assign n42337 =  ( n162 ) ? ( n7290 ) : ( n42336 ) ;
assign n42338 =  ( n7273 ) ? ( VREG_23_10 ) : ( n42337 ) ;
assign n42339 =  ( n3051 ) ? ( n42338 ) : ( VREG_23_10 ) ;
assign n42340 =  ( n3040 ) ? ( n42332 ) : ( n42339 ) ;
assign n42341 =  ( n192 ) ? ( VREG_23_10 ) : ( VREG_23_10 ) ;
assign n42342 =  ( n157 ) ? ( n42340 ) : ( n42341 ) ;
assign n42343 =  ( n6 ) ? ( n42327 ) : ( n42342 ) ;
assign n42344 =  ( n527 ) ? ( n42343 ) : ( VREG_23_10 ) ;
assign n42345 =  ( n148 ) ? ( n8351 ) : ( VREG_23_11 ) ;
assign n42346 =  ( n146 ) ? ( n8350 ) : ( n42345 ) ;
assign n42347 =  ( n144 ) ? ( n8349 ) : ( n42346 ) ;
assign n42348 =  ( n142 ) ? ( n8348 ) : ( n42347 ) ;
assign n42349 =  ( n10 ) ? ( n8347 ) : ( n42348 ) ;
assign n42350 =  ( n148 ) ? ( n9385 ) : ( VREG_23_11 ) ;
assign n42351 =  ( n146 ) ? ( n9384 ) : ( n42350 ) ;
assign n42352 =  ( n144 ) ? ( n9383 ) : ( n42351 ) ;
assign n42353 =  ( n142 ) ? ( n9382 ) : ( n42352 ) ;
assign n42354 =  ( n10 ) ? ( n9381 ) : ( n42353 ) ;
assign n42355 =  ( n9392 ) ? ( VREG_23_11 ) : ( n42349 ) ;
assign n42356 =  ( n9392 ) ? ( VREG_23_11 ) : ( n42354 ) ;
assign n42357 =  ( n3034 ) ? ( n42356 ) : ( VREG_23_11 ) ;
assign n42358 =  ( n2965 ) ? ( n42355 ) : ( n42357 ) ;
assign n42359 =  ( n1930 ) ? ( n42354 ) : ( n42358 ) ;
assign n42360 =  ( n879 ) ? ( n42349 ) : ( n42359 ) ;
assign n42361 =  ( n172 ) ? ( n9403 ) : ( VREG_23_11 ) ;
assign n42362 =  ( n170 ) ? ( n9402 ) : ( n42361 ) ;
assign n42363 =  ( n168 ) ? ( n9401 ) : ( n42362 ) ;
assign n42364 =  ( n166 ) ? ( n9400 ) : ( n42363 ) ;
assign n42365 =  ( n162 ) ? ( n9399 ) : ( n42364 ) ;
assign n42366 =  ( n172 ) ? ( n9413 ) : ( VREG_23_11 ) ;
assign n42367 =  ( n170 ) ? ( n9412 ) : ( n42366 ) ;
assign n42368 =  ( n168 ) ? ( n9411 ) : ( n42367 ) ;
assign n42369 =  ( n166 ) ? ( n9410 ) : ( n42368 ) ;
assign n42370 =  ( n162 ) ? ( n9409 ) : ( n42369 ) ;
assign n42371 =  ( n9392 ) ? ( VREG_23_11 ) : ( n42370 ) ;
assign n42372 =  ( n3051 ) ? ( n42371 ) : ( VREG_23_11 ) ;
assign n42373 =  ( n3040 ) ? ( n42365 ) : ( n42372 ) ;
assign n42374 =  ( n192 ) ? ( VREG_23_11 ) : ( VREG_23_11 ) ;
assign n42375 =  ( n157 ) ? ( n42373 ) : ( n42374 ) ;
assign n42376 =  ( n6 ) ? ( n42360 ) : ( n42375 ) ;
assign n42377 =  ( n527 ) ? ( n42376 ) : ( VREG_23_11 ) ;
assign n42378 =  ( n148 ) ? ( n10470 ) : ( VREG_23_12 ) ;
assign n42379 =  ( n146 ) ? ( n10469 ) : ( n42378 ) ;
assign n42380 =  ( n144 ) ? ( n10468 ) : ( n42379 ) ;
assign n42381 =  ( n142 ) ? ( n10467 ) : ( n42380 ) ;
assign n42382 =  ( n10 ) ? ( n10466 ) : ( n42381 ) ;
assign n42383 =  ( n148 ) ? ( n11504 ) : ( VREG_23_12 ) ;
assign n42384 =  ( n146 ) ? ( n11503 ) : ( n42383 ) ;
assign n42385 =  ( n144 ) ? ( n11502 ) : ( n42384 ) ;
assign n42386 =  ( n142 ) ? ( n11501 ) : ( n42385 ) ;
assign n42387 =  ( n10 ) ? ( n11500 ) : ( n42386 ) ;
assign n42388 =  ( n11511 ) ? ( VREG_23_12 ) : ( n42382 ) ;
assign n42389 =  ( n11511 ) ? ( VREG_23_12 ) : ( n42387 ) ;
assign n42390 =  ( n3034 ) ? ( n42389 ) : ( VREG_23_12 ) ;
assign n42391 =  ( n2965 ) ? ( n42388 ) : ( n42390 ) ;
assign n42392 =  ( n1930 ) ? ( n42387 ) : ( n42391 ) ;
assign n42393 =  ( n879 ) ? ( n42382 ) : ( n42392 ) ;
assign n42394 =  ( n172 ) ? ( n11522 ) : ( VREG_23_12 ) ;
assign n42395 =  ( n170 ) ? ( n11521 ) : ( n42394 ) ;
assign n42396 =  ( n168 ) ? ( n11520 ) : ( n42395 ) ;
assign n42397 =  ( n166 ) ? ( n11519 ) : ( n42396 ) ;
assign n42398 =  ( n162 ) ? ( n11518 ) : ( n42397 ) ;
assign n42399 =  ( n172 ) ? ( n11532 ) : ( VREG_23_12 ) ;
assign n42400 =  ( n170 ) ? ( n11531 ) : ( n42399 ) ;
assign n42401 =  ( n168 ) ? ( n11530 ) : ( n42400 ) ;
assign n42402 =  ( n166 ) ? ( n11529 ) : ( n42401 ) ;
assign n42403 =  ( n162 ) ? ( n11528 ) : ( n42402 ) ;
assign n42404 =  ( n11511 ) ? ( VREG_23_12 ) : ( n42403 ) ;
assign n42405 =  ( n3051 ) ? ( n42404 ) : ( VREG_23_12 ) ;
assign n42406 =  ( n3040 ) ? ( n42398 ) : ( n42405 ) ;
assign n42407 =  ( n192 ) ? ( VREG_23_12 ) : ( VREG_23_12 ) ;
assign n42408 =  ( n157 ) ? ( n42406 ) : ( n42407 ) ;
assign n42409 =  ( n6 ) ? ( n42393 ) : ( n42408 ) ;
assign n42410 =  ( n527 ) ? ( n42409 ) : ( VREG_23_12 ) ;
assign n42411 =  ( n148 ) ? ( n12589 ) : ( VREG_23_13 ) ;
assign n42412 =  ( n146 ) ? ( n12588 ) : ( n42411 ) ;
assign n42413 =  ( n144 ) ? ( n12587 ) : ( n42412 ) ;
assign n42414 =  ( n142 ) ? ( n12586 ) : ( n42413 ) ;
assign n42415 =  ( n10 ) ? ( n12585 ) : ( n42414 ) ;
assign n42416 =  ( n148 ) ? ( n13623 ) : ( VREG_23_13 ) ;
assign n42417 =  ( n146 ) ? ( n13622 ) : ( n42416 ) ;
assign n42418 =  ( n144 ) ? ( n13621 ) : ( n42417 ) ;
assign n42419 =  ( n142 ) ? ( n13620 ) : ( n42418 ) ;
assign n42420 =  ( n10 ) ? ( n13619 ) : ( n42419 ) ;
assign n42421 =  ( n13630 ) ? ( VREG_23_13 ) : ( n42415 ) ;
assign n42422 =  ( n13630 ) ? ( VREG_23_13 ) : ( n42420 ) ;
assign n42423 =  ( n3034 ) ? ( n42422 ) : ( VREG_23_13 ) ;
assign n42424 =  ( n2965 ) ? ( n42421 ) : ( n42423 ) ;
assign n42425 =  ( n1930 ) ? ( n42420 ) : ( n42424 ) ;
assign n42426 =  ( n879 ) ? ( n42415 ) : ( n42425 ) ;
assign n42427 =  ( n172 ) ? ( n13641 ) : ( VREG_23_13 ) ;
assign n42428 =  ( n170 ) ? ( n13640 ) : ( n42427 ) ;
assign n42429 =  ( n168 ) ? ( n13639 ) : ( n42428 ) ;
assign n42430 =  ( n166 ) ? ( n13638 ) : ( n42429 ) ;
assign n42431 =  ( n162 ) ? ( n13637 ) : ( n42430 ) ;
assign n42432 =  ( n172 ) ? ( n13651 ) : ( VREG_23_13 ) ;
assign n42433 =  ( n170 ) ? ( n13650 ) : ( n42432 ) ;
assign n42434 =  ( n168 ) ? ( n13649 ) : ( n42433 ) ;
assign n42435 =  ( n166 ) ? ( n13648 ) : ( n42434 ) ;
assign n42436 =  ( n162 ) ? ( n13647 ) : ( n42435 ) ;
assign n42437 =  ( n13630 ) ? ( VREG_23_13 ) : ( n42436 ) ;
assign n42438 =  ( n3051 ) ? ( n42437 ) : ( VREG_23_13 ) ;
assign n42439 =  ( n3040 ) ? ( n42431 ) : ( n42438 ) ;
assign n42440 =  ( n192 ) ? ( VREG_23_13 ) : ( VREG_23_13 ) ;
assign n42441 =  ( n157 ) ? ( n42439 ) : ( n42440 ) ;
assign n42442 =  ( n6 ) ? ( n42426 ) : ( n42441 ) ;
assign n42443 =  ( n527 ) ? ( n42442 ) : ( VREG_23_13 ) ;
assign n42444 =  ( n148 ) ? ( n14708 ) : ( VREG_23_14 ) ;
assign n42445 =  ( n146 ) ? ( n14707 ) : ( n42444 ) ;
assign n42446 =  ( n144 ) ? ( n14706 ) : ( n42445 ) ;
assign n42447 =  ( n142 ) ? ( n14705 ) : ( n42446 ) ;
assign n42448 =  ( n10 ) ? ( n14704 ) : ( n42447 ) ;
assign n42449 =  ( n148 ) ? ( n15742 ) : ( VREG_23_14 ) ;
assign n42450 =  ( n146 ) ? ( n15741 ) : ( n42449 ) ;
assign n42451 =  ( n144 ) ? ( n15740 ) : ( n42450 ) ;
assign n42452 =  ( n142 ) ? ( n15739 ) : ( n42451 ) ;
assign n42453 =  ( n10 ) ? ( n15738 ) : ( n42452 ) ;
assign n42454 =  ( n15749 ) ? ( VREG_23_14 ) : ( n42448 ) ;
assign n42455 =  ( n15749 ) ? ( VREG_23_14 ) : ( n42453 ) ;
assign n42456 =  ( n3034 ) ? ( n42455 ) : ( VREG_23_14 ) ;
assign n42457 =  ( n2965 ) ? ( n42454 ) : ( n42456 ) ;
assign n42458 =  ( n1930 ) ? ( n42453 ) : ( n42457 ) ;
assign n42459 =  ( n879 ) ? ( n42448 ) : ( n42458 ) ;
assign n42460 =  ( n172 ) ? ( n15760 ) : ( VREG_23_14 ) ;
assign n42461 =  ( n170 ) ? ( n15759 ) : ( n42460 ) ;
assign n42462 =  ( n168 ) ? ( n15758 ) : ( n42461 ) ;
assign n42463 =  ( n166 ) ? ( n15757 ) : ( n42462 ) ;
assign n42464 =  ( n162 ) ? ( n15756 ) : ( n42463 ) ;
assign n42465 =  ( n172 ) ? ( n15770 ) : ( VREG_23_14 ) ;
assign n42466 =  ( n170 ) ? ( n15769 ) : ( n42465 ) ;
assign n42467 =  ( n168 ) ? ( n15768 ) : ( n42466 ) ;
assign n42468 =  ( n166 ) ? ( n15767 ) : ( n42467 ) ;
assign n42469 =  ( n162 ) ? ( n15766 ) : ( n42468 ) ;
assign n42470 =  ( n15749 ) ? ( VREG_23_14 ) : ( n42469 ) ;
assign n42471 =  ( n3051 ) ? ( n42470 ) : ( VREG_23_14 ) ;
assign n42472 =  ( n3040 ) ? ( n42464 ) : ( n42471 ) ;
assign n42473 =  ( n192 ) ? ( VREG_23_14 ) : ( VREG_23_14 ) ;
assign n42474 =  ( n157 ) ? ( n42472 ) : ( n42473 ) ;
assign n42475 =  ( n6 ) ? ( n42459 ) : ( n42474 ) ;
assign n42476 =  ( n527 ) ? ( n42475 ) : ( VREG_23_14 ) ;
assign n42477 =  ( n148 ) ? ( n16827 ) : ( VREG_23_15 ) ;
assign n42478 =  ( n146 ) ? ( n16826 ) : ( n42477 ) ;
assign n42479 =  ( n144 ) ? ( n16825 ) : ( n42478 ) ;
assign n42480 =  ( n142 ) ? ( n16824 ) : ( n42479 ) ;
assign n42481 =  ( n10 ) ? ( n16823 ) : ( n42480 ) ;
assign n42482 =  ( n148 ) ? ( n17861 ) : ( VREG_23_15 ) ;
assign n42483 =  ( n146 ) ? ( n17860 ) : ( n42482 ) ;
assign n42484 =  ( n144 ) ? ( n17859 ) : ( n42483 ) ;
assign n42485 =  ( n142 ) ? ( n17858 ) : ( n42484 ) ;
assign n42486 =  ( n10 ) ? ( n17857 ) : ( n42485 ) ;
assign n42487 =  ( n17868 ) ? ( VREG_23_15 ) : ( n42481 ) ;
assign n42488 =  ( n17868 ) ? ( VREG_23_15 ) : ( n42486 ) ;
assign n42489 =  ( n3034 ) ? ( n42488 ) : ( VREG_23_15 ) ;
assign n42490 =  ( n2965 ) ? ( n42487 ) : ( n42489 ) ;
assign n42491 =  ( n1930 ) ? ( n42486 ) : ( n42490 ) ;
assign n42492 =  ( n879 ) ? ( n42481 ) : ( n42491 ) ;
assign n42493 =  ( n172 ) ? ( n17879 ) : ( VREG_23_15 ) ;
assign n42494 =  ( n170 ) ? ( n17878 ) : ( n42493 ) ;
assign n42495 =  ( n168 ) ? ( n17877 ) : ( n42494 ) ;
assign n42496 =  ( n166 ) ? ( n17876 ) : ( n42495 ) ;
assign n42497 =  ( n162 ) ? ( n17875 ) : ( n42496 ) ;
assign n42498 =  ( n172 ) ? ( n17889 ) : ( VREG_23_15 ) ;
assign n42499 =  ( n170 ) ? ( n17888 ) : ( n42498 ) ;
assign n42500 =  ( n168 ) ? ( n17887 ) : ( n42499 ) ;
assign n42501 =  ( n166 ) ? ( n17886 ) : ( n42500 ) ;
assign n42502 =  ( n162 ) ? ( n17885 ) : ( n42501 ) ;
assign n42503 =  ( n17868 ) ? ( VREG_23_15 ) : ( n42502 ) ;
assign n42504 =  ( n3051 ) ? ( n42503 ) : ( VREG_23_15 ) ;
assign n42505 =  ( n3040 ) ? ( n42497 ) : ( n42504 ) ;
assign n42506 =  ( n192 ) ? ( VREG_23_15 ) : ( VREG_23_15 ) ;
assign n42507 =  ( n157 ) ? ( n42505 ) : ( n42506 ) ;
assign n42508 =  ( n6 ) ? ( n42492 ) : ( n42507 ) ;
assign n42509 =  ( n527 ) ? ( n42508 ) : ( VREG_23_15 ) ;
assign n42510 =  ( n148 ) ? ( n18946 ) : ( VREG_23_2 ) ;
assign n42511 =  ( n146 ) ? ( n18945 ) : ( n42510 ) ;
assign n42512 =  ( n144 ) ? ( n18944 ) : ( n42511 ) ;
assign n42513 =  ( n142 ) ? ( n18943 ) : ( n42512 ) ;
assign n42514 =  ( n10 ) ? ( n18942 ) : ( n42513 ) ;
assign n42515 =  ( n148 ) ? ( n19980 ) : ( VREG_23_2 ) ;
assign n42516 =  ( n146 ) ? ( n19979 ) : ( n42515 ) ;
assign n42517 =  ( n144 ) ? ( n19978 ) : ( n42516 ) ;
assign n42518 =  ( n142 ) ? ( n19977 ) : ( n42517 ) ;
assign n42519 =  ( n10 ) ? ( n19976 ) : ( n42518 ) ;
assign n42520 =  ( n19987 ) ? ( VREG_23_2 ) : ( n42514 ) ;
assign n42521 =  ( n19987 ) ? ( VREG_23_2 ) : ( n42519 ) ;
assign n42522 =  ( n3034 ) ? ( n42521 ) : ( VREG_23_2 ) ;
assign n42523 =  ( n2965 ) ? ( n42520 ) : ( n42522 ) ;
assign n42524 =  ( n1930 ) ? ( n42519 ) : ( n42523 ) ;
assign n42525 =  ( n879 ) ? ( n42514 ) : ( n42524 ) ;
assign n42526 =  ( n172 ) ? ( n19998 ) : ( VREG_23_2 ) ;
assign n42527 =  ( n170 ) ? ( n19997 ) : ( n42526 ) ;
assign n42528 =  ( n168 ) ? ( n19996 ) : ( n42527 ) ;
assign n42529 =  ( n166 ) ? ( n19995 ) : ( n42528 ) ;
assign n42530 =  ( n162 ) ? ( n19994 ) : ( n42529 ) ;
assign n42531 =  ( n172 ) ? ( n20008 ) : ( VREG_23_2 ) ;
assign n42532 =  ( n170 ) ? ( n20007 ) : ( n42531 ) ;
assign n42533 =  ( n168 ) ? ( n20006 ) : ( n42532 ) ;
assign n42534 =  ( n166 ) ? ( n20005 ) : ( n42533 ) ;
assign n42535 =  ( n162 ) ? ( n20004 ) : ( n42534 ) ;
assign n42536 =  ( n19987 ) ? ( VREG_23_2 ) : ( n42535 ) ;
assign n42537 =  ( n3051 ) ? ( n42536 ) : ( VREG_23_2 ) ;
assign n42538 =  ( n3040 ) ? ( n42530 ) : ( n42537 ) ;
assign n42539 =  ( n192 ) ? ( VREG_23_2 ) : ( VREG_23_2 ) ;
assign n42540 =  ( n157 ) ? ( n42538 ) : ( n42539 ) ;
assign n42541 =  ( n6 ) ? ( n42525 ) : ( n42540 ) ;
assign n42542 =  ( n527 ) ? ( n42541 ) : ( VREG_23_2 ) ;
assign n42543 =  ( n148 ) ? ( n21065 ) : ( VREG_23_3 ) ;
assign n42544 =  ( n146 ) ? ( n21064 ) : ( n42543 ) ;
assign n42545 =  ( n144 ) ? ( n21063 ) : ( n42544 ) ;
assign n42546 =  ( n142 ) ? ( n21062 ) : ( n42545 ) ;
assign n42547 =  ( n10 ) ? ( n21061 ) : ( n42546 ) ;
assign n42548 =  ( n148 ) ? ( n22099 ) : ( VREG_23_3 ) ;
assign n42549 =  ( n146 ) ? ( n22098 ) : ( n42548 ) ;
assign n42550 =  ( n144 ) ? ( n22097 ) : ( n42549 ) ;
assign n42551 =  ( n142 ) ? ( n22096 ) : ( n42550 ) ;
assign n42552 =  ( n10 ) ? ( n22095 ) : ( n42551 ) ;
assign n42553 =  ( n22106 ) ? ( VREG_23_3 ) : ( n42547 ) ;
assign n42554 =  ( n22106 ) ? ( VREG_23_3 ) : ( n42552 ) ;
assign n42555 =  ( n3034 ) ? ( n42554 ) : ( VREG_23_3 ) ;
assign n42556 =  ( n2965 ) ? ( n42553 ) : ( n42555 ) ;
assign n42557 =  ( n1930 ) ? ( n42552 ) : ( n42556 ) ;
assign n42558 =  ( n879 ) ? ( n42547 ) : ( n42557 ) ;
assign n42559 =  ( n172 ) ? ( n22117 ) : ( VREG_23_3 ) ;
assign n42560 =  ( n170 ) ? ( n22116 ) : ( n42559 ) ;
assign n42561 =  ( n168 ) ? ( n22115 ) : ( n42560 ) ;
assign n42562 =  ( n166 ) ? ( n22114 ) : ( n42561 ) ;
assign n42563 =  ( n162 ) ? ( n22113 ) : ( n42562 ) ;
assign n42564 =  ( n172 ) ? ( n22127 ) : ( VREG_23_3 ) ;
assign n42565 =  ( n170 ) ? ( n22126 ) : ( n42564 ) ;
assign n42566 =  ( n168 ) ? ( n22125 ) : ( n42565 ) ;
assign n42567 =  ( n166 ) ? ( n22124 ) : ( n42566 ) ;
assign n42568 =  ( n162 ) ? ( n22123 ) : ( n42567 ) ;
assign n42569 =  ( n22106 ) ? ( VREG_23_3 ) : ( n42568 ) ;
assign n42570 =  ( n3051 ) ? ( n42569 ) : ( VREG_23_3 ) ;
assign n42571 =  ( n3040 ) ? ( n42563 ) : ( n42570 ) ;
assign n42572 =  ( n192 ) ? ( VREG_23_3 ) : ( VREG_23_3 ) ;
assign n42573 =  ( n157 ) ? ( n42571 ) : ( n42572 ) ;
assign n42574 =  ( n6 ) ? ( n42558 ) : ( n42573 ) ;
assign n42575 =  ( n527 ) ? ( n42574 ) : ( VREG_23_3 ) ;
assign n42576 =  ( n148 ) ? ( n23184 ) : ( VREG_23_4 ) ;
assign n42577 =  ( n146 ) ? ( n23183 ) : ( n42576 ) ;
assign n42578 =  ( n144 ) ? ( n23182 ) : ( n42577 ) ;
assign n42579 =  ( n142 ) ? ( n23181 ) : ( n42578 ) ;
assign n42580 =  ( n10 ) ? ( n23180 ) : ( n42579 ) ;
assign n42581 =  ( n148 ) ? ( n24218 ) : ( VREG_23_4 ) ;
assign n42582 =  ( n146 ) ? ( n24217 ) : ( n42581 ) ;
assign n42583 =  ( n144 ) ? ( n24216 ) : ( n42582 ) ;
assign n42584 =  ( n142 ) ? ( n24215 ) : ( n42583 ) ;
assign n42585 =  ( n10 ) ? ( n24214 ) : ( n42584 ) ;
assign n42586 =  ( n24225 ) ? ( VREG_23_4 ) : ( n42580 ) ;
assign n42587 =  ( n24225 ) ? ( VREG_23_4 ) : ( n42585 ) ;
assign n42588 =  ( n3034 ) ? ( n42587 ) : ( VREG_23_4 ) ;
assign n42589 =  ( n2965 ) ? ( n42586 ) : ( n42588 ) ;
assign n42590 =  ( n1930 ) ? ( n42585 ) : ( n42589 ) ;
assign n42591 =  ( n879 ) ? ( n42580 ) : ( n42590 ) ;
assign n42592 =  ( n172 ) ? ( n24236 ) : ( VREG_23_4 ) ;
assign n42593 =  ( n170 ) ? ( n24235 ) : ( n42592 ) ;
assign n42594 =  ( n168 ) ? ( n24234 ) : ( n42593 ) ;
assign n42595 =  ( n166 ) ? ( n24233 ) : ( n42594 ) ;
assign n42596 =  ( n162 ) ? ( n24232 ) : ( n42595 ) ;
assign n42597 =  ( n172 ) ? ( n24246 ) : ( VREG_23_4 ) ;
assign n42598 =  ( n170 ) ? ( n24245 ) : ( n42597 ) ;
assign n42599 =  ( n168 ) ? ( n24244 ) : ( n42598 ) ;
assign n42600 =  ( n166 ) ? ( n24243 ) : ( n42599 ) ;
assign n42601 =  ( n162 ) ? ( n24242 ) : ( n42600 ) ;
assign n42602 =  ( n24225 ) ? ( VREG_23_4 ) : ( n42601 ) ;
assign n42603 =  ( n3051 ) ? ( n42602 ) : ( VREG_23_4 ) ;
assign n42604 =  ( n3040 ) ? ( n42596 ) : ( n42603 ) ;
assign n42605 =  ( n192 ) ? ( VREG_23_4 ) : ( VREG_23_4 ) ;
assign n42606 =  ( n157 ) ? ( n42604 ) : ( n42605 ) ;
assign n42607 =  ( n6 ) ? ( n42591 ) : ( n42606 ) ;
assign n42608 =  ( n527 ) ? ( n42607 ) : ( VREG_23_4 ) ;
assign n42609 =  ( n148 ) ? ( n25303 ) : ( VREG_23_5 ) ;
assign n42610 =  ( n146 ) ? ( n25302 ) : ( n42609 ) ;
assign n42611 =  ( n144 ) ? ( n25301 ) : ( n42610 ) ;
assign n42612 =  ( n142 ) ? ( n25300 ) : ( n42611 ) ;
assign n42613 =  ( n10 ) ? ( n25299 ) : ( n42612 ) ;
assign n42614 =  ( n148 ) ? ( n26337 ) : ( VREG_23_5 ) ;
assign n42615 =  ( n146 ) ? ( n26336 ) : ( n42614 ) ;
assign n42616 =  ( n144 ) ? ( n26335 ) : ( n42615 ) ;
assign n42617 =  ( n142 ) ? ( n26334 ) : ( n42616 ) ;
assign n42618 =  ( n10 ) ? ( n26333 ) : ( n42617 ) ;
assign n42619 =  ( n26344 ) ? ( VREG_23_5 ) : ( n42613 ) ;
assign n42620 =  ( n26344 ) ? ( VREG_23_5 ) : ( n42618 ) ;
assign n42621 =  ( n3034 ) ? ( n42620 ) : ( VREG_23_5 ) ;
assign n42622 =  ( n2965 ) ? ( n42619 ) : ( n42621 ) ;
assign n42623 =  ( n1930 ) ? ( n42618 ) : ( n42622 ) ;
assign n42624 =  ( n879 ) ? ( n42613 ) : ( n42623 ) ;
assign n42625 =  ( n172 ) ? ( n26355 ) : ( VREG_23_5 ) ;
assign n42626 =  ( n170 ) ? ( n26354 ) : ( n42625 ) ;
assign n42627 =  ( n168 ) ? ( n26353 ) : ( n42626 ) ;
assign n42628 =  ( n166 ) ? ( n26352 ) : ( n42627 ) ;
assign n42629 =  ( n162 ) ? ( n26351 ) : ( n42628 ) ;
assign n42630 =  ( n172 ) ? ( n26365 ) : ( VREG_23_5 ) ;
assign n42631 =  ( n170 ) ? ( n26364 ) : ( n42630 ) ;
assign n42632 =  ( n168 ) ? ( n26363 ) : ( n42631 ) ;
assign n42633 =  ( n166 ) ? ( n26362 ) : ( n42632 ) ;
assign n42634 =  ( n162 ) ? ( n26361 ) : ( n42633 ) ;
assign n42635 =  ( n26344 ) ? ( VREG_23_5 ) : ( n42634 ) ;
assign n42636 =  ( n3051 ) ? ( n42635 ) : ( VREG_23_5 ) ;
assign n42637 =  ( n3040 ) ? ( n42629 ) : ( n42636 ) ;
assign n42638 =  ( n192 ) ? ( VREG_23_5 ) : ( VREG_23_5 ) ;
assign n42639 =  ( n157 ) ? ( n42637 ) : ( n42638 ) ;
assign n42640 =  ( n6 ) ? ( n42624 ) : ( n42639 ) ;
assign n42641 =  ( n527 ) ? ( n42640 ) : ( VREG_23_5 ) ;
assign n42642 =  ( n148 ) ? ( n27422 ) : ( VREG_23_6 ) ;
assign n42643 =  ( n146 ) ? ( n27421 ) : ( n42642 ) ;
assign n42644 =  ( n144 ) ? ( n27420 ) : ( n42643 ) ;
assign n42645 =  ( n142 ) ? ( n27419 ) : ( n42644 ) ;
assign n42646 =  ( n10 ) ? ( n27418 ) : ( n42645 ) ;
assign n42647 =  ( n148 ) ? ( n28456 ) : ( VREG_23_6 ) ;
assign n42648 =  ( n146 ) ? ( n28455 ) : ( n42647 ) ;
assign n42649 =  ( n144 ) ? ( n28454 ) : ( n42648 ) ;
assign n42650 =  ( n142 ) ? ( n28453 ) : ( n42649 ) ;
assign n42651 =  ( n10 ) ? ( n28452 ) : ( n42650 ) ;
assign n42652 =  ( n28463 ) ? ( VREG_23_6 ) : ( n42646 ) ;
assign n42653 =  ( n28463 ) ? ( VREG_23_6 ) : ( n42651 ) ;
assign n42654 =  ( n3034 ) ? ( n42653 ) : ( VREG_23_6 ) ;
assign n42655 =  ( n2965 ) ? ( n42652 ) : ( n42654 ) ;
assign n42656 =  ( n1930 ) ? ( n42651 ) : ( n42655 ) ;
assign n42657 =  ( n879 ) ? ( n42646 ) : ( n42656 ) ;
assign n42658 =  ( n172 ) ? ( n28474 ) : ( VREG_23_6 ) ;
assign n42659 =  ( n170 ) ? ( n28473 ) : ( n42658 ) ;
assign n42660 =  ( n168 ) ? ( n28472 ) : ( n42659 ) ;
assign n42661 =  ( n166 ) ? ( n28471 ) : ( n42660 ) ;
assign n42662 =  ( n162 ) ? ( n28470 ) : ( n42661 ) ;
assign n42663 =  ( n172 ) ? ( n28484 ) : ( VREG_23_6 ) ;
assign n42664 =  ( n170 ) ? ( n28483 ) : ( n42663 ) ;
assign n42665 =  ( n168 ) ? ( n28482 ) : ( n42664 ) ;
assign n42666 =  ( n166 ) ? ( n28481 ) : ( n42665 ) ;
assign n42667 =  ( n162 ) ? ( n28480 ) : ( n42666 ) ;
assign n42668 =  ( n28463 ) ? ( VREG_23_6 ) : ( n42667 ) ;
assign n42669 =  ( n3051 ) ? ( n42668 ) : ( VREG_23_6 ) ;
assign n42670 =  ( n3040 ) ? ( n42662 ) : ( n42669 ) ;
assign n42671 =  ( n192 ) ? ( VREG_23_6 ) : ( VREG_23_6 ) ;
assign n42672 =  ( n157 ) ? ( n42670 ) : ( n42671 ) ;
assign n42673 =  ( n6 ) ? ( n42657 ) : ( n42672 ) ;
assign n42674 =  ( n527 ) ? ( n42673 ) : ( VREG_23_6 ) ;
assign n42675 =  ( n148 ) ? ( n29541 ) : ( VREG_23_7 ) ;
assign n42676 =  ( n146 ) ? ( n29540 ) : ( n42675 ) ;
assign n42677 =  ( n144 ) ? ( n29539 ) : ( n42676 ) ;
assign n42678 =  ( n142 ) ? ( n29538 ) : ( n42677 ) ;
assign n42679 =  ( n10 ) ? ( n29537 ) : ( n42678 ) ;
assign n42680 =  ( n148 ) ? ( n30575 ) : ( VREG_23_7 ) ;
assign n42681 =  ( n146 ) ? ( n30574 ) : ( n42680 ) ;
assign n42682 =  ( n144 ) ? ( n30573 ) : ( n42681 ) ;
assign n42683 =  ( n142 ) ? ( n30572 ) : ( n42682 ) ;
assign n42684 =  ( n10 ) ? ( n30571 ) : ( n42683 ) ;
assign n42685 =  ( n30582 ) ? ( VREG_23_7 ) : ( n42679 ) ;
assign n42686 =  ( n30582 ) ? ( VREG_23_7 ) : ( n42684 ) ;
assign n42687 =  ( n3034 ) ? ( n42686 ) : ( VREG_23_7 ) ;
assign n42688 =  ( n2965 ) ? ( n42685 ) : ( n42687 ) ;
assign n42689 =  ( n1930 ) ? ( n42684 ) : ( n42688 ) ;
assign n42690 =  ( n879 ) ? ( n42679 ) : ( n42689 ) ;
assign n42691 =  ( n172 ) ? ( n30593 ) : ( VREG_23_7 ) ;
assign n42692 =  ( n170 ) ? ( n30592 ) : ( n42691 ) ;
assign n42693 =  ( n168 ) ? ( n30591 ) : ( n42692 ) ;
assign n42694 =  ( n166 ) ? ( n30590 ) : ( n42693 ) ;
assign n42695 =  ( n162 ) ? ( n30589 ) : ( n42694 ) ;
assign n42696 =  ( n172 ) ? ( n30603 ) : ( VREG_23_7 ) ;
assign n42697 =  ( n170 ) ? ( n30602 ) : ( n42696 ) ;
assign n42698 =  ( n168 ) ? ( n30601 ) : ( n42697 ) ;
assign n42699 =  ( n166 ) ? ( n30600 ) : ( n42698 ) ;
assign n42700 =  ( n162 ) ? ( n30599 ) : ( n42699 ) ;
assign n42701 =  ( n30582 ) ? ( VREG_23_7 ) : ( n42700 ) ;
assign n42702 =  ( n3051 ) ? ( n42701 ) : ( VREG_23_7 ) ;
assign n42703 =  ( n3040 ) ? ( n42695 ) : ( n42702 ) ;
assign n42704 =  ( n192 ) ? ( VREG_23_7 ) : ( VREG_23_7 ) ;
assign n42705 =  ( n157 ) ? ( n42703 ) : ( n42704 ) ;
assign n42706 =  ( n6 ) ? ( n42690 ) : ( n42705 ) ;
assign n42707 =  ( n527 ) ? ( n42706 ) : ( VREG_23_7 ) ;
assign n42708 =  ( n148 ) ? ( n31660 ) : ( VREG_23_8 ) ;
assign n42709 =  ( n146 ) ? ( n31659 ) : ( n42708 ) ;
assign n42710 =  ( n144 ) ? ( n31658 ) : ( n42709 ) ;
assign n42711 =  ( n142 ) ? ( n31657 ) : ( n42710 ) ;
assign n42712 =  ( n10 ) ? ( n31656 ) : ( n42711 ) ;
assign n42713 =  ( n148 ) ? ( n32694 ) : ( VREG_23_8 ) ;
assign n42714 =  ( n146 ) ? ( n32693 ) : ( n42713 ) ;
assign n42715 =  ( n144 ) ? ( n32692 ) : ( n42714 ) ;
assign n42716 =  ( n142 ) ? ( n32691 ) : ( n42715 ) ;
assign n42717 =  ( n10 ) ? ( n32690 ) : ( n42716 ) ;
assign n42718 =  ( n32701 ) ? ( VREG_23_8 ) : ( n42712 ) ;
assign n42719 =  ( n32701 ) ? ( VREG_23_8 ) : ( n42717 ) ;
assign n42720 =  ( n3034 ) ? ( n42719 ) : ( VREG_23_8 ) ;
assign n42721 =  ( n2965 ) ? ( n42718 ) : ( n42720 ) ;
assign n42722 =  ( n1930 ) ? ( n42717 ) : ( n42721 ) ;
assign n42723 =  ( n879 ) ? ( n42712 ) : ( n42722 ) ;
assign n42724 =  ( n172 ) ? ( n32712 ) : ( VREG_23_8 ) ;
assign n42725 =  ( n170 ) ? ( n32711 ) : ( n42724 ) ;
assign n42726 =  ( n168 ) ? ( n32710 ) : ( n42725 ) ;
assign n42727 =  ( n166 ) ? ( n32709 ) : ( n42726 ) ;
assign n42728 =  ( n162 ) ? ( n32708 ) : ( n42727 ) ;
assign n42729 =  ( n172 ) ? ( n32722 ) : ( VREG_23_8 ) ;
assign n42730 =  ( n170 ) ? ( n32721 ) : ( n42729 ) ;
assign n42731 =  ( n168 ) ? ( n32720 ) : ( n42730 ) ;
assign n42732 =  ( n166 ) ? ( n32719 ) : ( n42731 ) ;
assign n42733 =  ( n162 ) ? ( n32718 ) : ( n42732 ) ;
assign n42734 =  ( n32701 ) ? ( VREG_23_8 ) : ( n42733 ) ;
assign n42735 =  ( n3051 ) ? ( n42734 ) : ( VREG_23_8 ) ;
assign n42736 =  ( n3040 ) ? ( n42728 ) : ( n42735 ) ;
assign n42737 =  ( n192 ) ? ( VREG_23_8 ) : ( VREG_23_8 ) ;
assign n42738 =  ( n157 ) ? ( n42736 ) : ( n42737 ) ;
assign n42739 =  ( n6 ) ? ( n42723 ) : ( n42738 ) ;
assign n42740 =  ( n527 ) ? ( n42739 ) : ( VREG_23_8 ) ;
assign n42741 =  ( n148 ) ? ( n33779 ) : ( VREG_23_9 ) ;
assign n42742 =  ( n146 ) ? ( n33778 ) : ( n42741 ) ;
assign n42743 =  ( n144 ) ? ( n33777 ) : ( n42742 ) ;
assign n42744 =  ( n142 ) ? ( n33776 ) : ( n42743 ) ;
assign n42745 =  ( n10 ) ? ( n33775 ) : ( n42744 ) ;
assign n42746 =  ( n148 ) ? ( n34813 ) : ( VREG_23_9 ) ;
assign n42747 =  ( n146 ) ? ( n34812 ) : ( n42746 ) ;
assign n42748 =  ( n144 ) ? ( n34811 ) : ( n42747 ) ;
assign n42749 =  ( n142 ) ? ( n34810 ) : ( n42748 ) ;
assign n42750 =  ( n10 ) ? ( n34809 ) : ( n42749 ) ;
assign n42751 =  ( n34820 ) ? ( VREG_23_9 ) : ( n42745 ) ;
assign n42752 =  ( n34820 ) ? ( VREG_23_9 ) : ( n42750 ) ;
assign n42753 =  ( n3034 ) ? ( n42752 ) : ( VREG_23_9 ) ;
assign n42754 =  ( n2965 ) ? ( n42751 ) : ( n42753 ) ;
assign n42755 =  ( n1930 ) ? ( n42750 ) : ( n42754 ) ;
assign n42756 =  ( n879 ) ? ( n42745 ) : ( n42755 ) ;
assign n42757 =  ( n172 ) ? ( n34831 ) : ( VREG_23_9 ) ;
assign n42758 =  ( n170 ) ? ( n34830 ) : ( n42757 ) ;
assign n42759 =  ( n168 ) ? ( n34829 ) : ( n42758 ) ;
assign n42760 =  ( n166 ) ? ( n34828 ) : ( n42759 ) ;
assign n42761 =  ( n162 ) ? ( n34827 ) : ( n42760 ) ;
assign n42762 =  ( n172 ) ? ( n34841 ) : ( VREG_23_9 ) ;
assign n42763 =  ( n170 ) ? ( n34840 ) : ( n42762 ) ;
assign n42764 =  ( n168 ) ? ( n34839 ) : ( n42763 ) ;
assign n42765 =  ( n166 ) ? ( n34838 ) : ( n42764 ) ;
assign n42766 =  ( n162 ) ? ( n34837 ) : ( n42765 ) ;
assign n42767 =  ( n34820 ) ? ( VREG_23_9 ) : ( n42766 ) ;
assign n42768 =  ( n3051 ) ? ( n42767 ) : ( VREG_23_9 ) ;
assign n42769 =  ( n3040 ) ? ( n42761 ) : ( n42768 ) ;
assign n42770 =  ( n192 ) ? ( VREG_23_9 ) : ( VREG_23_9 ) ;
assign n42771 =  ( n157 ) ? ( n42769 ) : ( n42770 ) ;
assign n42772 =  ( n6 ) ? ( n42756 ) : ( n42771 ) ;
assign n42773 =  ( n527 ) ? ( n42772 ) : ( VREG_23_9 ) ;
assign n42774 =  ( n148 ) ? ( n1924 ) : ( VREG_24_0 ) ;
assign n42775 =  ( n146 ) ? ( n1923 ) : ( n42774 ) ;
assign n42776 =  ( n144 ) ? ( n1922 ) : ( n42775 ) ;
assign n42777 =  ( n142 ) ? ( n1921 ) : ( n42776 ) ;
assign n42778 =  ( n10 ) ? ( n1920 ) : ( n42777 ) ;
assign n42779 =  ( n148 ) ? ( n2959 ) : ( VREG_24_0 ) ;
assign n42780 =  ( n146 ) ? ( n2958 ) : ( n42779 ) ;
assign n42781 =  ( n144 ) ? ( n2957 ) : ( n42780 ) ;
assign n42782 =  ( n142 ) ? ( n2956 ) : ( n42781 ) ;
assign n42783 =  ( n10 ) ? ( n2955 ) : ( n42782 ) ;
assign n42784 =  ( n3032 ) ? ( VREG_24_0 ) : ( n42778 ) ;
assign n42785 =  ( n3032 ) ? ( VREG_24_0 ) : ( n42783 ) ;
assign n42786 =  ( n3034 ) ? ( n42785 ) : ( VREG_24_0 ) ;
assign n42787 =  ( n2965 ) ? ( n42784 ) : ( n42786 ) ;
assign n42788 =  ( n1930 ) ? ( n42783 ) : ( n42787 ) ;
assign n42789 =  ( n879 ) ? ( n42778 ) : ( n42788 ) ;
assign n42790 =  ( n172 ) ? ( n3045 ) : ( VREG_24_0 ) ;
assign n42791 =  ( n170 ) ? ( n3044 ) : ( n42790 ) ;
assign n42792 =  ( n168 ) ? ( n3043 ) : ( n42791 ) ;
assign n42793 =  ( n166 ) ? ( n3042 ) : ( n42792 ) ;
assign n42794 =  ( n162 ) ? ( n3041 ) : ( n42793 ) ;
assign n42795 =  ( n172 ) ? ( n3056 ) : ( VREG_24_0 ) ;
assign n42796 =  ( n170 ) ? ( n3055 ) : ( n42795 ) ;
assign n42797 =  ( n168 ) ? ( n3054 ) : ( n42796 ) ;
assign n42798 =  ( n166 ) ? ( n3053 ) : ( n42797 ) ;
assign n42799 =  ( n162 ) ? ( n3052 ) : ( n42798 ) ;
assign n42800 =  ( n3032 ) ? ( VREG_24_0 ) : ( n42799 ) ;
assign n42801 =  ( n3051 ) ? ( n42800 ) : ( VREG_24_0 ) ;
assign n42802 =  ( n3040 ) ? ( n42794 ) : ( n42801 ) ;
assign n42803 =  ( n192 ) ? ( VREG_24_0 ) : ( VREG_24_0 ) ;
assign n42804 =  ( n157 ) ? ( n42802 ) : ( n42803 ) ;
assign n42805 =  ( n6 ) ? ( n42789 ) : ( n42804 ) ;
assign n42806 =  ( n549 ) ? ( n42805 ) : ( VREG_24_0 ) ;
assign n42807 =  ( n148 ) ? ( n4113 ) : ( VREG_24_1 ) ;
assign n42808 =  ( n146 ) ? ( n4112 ) : ( n42807 ) ;
assign n42809 =  ( n144 ) ? ( n4111 ) : ( n42808 ) ;
assign n42810 =  ( n142 ) ? ( n4110 ) : ( n42809 ) ;
assign n42811 =  ( n10 ) ? ( n4109 ) : ( n42810 ) ;
assign n42812 =  ( n148 ) ? ( n5147 ) : ( VREG_24_1 ) ;
assign n42813 =  ( n146 ) ? ( n5146 ) : ( n42812 ) ;
assign n42814 =  ( n144 ) ? ( n5145 ) : ( n42813 ) ;
assign n42815 =  ( n142 ) ? ( n5144 ) : ( n42814 ) ;
assign n42816 =  ( n10 ) ? ( n5143 ) : ( n42815 ) ;
assign n42817 =  ( n5154 ) ? ( VREG_24_1 ) : ( n42811 ) ;
assign n42818 =  ( n5154 ) ? ( VREG_24_1 ) : ( n42816 ) ;
assign n42819 =  ( n3034 ) ? ( n42818 ) : ( VREG_24_1 ) ;
assign n42820 =  ( n2965 ) ? ( n42817 ) : ( n42819 ) ;
assign n42821 =  ( n1930 ) ? ( n42816 ) : ( n42820 ) ;
assign n42822 =  ( n879 ) ? ( n42811 ) : ( n42821 ) ;
assign n42823 =  ( n172 ) ? ( n5165 ) : ( VREG_24_1 ) ;
assign n42824 =  ( n170 ) ? ( n5164 ) : ( n42823 ) ;
assign n42825 =  ( n168 ) ? ( n5163 ) : ( n42824 ) ;
assign n42826 =  ( n166 ) ? ( n5162 ) : ( n42825 ) ;
assign n42827 =  ( n162 ) ? ( n5161 ) : ( n42826 ) ;
assign n42828 =  ( n172 ) ? ( n5175 ) : ( VREG_24_1 ) ;
assign n42829 =  ( n170 ) ? ( n5174 ) : ( n42828 ) ;
assign n42830 =  ( n168 ) ? ( n5173 ) : ( n42829 ) ;
assign n42831 =  ( n166 ) ? ( n5172 ) : ( n42830 ) ;
assign n42832 =  ( n162 ) ? ( n5171 ) : ( n42831 ) ;
assign n42833 =  ( n5154 ) ? ( VREG_24_1 ) : ( n42832 ) ;
assign n42834 =  ( n3051 ) ? ( n42833 ) : ( VREG_24_1 ) ;
assign n42835 =  ( n3040 ) ? ( n42827 ) : ( n42834 ) ;
assign n42836 =  ( n192 ) ? ( VREG_24_1 ) : ( VREG_24_1 ) ;
assign n42837 =  ( n157 ) ? ( n42835 ) : ( n42836 ) ;
assign n42838 =  ( n6 ) ? ( n42822 ) : ( n42837 ) ;
assign n42839 =  ( n549 ) ? ( n42838 ) : ( VREG_24_1 ) ;
assign n42840 =  ( n148 ) ? ( n6232 ) : ( VREG_24_10 ) ;
assign n42841 =  ( n146 ) ? ( n6231 ) : ( n42840 ) ;
assign n42842 =  ( n144 ) ? ( n6230 ) : ( n42841 ) ;
assign n42843 =  ( n142 ) ? ( n6229 ) : ( n42842 ) ;
assign n42844 =  ( n10 ) ? ( n6228 ) : ( n42843 ) ;
assign n42845 =  ( n148 ) ? ( n7266 ) : ( VREG_24_10 ) ;
assign n42846 =  ( n146 ) ? ( n7265 ) : ( n42845 ) ;
assign n42847 =  ( n144 ) ? ( n7264 ) : ( n42846 ) ;
assign n42848 =  ( n142 ) ? ( n7263 ) : ( n42847 ) ;
assign n42849 =  ( n10 ) ? ( n7262 ) : ( n42848 ) ;
assign n42850 =  ( n7273 ) ? ( VREG_24_10 ) : ( n42844 ) ;
assign n42851 =  ( n7273 ) ? ( VREG_24_10 ) : ( n42849 ) ;
assign n42852 =  ( n3034 ) ? ( n42851 ) : ( VREG_24_10 ) ;
assign n42853 =  ( n2965 ) ? ( n42850 ) : ( n42852 ) ;
assign n42854 =  ( n1930 ) ? ( n42849 ) : ( n42853 ) ;
assign n42855 =  ( n879 ) ? ( n42844 ) : ( n42854 ) ;
assign n42856 =  ( n172 ) ? ( n7284 ) : ( VREG_24_10 ) ;
assign n42857 =  ( n170 ) ? ( n7283 ) : ( n42856 ) ;
assign n42858 =  ( n168 ) ? ( n7282 ) : ( n42857 ) ;
assign n42859 =  ( n166 ) ? ( n7281 ) : ( n42858 ) ;
assign n42860 =  ( n162 ) ? ( n7280 ) : ( n42859 ) ;
assign n42861 =  ( n172 ) ? ( n7294 ) : ( VREG_24_10 ) ;
assign n42862 =  ( n170 ) ? ( n7293 ) : ( n42861 ) ;
assign n42863 =  ( n168 ) ? ( n7292 ) : ( n42862 ) ;
assign n42864 =  ( n166 ) ? ( n7291 ) : ( n42863 ) ;
assign n42865 =  ( n162 ) ? ( n7290 ) : ( n42864 ) ;
assign n42866 =  ( n7273 ) ? ( VREG_24_10 ) : ( n42865 ) ;
assign n42867 =  ( n3051 ) ? ( n42866 ) : ( VREG_24_10 ) ;
assign n42868 =  ( n3040 ) ? ( n42860 ) : ( n42867 ) ;
assign n42869 =  ( n192 ) ? ( VREG_24_10 ) : ( VREG_24_10 ) ;
assign n42870 =  ( n157 ) ? ( n42868 ) : ( n42869 ) ;
assign n42871 =  ( n6 ) ? ( n42855 ) : ( n42870 ) ;
assign n42872 =  ( n549 ) ? ( n42871 ) : ( VREG_24_10 ) ;
assign n42873 =  ( n148 ) ? ( n8351 ) : ( VREG_24_11 ) ;
assign n42874 =  ( n146 ) ? ( n8350 ) : ( n42873 ) ;
assign n42875 =  ( n144 ) ? ( n8349 ) : ( n42874 ) ;
assign n42876 =  ( n142 ) ? ( n8348 ) : ( n42875 ) ;
assign n42877 =  ( n10 ) ? ( n8347 ) : ( n42876 ) ;
assign n42878 =  ( n148 ) ? ( n9385 ) : ( VREG_24_11 ) ;
assign n42879 =  ( n146 ) ? ( n9384 ) : ( n42878 ) ;
assign n42880 =  ( n144 ) ? ( n9383 ) : ( n42879 ) ;
assign n42881 =  ( n142 ) ? ( n9382 ) : ( n42880 ) ;
assign n42882 =  ( n10 ) ? ( n9381 ) : ( n42881 ) ;
assign n42883 =  ( n9392 ) ? ( VREG_24_11 ) : ( n42877 ) ;
assign n42884 =  ( n9392 ) ? ( VREG_24_11 ) : ( n42882 ) ;
assign n42885 =  ( n3034 ) ? ( n42884 ) : ( VREG_24_11 ) ;
assign n42886 =  ( n2965 ) ? ( n42883 ) : ( n42885 ) ;
assign n42887 =  ( n1930 ) ? ( n42882 ) : ( n42886 ) ;
assign n42888 =  ( n879 ) ? ( n42877 ) : ( n42887 ) ;
assign n42889 =  ( n172 ) ? ( n9403 ) : ( VREG_24_11 ) ;
assign n42890 =  ( n170 ) ? ( n9402 ) : ( n42889 ) ;
assign n42891 =  ( n168 ) ? ( n9401 ) : ( n42890 ) ;
assign n42892 =  ( n166 ) ? ( n9400 ) : ( n42891 ) ;
assign n42893 =  ( n162 ) ? ( n9399 ) : ( n42892 ) ;
assign n42894 =  ( n172 ) ? ( n9413 ) : ( VREG_24_11 ) ;
assign n42895 =  ( n170 ) ? ( n9412 ) : ( n42894 ) ;
assign n42896 =  ( n168 ) ? ( n9411 ) : ( n42895 ) ;
assign n42897 =  ( n166 ) ? ( n9410 ) : ( n42896 ) ;
assign n42898 =  ( n162 ) ? ( n9409 ) : ( n42897 ) ;
assign n42899 =  ( n9392 ) ? ( VREG_24_11 ) : ( n42898 ) ;
assign n42900 =  ( n3051 ) ? ( n42899 ) : ( VREG_24_11 ) ;
assign n42901 =  ( n3040 ) ? ( n42893 ) : ( n42900 ) ;
assign n42902 =  ( n192 ) ? ( VREG_24_11 ) : ( VREG_24_11 ) ;
assign n42903 =  ( n157 ) ? ( n42901 ) : ( n42902 ) ;
assign n42904 =  ( n6 ) ? ( n42888 ) : ( n42903 ) ;
assign n42905 =  ( n549 ) ? ( n42904 ) : ( VREG_24_11 ) ;
assign n42906 =  ( n148 ) ? ( n10470 ) : ( VREG_24_12 ) ;
assign n42907 =  ( n146 ) ? ( n10469 ) : ( n42906 ) ;
assign n42908 =  ( n144 ) ? ( n10468 ) : ( n42907 ) ;
assign n42909 =  ( n142 ) ? ( n10467 ) : ( n42908 ) ;
assign n42910 =  ( n10 ) ? ( n10466 ) : ( n42909 ) ;
assign n42911 =  ( n148 ) ? ( n11504 ) : ( VREG_24_12 ) ;
assign n42912 =  ( n146 ) ? ( n11503 ) : ( n42911 ) ;
assign n42913 =  ( n144 ) ? ( n11502 ) : ( n42912 ) ;
assign n42914 =  ( n142 ) ? ( n11501 ) : ( n42913 ) ;
assign n42915 =  ( n10 ) ? ( n11500 ) : ( n42914 ) ;
assign n42916 =  ( n11511 ) ? ( VREG_24_12 ) : ( n42910 ) ;
assign n42917 =  ( n11511 ) ? ( VREG_24_12 ) : ( n42915 ) ;
assign n42918 =  ( n3034 ) ? ( n42917 ) : ( VREG_24_12 ) ;
assign n42919 =  ( n2965 ) ? ( n42916 ) : ( n42918 ) ;
assign n42920 =  ( n1930 ) ? ( n42915 ) : ( n42919 ) ;
assign n42921 =  ( n879 ) ? ( n42910 ) : ( n42920 ) ;
assign n42922 =  ( n172 ) ? ( n11522 ) : ( VREG_24_12 ) ;
assign n42923 =  ( n170 ) ? ( n11521 ) : ( n42922 ) ;
assign n42924 =  ( n168 ) ? ( n11520 ) : ( n42923 ) ;
assign n42925 =  ( n166 ) ? ( n11519 ) : ( n42924 ) ;
assign n42926 =  ( n162 ) ? ( n11518 ) : ( n42925 ) ;
assign n42927 =  ( n172 ) ? ( n11532 ) : ( VREG_24_12 ) ;
assign n42928 =  ( n170 ) ? ( n11531 ) : ( n42927 ) ;
assign n42929 =  ( n168 ) ? ( n11530 ) : ( n42928 ) ;
assign n42930 =  ( n166 ) ? ( n11529 ) : ( n42929 ) ;
assign n42931 =  ( n162 ) ? ( n11528 ) : ( n42930 ) ;
assign n42932 =  ( n11511 ) ? ( VREG_24_12 ) : ( n42931 ) ;
assign n42933 =  ( n3051 ) ? ( n42932 ) : ( VREG_24_12 ) ;
assign n42934 =  ( n3040 ) ? ( n42926 ) : ( n42933 ) ;
assign n42935 =  ( n192 ) ? ( VREG_24_12 ) : ( VREG_24_12 ) ;
assign n42936 =  ( n157 ) ? ( n42934 ) : ( n42935 ) ;
assign n42937 =  ( n6 ) ? ( n42921 ) : ( n42936 ) ;
assign n42938 =  ( n549 ) ? ( n42937 ) : ( VREG_24_12 ) ;
assign n42939 =  ( n148 ) ? ( n12589 ) : ( VREG_24_13 ) ;
assign n42940 =  ( n146 ) ? ( n12588 ) : ( n42939 ) ;
assign n42941 =  ( n144 ) ? ( n12587 ) : ( n42940 ) ;
assign n42942 =  ( n142 ) ? ( n12586 ) : ( n42941 ) ;
assign n42943 =  ( n10 ) ? ( n12585 ) : ( n42942 ) ;
assign n42944 =  ( n148 ) ? ( n13623 ) : ( VREG_24_13 ) ;
assign n42945 =  ( n146 ) ? ( n13622 ) : ( n42944 ) ;
assign n42946 =  ( n144 ) ? ( n13621 ) : ( n42945 ) ;
assign n42947 =  ( n142 ) ? ( n13620 ) : ( n42946 ) ;
assign n42948 =  ( n10 ) ? ( n13619 ) : ( n42947 ) ;
assign n42949 =  ( n13630 ) ? ( VREG_24_13 ) : ( n42943 ) ;
assign n42950 =  ( n13630 ) ? ( VREG_24_13 ) : ( n42948 ) ;
assign n42951 =  ( n3034 ) ? ( n42950 ) : ( VREG_24_13 ) ;
assign n42952 =  ( n2965 ) ? ( n42949 ) : ( n42951 ) ;
assign n42953 =  ( n1930 ) ? ( n42948 ) : ( n42952 ) ;
assign n42954 =  ( n879 ) ? ( n42943 ) : ( n42953 ) ;
assign n42955 =  ( n172 ) ? ( n13641 ) : ( VREG_24_13 ) ;
assign n42956 =  ( n170 ) ? ( n13640 ) : ( n42955 ) ;
assign n42957 =  ( n168 ) ? ( n13639 ) : ( n42956 ) ;
assign n42958 =  ( n166 ) ? ( n13638 ) : ( n42957 ) ;
assign n42959 =  ( n162 ) ? ( n13637 ) : ( n42958 ) ;
assign n42960 =  ( n172 ) ? ( n13651 ) : ( VREG_24_13 ) ;
assign n42961 =  ( n170 ) ? ( n13650 ) : ( n42960 ) ;
assign n42962 =  ( n168 ) ? ( n13649 ) : ( n42961 ) ;
assign n42963 =  ( n166 ) ? ( n13648 ) : ( n42962 ) ;
assign n42964 =  ( n162 ) ? ( n13647 ) : ( n42963 ) ;
assign n42965 =  ( n13630 ) ? ( VREG_24_13 ) : ( n42964 ) ;
assign n42966 =  ( n3051 ) ? ( n42965 ) : ( VREG_24_13 ) ;
assign n42967 =  ( n3040 ) ? ( n42959 ) : ( n42966 ) ;
assign n42968 =  ( n192 ) ? ( VREG_24_13 ) : ( VREG_24_13 ) ;
assign n42969 =  ( n157 ) ? ( n42967 ) : ( n42968 ) ;
assign n42970 =  ( n6 ) ? ( n42954 ) : ( n42969 ) ;
assign n42971 =  ( n549 ) ? ( n42970 ) : ( VREG_24_13 ) ;
assign n42972 =  ( n148 ) ? ( n14708 ) : ( VREG_24_14 ) ;
assign n42973 =  ( n146 ) ? ( n14707 ) : ( n42972 ) ;
assign n42974 =  ( n144 ) ? ( n14706 ) : ( n42973 ) ;
assign n42975 =  ( n142 ) ? ( n14705 ) : ( n42974 ) ;
assign n42976 =  ( n10 ) ? ( n14704 ) : ( n42975 ) ;
assign n42977 =  ( n148 ) ? ( n15742 ) : ( VREG_24_14 ) ;
assign n42978 =  ( n146 ) ? ( n15741 ) : ( n42977 ) ;
assign n42979 =  ( n144 ) ? ( n15740 ) : ( n42978 ) ;
assign n42980 =  ( n142 ) ? ( n15739 ) : ( n42979 ) ;
assign n42981 =  ( n10 ) ? ( n15738 ) : ( n42980 ) ;
assign n42982 =  ( n15749 ) ? ( VREG_24_14 ) : ( n42976 ) ;
assign n42983 =  ( n15749 ) ? ( VREG_24_14 ) : ( n42981 ) ;
assign n42984 =  ( n3034 ) ? ( n42983 ) : ( VREG_24_14 ) ;
assign n42985 =  ( n2965 ) ? ( n42982 ) : ( n42984 ) ;
assign n42986 =  ( n1930 ) ? ( n42981 ) : ( n42985 ) ;
assign n42987 =  ( n879 ) ? ( n42976 ) : ( n42986 ) ;
assign n42988 =  ( n172 ) ? ( n15760 ) : ( VREG_24_14 ) ;
assign n42989 =  ( n170 ) ? ( n15759 ) : ( n42988 ) ;
assign n42990 =  ( n168 ) ? ( n15758 ) : ( n42989 ) ;
assign n42991 =  ( n166 ) ? ( n15757 ) : ( n42990 ) ;
assign n42992 =  ( n162 ) ? ( n15756 ) : ( n42991 ) ;
assign n42993 =  ( n172 ) ? ( n15770 ) : ( VREG_24_14 ) ;
assign n42994 =  ( n170 ) ? ( n15769 ) : ( n42993 ) ;
assign n42995 =  ( n168 ) ? ( n15768 ) : ( n42994 ) ;
assign n42996 =  ( n166 ) ? ( n15767 ) : ( n42995 ) ;
assign n42997 =  ( n162 ) ? ( n15766 ) : ( n42996 ) ;
assign n42998 =  ( n15749 ) ? ( VREG_24_14 ) : ( n42997 ) ;
assign n42999 =  ( n3051 ) ? ( n42998 ) : ( VREG_24_14 ) ;
assign n43000 =  ( n3040 ) ? ( n42992 ) : ( n42999 ) ;
assign n43001 =  ( n192 ) ? ( VREG_24_14 ) : ( VREG_24_14 ) ;
assign n43002 =  ( n157 ) ? ( n43000 ) : ( n43001 ) ;
assign n43003 =  ( n6 ) ? ( n42987 ) : ( n43002 ) ;
assign n43004 =  ( n549 ) ? ( n43003 ) : ( VREG_24_14 ) ;
assign n43005 =  ( n148 ) ? ( n16827 ) : ( VREG_24_15 ) ;
assign n43006 =  ( n146 ) ? ( n16826 ) : ( n43005 ) ;
assign n43007 =  ( n144 ) ? ( n16825 ) : ( n43006 ) ;
assign n43008 =  ( n142 ) ? ( n16824 ) : ( n43007 ) ;
assign n43009 =  ( n10 ) ? ( n16823 ) : ( n43008 ) ;
assign n43010 =  ( n148 ) ? ( n17861 ) : ( VREG_24_15 ) ;
assign n43011 =  ( n146 ) ? ( n17860 ) : ( n43010 ) ;
assign n43012 =  ( n144 ) ? ( n17859 ) : ( n43011 ) ;
assign n43013 =  ( n142 ) ? ( n17858 ) : ( n43012 ) ;
assign n43014 =  ( n10 ) ? ( n17857 ) : ( n43013 ) ;
assign n43015 =  ( n17868 ) ? ( VREG_24_15 ) : ( n43009 ) ;
assign n43016 =  ( n17868 ) ? ( VREG_24_15 ) : ( n43014 ) ;
assign n43017 =  ( n3034 ) ? ( n43016 ) : ( VREG_24_15 ) ;
assign n43018 =  ( n2965 ) ? ( n43015 ) : ( n43017 ) ;
assign n43019 =  ( n1930 ) ? ( n43014 ) : ( n43018 ) ;
assign n43020 =  ( n879 ) ? ( n43009 ) : ( n43019 ) ;
assign n43021 =  ( n172 ) ? ( n17879 ) : ( VREG_24_15 ) ;
assign n43022 =  ( n170 ) ? ( n17878 ) : ( n43021 ) ;
assign n43023 =  ( n168 ) ? ( n17877 ) : ( n43022 ) ;
assign n43024 =  ( n166 ) ? ( n17876 ) : ( n43023 ) ;
assign n43025 =  ( n162 ) ? ( n17875 ) : ( n43024 ) ;
assign n43026 =  ( n172 ) ? ( n17889 ) : ( VREG_24_15 ) ;
assign n43027 =  ( n170 ) ? ( n17888 ) : ( n43026 ) ;
assign n43028 =  ( n168 ) ? ( n17887 ) : ( n43027 ) ;
assign n43029 =  ( n166 ) ? ( n17886 ) : ( n43028 ) ;
assign n43030 =  ( n162 ) ? ( n17885 ) : ( n43029 ) ;
assign n43031 =  ( n17868 ) ? ( VREG_24_15 ) : ( n43030 ) ;
assign n43032 =  ( n3051 ) ? ( n43031 ) : ( VREG_24_15 ) ;
assign n43033 =  ( n3040 ) ? ( n43025 ) : ( n43032 ) ;
assign n43034 =  ( n192 ) ? ( VREG_24_15 ) : ( VREG_24_15 ) ;
assign n43035 =  ( n157 ) ? ( n43033 ) : ( n43034 ) ;
assign n43036 =  ( n6 ) ? ( n43020 ) : ( n43035 ) ;
assign n43037 =  ( n549 ) ? ( n43036 ) : ( VREG_24_15 ) ;
assign n43038 =  ( n148 ) ? ( n18946 ) : ( VREG_24_2 ) ;
assign n43039 =  ( n146 ) ? ( n18945 ) : ( n43038 ) ;
assign n43040 =  ( n144 ) ? ( n18944 ) : ( n43039 ) ;
assign n43041 =  ( n142 ) ? ( n18943 ) : ( n43040 ) ;
assign n43042 =  ( n10 ) ? ( n18942 ) : ( n43041 ) ;
assign n43043 =  ( n148 ) ? ( n19980 ) : ( VREG_24_2 ) ;
assign n43044 =  ( n146 ) ? ( n19979 ) : ( n43043 ) ;
assign n43045 =  ( n144 ) ? ( n19978 ) : ( n43044 ) ;
assign n43046 =  ( n142 ) ? ( n19977 ) : ( n43045 ) ;
assign n43047 =  ( n10 ) ? ( n19976 ) : ( n43046 ) ;
assign n43048 =  ( n19987 ) ? ( VREG_24_2 ) : ( n43042 ) ;
assign n43049 =  ( n19987 ) ? ( VREG_24_2 ) : ( n43047 ) ;
assign n43050 =  ( n3034 ) ? ( n43049 ) : ( VREG_24_2 ) ;
assign n43051 =  ( n2965 ) ? ( n43048 ) : ( n43050 ) ;
assign n43052 =  ( n1930 ) ? ( n43047 ) : ( n43051 ) ;
assign n43053 =  ( n879 ) ? ( n43042 ) : ( n43052 ) ;
assign n43054 =  ( n172 ) ? ( n19998 ) : ( VREG_24_2 ) ;
assign n43055 =  ( n170 ) ? ( n19997 ) : ( n43054 ) ;
assign n43056 =  ( n168 ) ? ( n19996 ) : ( n43055 ) ;
assign n43057 =  ( n166 ) ? ( n19995 ) : ( n43056 ) ;
assign n43058 =  ( n162 ) ? ( n19994 ) : ( n43057 ) ;
assign n43059 =  ( n172 ) ? ( n20008 ) : ( VREG_24_2 ) ;
assign n43060 =  ( n170 ) ? ( n20007 ) : ( n43059 ) ;
assign n43061 =  ( n168 ) ? ( n20006 ) : ( n43060 ) ;
assign n43062 =  ( n166 ) ? ( n20005 ) : ( n43061 ) ;
assign n43063 =  ( n162 ) ? ( n20004 ) : ( n43062 ) ;
assign n43064 =  ( n19987 ) ? ( VREG_24_2 ) : ( n43063 ) ;
assign n43065 =  ( n3051 ) ? ( n43064 ) : ( VREG_24_2 ) ;
assign n43066 =  ( n3040 ) ? ( n43058 ) : ( n43065 ) ;
assign n43067 =  ( n192 ) ? ( VREG_24_2 ) : ( VREG_24_2 ) ;
assign n43068 =  ( n157 ) ? ( n43066 ) : ( n43067 ) ;
assign n43069 =  ( n6 ) ? ( n43053 ) : ( n43068 ) ;
assign n43070 =  ( n549 ) ? ( n43069 ) : ( VREG_24_2 ) ;
assign n43071 =  ( n148 ) ? ( n21065 ) : ( VREG_24_3 ) ;
assign n43072 =  ( n146 ) ? ( n21064 ) : ( n43071 ) ;
assign n43073 =  ( n144 ) ? ( n21063 ) : ( n43072 ) ;
assign n43074 =  ( n142 ) ? ( n21062 ) : ( n43073 ) ;
assign n43075 =  ( n10 ) ? ( n21061 ) : ( n43074 ) ;
assign n43076 =  ( n148 ) ? ( n22099 ) : ( VREG_24_3 ) ;
assign n43077 =  ( n146 ) ? ( n22098 ) : ( n43076 ) ;
assign n43078 =  ( n144 ) ? ( n22097 ) : ( n43077 ) ;
assign n43079 =  ( n142 ) ? ( n22096 ) : ( n43078 ) ;
assign n43080 =  ( n10 ) ? ( n22095 ) : ( n43079 ) ;
assign n43081 =  ( n22106 ) ? ( VREG_24_3 ) : ( n43075 ) ;
assign n43082 =  ( n22106 ) ? ( VREG_24_3 ) : ( n43080 ) ;
assign n43083 =  ( n3034 ) ? ( n43082 ) : ( VREG_24_3 ) ;
assign n43084 =  ( n2965 ) ? ( n43081 ) : ( n43083 ) ;
assign n43085 =  ( n1930 ) ? ( n43080 ) : ( n43084 ) ;
assign n43086 =  ( n879 ) ? ( n43075 ) : ( n43085 ) ;
assign n43087 =  ( n172 ) ? ( n22117 ) : ( VREG_24_3 ) ;
assign n43088 =  ( n170 ) ? ( n22116 ) : ( n43087 ) ;
assign n43089 =  ( n168 ) ? ( n22115 ) : ( n43088 ) ;
assign n43090 =  ( n166 ) ? ( n22114 ) : ( n43089 ) ;
assign n43091 =  ( n162 ) ? ( n22113 ) : ( n43090 ) ;
assign n43092 =  ( n172 ) ? ( n22127 ) : ( VREG_24_3 ) ;
assign n43093 =  ( n170 ) ? ( n22126 ) : ( n43092 ) ;
assign n43094 =  ( n168 ) ? ( n22125 ) : ( n43093 ) ;
assign n43095 =  ( n166 ) ? ( n22124 ) : ( n43094 ) ;
assign n43096 =  ( n162 ) ? ( n22123 ) : ( n43095 ) ;
assign n43097 =  ( n22106 ) ? ( VREG_24_3 ) : ( n43096 ) ;
assign n43098 =  ( n3051 ) ? ( n43097 ) : ( VREG_24_3 ) ;
assign n43099 =  ( n3040 ) ? ( n43091 ) : ( n43098 ) ;
assign n43100 =  ( n192 ) ? ( VREG_24_3 ) : ( VREG_24_3 ) ;
assign n43101 =  ( n157 ) ? ( n43099 ) : ( n43100 ) ;
assign n43102 =  ( n6 ) ? ( n43086 ) : ( n43101 ) ;
assign n43103 =  ( n549 ) ? ( n43102 ) : ( VREG_24_3 ) ;
assign n43104 =  ( n148 ) ? ( n23184 ) : ( VREG_24_4 ) ;
assign n43105 =  ( n146 ) ? ( n23183 ) : ( n43104 ) ;
assign n43106 =  ( n144 ) ? ( n23182 ) : ( n43105 ) ;
assign n43107 =  ( n142 ) ? ( n23181 ) : ( n43106 ) ;
assign n43108 =  ( n10 ) ? ( n23180 ) : ( n43107 ) ;
assign n43109 =  ( n148 ) ? ( n24218 ) : ( VREG_24_4 ) ;
assign n43110 =  ( n146 ) ? ( n24217 ) : ( n43109 ) ;
assign n43111 =  ( n144 ) ? ( n24216 ) : ( n43110 ) ;
assign n43112 =  ( n142 ) ? ( n24215 ) : ( n43111 ) ;
assign n43113 =  ( n10 ) ? ( n24214 ) : ( n43112 ) ;
assign n43114 =  ( n24225 ) ? ( VREG_24_4 ) : ( n43108 ) ;
assign n43115 =  ( n24225 ) ? ( VREG_24_4 ) : ( n43113 ) ;
assign n43116 =  ( n3034 ) ? ( n43115 ) : ( VREG_24_4 ) ;
assign n43117 =  ( n2965 ) ? ( n43114 ) : ( n43116 ) ;
assign n43118 =  ( n1930 ) ? ( n43113 ) : ( n43117 ) ;
assign n43119 =  ( n879 ) ? ( n43108 ) : ( n43118 ) ;
assign n43120 =  ( n172 ) ? ( n24236 ) : ( VREG_24_4 ) ;
assign n43121 =  ( n170 ) ? ( n24235 ) : ( n43120 ) ;
assign n43122 =  ( n168 ) ? ( n24234 ) : ( n43121 ) ;
assign n43123 =  ( n166 ) ? ( n24233 ) : ( n43122 ) ;
assign n43124 =  ( n162 ) ? ( n24232 ) : ( n43123 ) ;
assign n43125 =  ( n172 ) ? ( n24246 ) : ( VREG_24_4 ) ;
assign n43126 =  ( n170 ) ? ( n24245 ) : ( n43125 ) ;
assign n43127 =  ( n168 ) ? ( n24244 ) : ( n43126 ) ;
assign n43128 =  ( n166 ) ? ( n24243 ) : ( n43127 ) ;
assign n43129 =  ( n162 ) ? ( n24242 ) : ( n43128 ) ;
assign n43130 =  ( n24225 ) ? ( VREG_24_4 ) : ( n43129 ) ;
assign n43131 =  ( n3051 ) ? ( n43130 ) : ( VREG_24_4 ) ;
assign n43132 =  ( n3040 ) ? ( n43124 ) : ( n43131 ) ;
assign n43133 =  ( n192 ) ? ( VREG_24_4 ) : ( VREG_24_4 ) ;
assign n43134 =  ( n157 ) ? ( n43132 ) : ( n43133 ) ;
assign n43135 =  ( n6 ) ? ( n43119 ) : ( n43134 ) ;
assign n43136 =  ( n549 ) ? ( n43135 ) : ( VREG_24_4 ) ;
assign n43137 =  ( n148 ) ? ( n25303 ) : ( VREG_24_5 ) ;
assign n43138 =  ( n146 ) ? ( n25302 ) : ( n43137 ) ;
assign n43139 =  ( n144 ) ? ( n25301 ) : ( n43138 ) ;
assign n43140 =  ( n142 ) ? ( n25300 ) : ( n43139 ) ;
assign n43141 =  ( n10 ) ? ( n25299 ) : ( n43140 ) ;
assign n43142 =  ( n148 ) ? ( n26337 ) : ( VREG_24_5 ) ;
assign n43143 =  ( n146 ) ? ( n26336 ) : ( n43142 ) ;
assign n43144 =  ( n144 ) ? ( n26335 ) : ( n43143 ) ;
assign n43145 =  ( n142 ) ? ( n26334 ) : ( n43144 ) ;
assign n43146 =  ( n10 ) ? ( n26333 ) : ( n43145 ) ;
assign n43147 =  ( n26344 ) ? ( VREG_24_5 ) : ( n43141 ) ;
assign n43148 =  ( n26344 ) ? ( VREG_24_5 ) : ( n43146 ) ;
assign n43149 =  ( n3034 ) ? ( n43148 ) : ( VREG_24_5 ) ;
assign n43150 =  ( n2965 ) ? ( n43147 ) : ( n43149 ) ;
assign n43151 =  ( n1930 ) ? ( n43146 ) : ( n43150 ) ;
assign n43152 =  ( n879 ) ? ( n43141 ) : ( n43151 ) ;
assign n43153 =  ( n172 ) ? ( n26355 ) : ( VREG_24_5 ) ;
assign n43154 =  ( n170 ) ? ( n26354 ) : ( n43153 ) ;
assign n43155 =  ( n168 ) ? ( n26353 ) : ( n43154 ) ;
assign n43156 =  ( n166 ) ? ( n26352 ) : ( n43155 ) ;
assign n43157 =  ( n162 ) ? ( n26351 ) : ( n43156 ) ;
assign n43158 =  ( n172 ) ? ( n26365 ) : ( VREG_24_5 ) ;
assign n43159 =  ( n170 ) ? ( n26364 ) : ( n43158 ) ;
assign n43160 =  ( n168 ) ? ( n26363 ) : ( n43159 ) ;
assign n43161 =  ( n166 ) ? ( n26362 ) : ( n43160 ) ;
assign n43162 =  ( n162 ) ? ( n26361 ) : ( n43161 ) ;
assign n43163 =  ( n26344 ) ? ( VREG_24_5 ) : ( n43162 ) ;
assign n43164 =  ( n3051 ) ? ( n43163 ) : ( VREG_24_5 ) ;
assign n43165 =  ( n3040 ) ? ( n43157 ) : ( n43164 ) ;
assign n43166 =  ( n192 ) ? ( VREG_24_5 ) : ( VREG_24_5 ) ;
assign n43167 =  ( n157 ) ? ( n43165 ) : ( n43166 ) ;
assign n43168 =  ( n6 ) ? ( n43152 ) : ( n43167 ) ;
assign n43169 =  ( n549 ) ? ( n43168 ) : ( VREG_24_5 ) ;
assign n43170 =  ( n148 ) ? ( n27422 ) : ( VREG_24_6 ) ;
assign n43171 =  ( n146 ) ? ( n27421 ) : ( n43170 ) ;
assign n43172 =  ( n144 ) ? ( n27420 ) : ( n43171 ) ;
assign n43173 =  ( n142 ) ? ( n27419 ) : ( n43172 ) ;
assign n43174 =  ( n10 ) ? ( n27418 ) : ( n43173 ) ;
assign n43175 =  ( n148 ) ? ( n28456 ) : ( VREG_24_6 ) ;
assign n43176 =  ( n146 ) ? ( n28455 ) : ( n43175 ) ;
assign n43177 =  ( n144 ) ? ( n28454 ) : ( n43176 ) ;
assign n43178 =  ( n142 ) ? ( n28453 ) : ( n43177 ) ;
assign n43179 =  ( n10 ) ? ( n28452 ) : ( n43178 ) ;
assign n43180 =  ( n28463 ) ? ( VREG_24_6 ) : ( n43174 ) ;
assign n43181 =  ( n28463 ) ? ( VREG_24_6 ) : ( n43179 ) ;
assign n43182 =  ( n3034 ) ? ( n43181 ) : ( VREG_24_6 ) ;
assign n43183 =  ( n2965 ) ? ( n43180 ) : ( n43182 ) ;
assign n43184 =  ( n1930 ) ? ( n43179 ) : ( n43183 ) ;
assign n43185 =  ( n879 ) ? ( n43174 ) : ( n43184 ) ;
assign n43186 =  ( n172 ) ? ( n28474 ) : ( VREG_24_6 ) ;
assign n43187 =  ( n170 ) ? ( n28473 ) : ( n43186 ) ;
assign n43188 =  ( n168 ) ? ( n28472 ) : ( n43187 ) ;
assign n43189 =  ( n166 ) ? ( n28471 ) : ( n43188 ) ;
assign n43190 =  ( n162 ) ? ( n28470 ) : ( n43189 ) ;
assign n43191 =  ( n172 ) ? ( n28484 ) : ( VREG_24_6 ) ;
assign n43192 =  ( n170 ) ? ( n28483 ) : ( n43191 ) ;
assign n43193 =  ( n168 ) ? ( n28482 ) : ( n43192 ) ;
assign n43194 =  ( n166 ) ? ( n28481 ) : ( n43193 ) ;
assign n43195 =  ( n162 ) ? ( n28480 ) : ( n43194 ) ;
assign n43196 =  ( n28463 ) ? ( VREG_24_6 ) : ( n43195 ) ;
assign n43197 =  ( n3051 ) ? ( n43196 ) : ( VREG_24_6 ) ;
assign n43198 =  ( n3040 ) ? ( n43190 ) : ( n43197 ) ;
assign n43199 =  ( n192 ) ? ( VREG_24_6 ) : ( VREG_24_6 ) ;
assign n43200 =  ( n157 ) ? ( n43198 ) : ( n43199 ) ;
assign n43201 =  ( n6 ) ? ( n43185 ) : ( n43200 ) ;
assign n43202 =  ( n549 ) ? ( n43201 ) : ( VREG_24_6 ) ;
assign n43203 =  ( n148 ) ? ( n29541 ) : ( VREG_24_7 ) ;
assign n43204 =  ( n146 ) ? ( n29540 ) : ( n43203 ) ;
assign n43205 =  ( n144 ) ? ( n29539 ) : ( n43204 ) ;
assign n43206 =  ( n142 ) ? ( n29538 ) : ( n43205 ) ;
assign n43207 =  ( n10 ) ? ( n29537 ) : ( n43206 ) ;
assign n43208 =  ( n148 ) ? ( n30575 ) : ( VREG_24_7 ) ;
assign n43209 =  ( n146 ) ? ( n30574 ) : ( n43208 ) ;
assign n43210 =  ( n144 ) ? ( n30573 ) : ( n43209 ) ;
assign n43211 =  ( n142 ) ? ( n30572 ) : ( n43210 ) ;
assign n43212 =  ( n10 ) ? ( n30571 ) : ( n43211 ) ;
assign n43213 =  ( n30582 ) ? ( VREG_24_7 ) : ( n43207 ) ;
assign n43214 =  ( n30582 ) ? ( VREG_24_7 ) : ( n43212 ) ;
assign n43215 =  ( n3034 ) ? ( n43214 ) : ( VREG_24_7 ) ;
assign n43216 =  ( n2965 ) ? ( n43213 ) : ( n43215 ) ;
assign n43217 =  ( n1930 ) ? ( n43212 ) : ( n43216 ) ;
assign n43218 =  ( n879 ) ? ( n43207 ) : ( n43217 ) ;
assign n43219 =  ( n172 ) ? ( n30593 ) : ( VREG_24_7 ) ;
assign n43220 =  ( n170 ) ? ( n30592 ) : ( n43219 ) ;
assign n43221 =  ( n168 ) ? ( n30591 ) : ( n43220 ) ;
assign n43222 =  ( n166 ) ? ( n30590 ) : ( n43221 ) ;
assign n43223 =  ( n162 ) ? ( n30589 ) : ( n43222 ) ;
assign n43224 =  ( n172 ) ? ( n30603 ) : ( VREG_24_7 ) ;
assign n43225 =  ( n170 ) ? ( n30602 ) : ( n43224 ) ;
assign n43226 =  ( n168 ) ? ( n30601 ) : ( n43225 ) ;
assign n43227 =  ( n166 ) ? ( n30600 ) : ( n43226 ) ;
assign n43228 =  ( n162 ) ? ( n30599 ) : ( n43227 ) ;
assign n43229 =  ( n30582 ) ? ( VREG_24_7 ) : ( n43228 ) ;
assign n43230 =  ( n3051 ) ? ( n43229 ) : ( VREG_24_7 ) ;
assign n43231 =  ( n3040 ) ? ( n43223 ) : ( n43230 ) ;
assign n43232 =  ( n192 ) ? ( VREG_24_7 ) : ( VREG_24_7 ) ;
assign n43233 =  ( n157 ) ? ( n43231 ) : ( n43232 ) ;
assign n43234 =  ( n6 ) ? ( n43218 ) : ( n43233 ) ;
assign n43235 =  ( n549 ) ? ( n43234 ) : ( VREG_24_7 ) ;
assign n43236 =  ( n148 ) ? ( n31660 ) : ( VREG_24_8 ) ;
assign n43237 =  ( n146 ) ? ( n31659 ) : ( n43236 ) ;
assign n43238 =  ( n144 ) ? ( n31658 ) : ( n43237 ) ;
assign n43239 =  ( n142 ) ? ( n31657 ) : ( n43238 ) ;
assign n43240 =  ( n10 ) ? ( n31656 ) : ( n43239 ) ;
assign n43241 =  ( n148 ) ? ( n32694 ) : ( VREG_24_8 ) ;
assign n43242 =  ( n146 ) ? ( n32693 ) : ( n43241 ) ;
assign n43243 =  ( n144 ) ? ( n32692 ) : ( n43242 ) ;
assign n43244 =  ( n142 ) ? ( n32691 ) : ( n43243 ) ;
assign n43245 =  ( n10 ) ? ( n32690 ) : ( n43244 ) ;
assign n43246 =  ( n32701 ) ? ( VREG_24_8 ) : ( n43240 ) ;
assign n43247 =  ( n32701 ) ? ( VREG_24_8 ) : ( n43245 ) ;
assign n43248 =  ( n3034 ) ? ( n43247 ) : ( VREG_24_8 ) ;
assign n43249 =  ( n2965 ) ? ( n43246 ) : ( n43248 ) ;
assign n43250 =  ( n1930 ) ? ( n43245 ) : ( n43249 ) ;
assign n43251 =  ( n879 ) ? ( n43240 ) : ( n43250 ) ;
assign n43252 =  ( n172 ) ? ( n32712 ) : ( VREG_24_8 ) ;
assign n43253 =  ( n170 ) ? ( n32711 ) : ( n43252 ) ;
assign n43254 =  ( n168 ) ? ( n32710 ) : ( n43253 ) ;
assign n43255 =  ( n166 ) ? ( n32709 ) : ( n43254 ) ;
assign n43256 =  ( n162 ) ? ( n32708 ) : ( n43255 ) ;
assign n43257 =  ( n172 ) ? ( n32722 ) : ( VREG_24_8 ) ;
assign n43258 =  ( n170 ) ? ( n32721 ) : ( n43257 ) ;
assign n43259 =  ( n168 ) ? ( n32720 ) : ( n43258 ) ;
assign n43260 =  ( n166 ) ? ( n32719 ) : ( n43259 ) ;
assign n43261 =  ( n162 ) ? ( n32718 ) : ( n43260 ) ;
assign n43262 =  ( n32701 ) ? ( VREG_24_8 ) : ( n43261 ) ;
assign n43263 =  ( n3051 ) ? ( n43262 ) : ( VREG_24_8 ) ;
assign n43264 =  ( n3040 ) ? ( n43256 ) : ( n43263 ) ;
assign n43265 =  ( n192 ) ? ( VREG_24_8 ) : ( VREG_24_8 ) ;
assign n43266 =  ( n157 ) ? ( n43264 ) : ( n43265 ) ;
assign n43267 =  ( n6 ) ? ( n43251 ) : ( n43266 ) ;
assign n43268 =  ( n549 ) ? ( n43267 ) : ( VREG_24_8 ) ;
assign n43269 =  ( n148 ) ? ( n33779 ) : ( VREG_24_9 ) ;
assign n43270 =  ( n146 ) ? ( n33778 ) : ( n43269 ) ;
assign n43271 =  ( n144 ) ? ( n33777 ) : ( n43270 ) ;
assign n43272 =  ( n142 ) ? ( n33776 ) : ( n43271 ) ;
assign n43273 =  ( n10 ) ? ( n33775 ) : ( n43272 ) ;
assign n43274 =  ( n148 ) ? ( n34813 ) : ( VREG_24_9 ) ;
assign n43275 =  ( n146 ) ? ( n34812 ) : ( n43274 ) ;
assign n43276 =  ( n144 ) ? ( n34811 ) : ( n43275 ) ;
assign n43277 =  ( n142 ) ? ( n34810 ) : ( n43276 ) ;
assign n43278 =  ( n10 ) ? ( n34809 ) : ( n43277 ) ;
assign n43279 =  ( n34820 ) ? ( VREG_24_9 ) : ( n43273 ) ;
assign n43280 =  ( n34820 ) ? ( VREG_24_9 ) : ( n43278 ) ;
assign n43281 =  ( n3034 ) ? ( n43280 ) : ( VREG_24_9 ) ;
assign n43282 =  ( n2965 ) ? ( n43279 ) : ( n43281 ) ;
assign n43283 =  ( n1930 ) ? ( n43278 ) : ( n43282 ) ;
assign n43284 =  ( n879 ) ? ( n43273 ) : ( n43283 ) ;
assign n43285 =  ( n172 ) ? ( n34831 ) : ( VREG_24_9 ) ;
assign n43286 =  ( n170 ) ? ( n34830 ) : ( n43285 ) ;
assign n43287 =  ( n168 ) ? ( n34829 ) : ( n43286 ) ;
assign n43288 =  ( n166 ) ? ( n34828 ) : ( n43287 ) ;
assign n43289 =  ( n162 ) ? ( n34827 ) : ( n43288 ) ;
assign n43290 =  ( n172 ) ? ( n34841 ) : ( VREG_24_9 ) ;
assign n43291 =  ( n170 ) ? ( n34840 ) : ( n43290 ) ;
assign n43292 =  ( n168 ) ? ( n34839 ) : ( n43291 ) ;
assign n43293 =  ( n166 ) ? ( n34838 ) : ( n43292 ) ;
assign n43294 =  ( n162 ) ? ( n34837 ) : ( n43293 ) ;
assign n43295 =  ( n34820 ) ? ( VREG_24_9 ) : ( n43294 ) ;
assign n43296 =  ( n3051 ) ? ( n43295 ) : ( VREG_24_9 ) ;
assign n43297 =  ( n3040 ) ? ( n43289 ) : ( n43296 ) ;
assign n43298 =  ( n192 ) ? ( VREG_24_9 ) : ( VREG_24_9 ) ;
assign n43299 =  ( n157 ) ? ( n43297 ) : ( n43298 ) ;
assign n43300 =  ( n6 ) ? ( n43284 ) : ( n43299 ) ;
assign n43301 =  ( n549 ) ? ( n43300 ) : ( VREG_24_9 ) ;
assign n43302 =  ( n148 ) ? ( n1924 ) : ( VREG_25_0 ) ;
assign n43303 =  ( n146 ) ? ( n1923 ) : ( n43302 ) ;
assign n43304 =  ( n144 ) ? ( n1922 ) : ( n43303 ) ;
assign n43305 =  ( n142 ) ? ( n1921 ) : ( n43304 ) ;
assign n43306 =  ( n10 ) ? ( n1920 ) : ( n43305 ) ;
assign n43307 =  ( n148 ) ? ( n2959 ) : ( VREG_25_0 ) ;
assign n43308 =  ( n146 ) ? ( n2958 ) : ( n43307 ) ;
assign n43309 =  ( n144 ) ? ( n2957 ) : ( n43308 ) ;
assign n43310 =  ( n142 ) ? ( n2956 ) : ( n43309 ) ;
assign n43311 =  ( n10 ) ? ( n2955 ) : ( n43310 ) ;
assign n43312 =  ( n3032 ) ? ( VREG_25_0 ) : ( n43306 ) ;
assign n43313 =  ( n3032 ) ? ( VREG_25_0 ) : ( n43311 ) ;
assign n43314 =  ( n3034 ) ? ( n43313 ) : ( VREG_25_0 ) ;
assign n43315 =  ( n2965 ) ? ( n43312 ) : ( n43314 ) ;
assign n43316 =  ( n1930 ) ? ( n43311 ) : ( n43315 ) ;
assign n43317 =  ( n879 ) ? ( n43306 ) : ( n43316 ) ;
assign n43318 =  ( n172 ) ? ( n3045 ) : ( VREG_25_0 ) ;
assign n43319 =  ( n170 ) ? ( n3044 ) : ( n43318 ) ;
assign n43320 =  ( n168 ) ? ( n3043 ) : ( n43319 ) ;
assign n43321 =  ( n166 ) ? ( n3042 ) : ( n43320 ) ;
assign n43322 =  ( n162 ) ? ( n3041 ) : ( n43321 ) ;
assign n43323 =  ( n172 ) ? ( n3056 ) : ( VREG_25_0 ) ;
assign n43324 =  ( n170 ) ? ( n3055 ) : ( n43323 ) ;
assign n43325 =  ( n168 ) ? ( n3054 ) : ( n43324 ) ;
assign n43326 =  ( n166 ) ? ( n3053 ) : ( n43325 ) ;
assign n43327 =  ( n162 ) ? ( n3052 ) : ( n43326 ) ;
assign n43328 =  ( n3032 ) ? ( VREG_25_0 ) : ( n43327 ) ;
assign n43329 =  ( n3051 ) ? ( n43328 ) : ( VREG_25_0 ) ;
assign n43330 =  ( n3040 ) ? ( n43322 ) : ( n43329 ) ;
assign n43331 =  ( n192 ) ? ( VREG_25_0 ) : ( VREG_25_0 ) ;
assign n43332 =  ( n157 ) ? ( n43330 ) : ( n43331 ) ;
assign n43333 =  ( n6 ) ? ( n43317 ) : ( n43332 ) ;
assign n43334 =  ( n571 ) ? ( n43333 ) : ( VREG_25_0 ) ;
assign n43335 =  ( n148 ) ? ( n4113 ) : ( VREG_25_1 ) ;
assign n43336 =  ( n146 ) ? ( n4112 ) : ( n43335 ) ;
assign n43337 =  ( n144 ) ? ( n4111 ) : ( n43336 ) ;
assign n43338 =  ( n142 ) ? ( n4110 ) : ( n43337 ) ;
assign n43339 =  ( n10 ) ? ( n4109 ) : ( n43338 ) ;
assign n43340 =  ( n148 ) ? ( n5147 ) : ( VREG_25_1 ) ;
assign n43341 =  ( n146 ) ? ( n5146 ) : ( n43340 ) ;
assign n43342 =  ( n144 ) ? ( n5145 ) : ( n43341 ) ;
assign n43343 =  ( n142 ) ? ( n5144 ) : ( n43342 ) ;
assign n43344 =  ( n10 ) ? ( n5143 ) : ( n43343 ) ;
assign n43345 =  ( n5154 ) ? ( VREG_25_1 ) : ( n43339 ) ;
assign n43346 =  ( n5154 ) ? ( VREG_25_1 ) : ( n43344 ) ;
assign n43347 =  ( n3034 ) ? ( n43346 ) : ( VREG_25_1 ) ;
assign n43348 =  ( n2965 ) ? ( n43345 ) : ( n43347 ) ;
assign n43349 =  ( n1930 ) ? ( n43344 ) : ( n43348 ) ;
assign n43350 =  ( n879 ) ? ( n43339 ) : ( n43349 ) ;
assign n43351 =  ( n172 ) ? ( n5165 ) : ( VREG_25_1 ) ;
assign n43352 =  ( n170 ) ? ( n5164 ) : ( n43351 ) ;
assign n43353 =  ( n168 ) ? ( n5163 ) : ( n43352 ) ;
assign n43354 =  ( n166 ) ? ( n5162 ) : ( n43353 ) ;
assign n43355 =  ( n162 ) ? ( n5161 ) : ( n43354 ) ;
assign n43356 =  ( n172 ) ? ( n5175 ) : ( VREG_25_1 ) ;
assign n43357 =  ( n170 ) ? ( n5174 ) : ( n43356 ) ;
assign n43358 =  ( n168 ) ? ( n5173 ) : ( n43357 ) ;
assign n43359 =  ( n166 ) ? ( n5172 ) : ( n43358 ) ;
assign n43360 =  ( n162 ) ? ( n5171 ) : ( n43359 ) ;
assign n43361 =  ( n5154 ) ? ( VREG_25_1 ) : ( n43360 ) ;
assign n43362 =  ( n3051 ) ? ( n43361 ) : ( VREG_25_1 ) ;
assign n43363 =  ( n3040 ) ? ( n43355 ) : ( n43362 ) ;
assign n43364 =  ( n192 ) ? ( VREG_25_1 ) : ( VREG_25_1 ) ;
assign n43365 =  ( n157 ) ? ( n43363 ) : ( n43364 ) ;
assign n43366 =  ( n6 ) ? ( n43350 ) : ( n43365 ) ;
assign n43367 =  ( n571 ) ? ( n43366 ) : ( VREG_25_1 ) ;
assign n43368 =  ( n148 ) ? ( n6232 ) : ( VREG_25_10 ) ;
assign n43369 =  ( n146 ) ? ( n6231 ) : ( n43368 ) ;
assign n43370 =  ( n144 ) ? ( n6230 ) : ( n43369 ) ;
assign n43371 =  ( n142 ) ? ( n6229 ) : ( n43370 ) ;
assign n43372 =  ( n10 ) ? ( n6228 ) : ( n43371 ) ;
assign n43373 =  ( n148 ) ? ( n7266 ) : ( VREG_25_10 ) ;
assign n43374 =  ( n146 ) ? ( n7265 ) : ( n43373 ) ;
assign n43375 =  ( n144 ) ? ( n7264 ) : ( n43374 ) ;
assign n43376 =  ( n142 ) ? ( n7263 ) : ( n43375 ) ;
assign n43377 =  ( n10 ) ? ( n7262 ) : ( n43376 ) ;
assign n43378 =  ( n7273 ) ? ( VREG_25_10 ) : ( n43372 ) ;
assign n43379 =  ( n7273 ) ? ( VREG_25_10 ) : ( n43377 ) ;
assign n43380 =  ( n3034 ) ? ( n43379 ) : ( VREG_25_10 ) ;
assign n43381 =  ( n2965 ) ? ( n43378 ) : ( n43380 ) ;
assign n43382 =  ( n1930 ) ? ( n43377 ) : ( n43381 ) ;
assign n43383 =  ( n879 ) ? ( n43372 ) : ( n43382 ) ;
assign n43384 =  ( n172 ) ? ( n7284 ) : ( VREG_25_10 ) ;
assign n43385 =  ( n170 ) ? ( n7283 ) : ( n43384 ) ;
assign n43386 =  ( n168 ) ? ( n7282 ) : ( n43385 ) ;
assign n43387 =  ( n166 ) ? ( n7281 ) : ( n43386 ) ;
assign n43388 =  ( n162 ) ? ( n7280 ) : ( n43387 ) ;
assign n43389 =  ( n172 ) ? ( n7294 ) : ( VREG_25_10 ) ;
assign n43390 =  ( n170 ) ? ( n7293 ) : ( n43389 ) ;
assign n43391 =  ( n168 ) ? ( n7292 ) : ( n43390 ) ;
assign n43392 =  ( n166 ) ? ( n7291 ) : ( n43391 ) ;
assign n43393 =  ( n162 ) ? ( n7290 ) : ( n43392 ) ;
assign n43394 =  ( n7273 ) ? ( VREG_25_10 ) : ( n43393 ) ;
assign n43395 =  ( n3051 ) ? ( n43394 ) : ( VREG_25_10 ) ;
assign n43396 =  ( n3040 ) ? ( n43388 ) : ( n43395 ) ;
assign n43397 =  ( n192 ) ? ( VREG_25_10 ) : ( VREG_25_10 ) ;
assign n43398 =  ( n157 ) ? ( n43396 ) : ( n43397 ) ;
assign n43399 =  ( n6 ) ? ( n43383 ) : ( n43398 ) ;
assign n43400 =  ( n571 ) ? ( n43399 ) : ( VREG_25_10 ) ;
assign n43401 =  ( n148 ) ? ( n8351 ) : ( VREG_25_11 ) ;
assign n43402 =  ( n146 ) ? ( n8350 ) : ( n43401 ) ;
assign n43403 =  ( n144 ) ? ( n8349 ) : ( n43402 ) ;
assign n43404 =  ( n142 ) ? ( n8348 ) : ( n43403 ) ;
assign n43405 =  ( n10 ) ? ( n8347 ) : ( n43404 ) ;
assign n43406 =  ( n148 ) ? ( n9385 ) : ( VREG_25_11 ) ;
assign n43407 =  ( n146 ) ? ( n9384 ) : ( n43406 ) ;
assign n43408 =  ( n144 ) ? ( n9383 ) : ( n43407 ) ;
assign n43409 =  ( n142 ) ? ( n9382 ) : ( n43408 ) ;
assign n43410 =  ( n10 ) ? ( n9381 ) : ( n43409 ) ;
assign n43411 =  ( n9392 ) ? ( VREG_25_11 ) : ( n43405 ) ;
assign n43412 =  ( n9392 ) ? ( VREG_25_11 ) : ( n43410 ) ;
assign n43413 =  ( n3034 ) ? ( n43412 ) : ( VREG_25_11 ) ;
assign n43414 =  ( n2965 ) ? ( n43411 ) : ( n43413 ) ;
assign n43415 =  ( n1930 ) ? ( n43410 ) : ( n43414 ) ;
assign n43416 =  ( n879 ) ? ( n43405 ) : ( n43415 ) ;
assign n43417 =  ( n172 ) ? ( n9403 ) : ( VREG_25_11 ) ;
assign n43418 =  ( n170 ) ? ( n9402 ) : ( n43417 ) ;
assign n43419 =  ( n168 ) ? ( n9401 ) : ( n43418 ) ;
assign n43420 =  ( n166 ) ? ( n9400 ) : ( n43419 ) ;
assign n43421 =  ( n162 ) ? ( n9399 ) : ( n43420 ) ;
assign n43422 =  ( n172 ) ? ( n9413 ) : ( VREG_25_11 ) ;
assign n43423 =  ( n170 ) ? ( n9412 ) : ( n43422 ) ;
assign n43424 =  ( n168 ) ? ( n9411 ) : ( n43423 ) ;
assign n43425 =  ( n166 ) ? ( n9410 ) : ( n43424 ) ;
assign n43426 =  ( n162 ) ? ( n9409 ) : ( n43425 ) ;
assign n43427 =  ( n9392 ) ? ( VREG_25_11 ) : ( n43426 ) ;
assign n43428 =  ( n3051 ) ? ( n43427 ) : ( VREG_25_11 ) ;
assign n43429 =  ( n3040 ) ? ( n43421 ) : ( n43428 ) ;
assign n43430 =  ( n192 ) ? ( VREG_25_11 ) : ( VREG_25_11 ) ;
assign n43431 =  ( n157 ) ? ( n43429 ) : ( n43430 ) ;
assign n43432 =  ( n6 ) ? ( n43416 ) : ( n43431 ) ;
assign n43433 =  ( n571 ) ? ( n43432 ) : ( VREG_25_11 ) ;
assign n43434 =  ( n148 ) ? ( n10470 ) : ( VREG_25_12 ) ;
assign n43435 =  ( n146 ) ? ( n10469 ) : ( n43434 ) ;
assign n43436 =  ( n144 ) ? ( n10468 ) : ( n43435 ) ;
assign n43437 =  ( n142 ) ? ( n10467 ) : ( n43436 ) ;
assign n43438 =  ( n10 ) ? ( n10466 ) : ( n43437 ) ;
assign n43439 =  ( n148 ) ? ( n11504 ) : ( VREG_25_12 ) ;
assign n43440 =  ( n146 ) ? ( n11503 ) : ( n43439 ) ;
assign n43441 =  ( n144 ) ? ( n11502 ) : ( n43440 ) ;
assign n43442 =  ( n142 ) ? ( n11501 ) : ( n43441 ) ;
assign n43443 =  ( n10 ) ? ( n11500 ) : ( n43442 ) ;
assign n43444 =  ( n11511 ) ? ( VREG_25_12 ) : ( n43438 ) ;
assign n43445 =  ( n11511 ) ? ( VREG_25_12 ) : ( n43443 ) ;
assign n43446 =  ( n3034 ) ? ( n43445 ) : ( VREG_25_12 ) ;
assign n43447 =  ( n2965 ) ? ( n43444 ) : ( n43446 ) ;
assign n43448 =  ( n1930 ) ? ( n43443 ) : ( n43447 ) ;
assign n43449 =  ( n879 ) ? ( n43438 ) : ( n43448 ) ;
assign n43450 =  ( n172 ) ? ( n11522 ) : ( VREG_25_12 ) ;
assign n43451 =  ( n170 ) ? ( n11521 ) : ( n43450 ) ;
assign n43452 =  ( n168 ) ? ( n11520 ) : ( n43451 ) ;
assign n43453 =  ( n166 ) ? ( n11519 ) : ( n43452 ) ;
assign n43454 =  ( n162 ) ? ( n11518 ) : ( n43453 ) ;
assign n43455 =  ( n172 ) ? ( n11532 ) : ( VREG_25_12 ) ;
assign n43456 =  ( n170 ) ? ( n11531 ) : ( n43455 ) ;
assign n43457 =  ( n168 ) ? ( n11530 ) : ( n43456 ) ;
assign n43458 =  ( n166 ) ? ( n11529 ) : ( n43457 ) ;
assign n43459 =  ( n162 ) ? ( n11528 ) : ( n43458 ) ;
assign n43460 =  ( n11511 ) ? ( VREG_25_12 ) : ( n43459 ) ;
assign n43461 =  ( n3051 ) ? ( n43460 ) : ( VREG_25_12 ) ;
assign n43462 =  ( n3040 ) ? ( n43454 ) : ( n43461 ) ;
assign n43463 =  ( n192 ) ? ( VREG_25_12 ) : ( VREG_25_12 ) ;
assign n43464 =  ( n157 ) ? ( n43462 ) : ( n43463 ) ;
assign n43465 =  ( n6 ) ? ( n43449 ) : ( n43464 ) ;
assign n43466 =  ( n571 ) ? ( n43465 ) : ( VREG_25_12 ) ;
assign n43467 =  ( n148 ) ? ( n12589 ) : ( VREG_25_13 ) ;
assign n43468 =  ( n146 ) ? ( n12588 ) : ( n43467 ) ;
assign n43469 =  ( n144 ) ? ( n12587 ) : ( n43468 ) ;
assign n43470 =  ( n142 ) ? ( n12586 ) : ( n43469 ) ;
assign n43471 =  ( n10 ) ? ( n12585 ) : ( n43470 ) ;
assign n43472 =  ( n148 ) ? ( n13623 ) : ( VREG_25_13 ) ;
assign n43473 =  ( n146 ) ? ( n13622 ) : ( n43472 ) ;
assign n43474 =  ( n144 ) ? ( n13621 ) : ( n43473 ) ;
assign n43475 =  ( n142 ) ? ( n13620 ) : ( n43474 ) ;
assign n43476 =  ( n10 ) ? ( n13619 ) : ( n43475 ) ;
assign n43477 =  ( n13630 ) ? ( VREG_25_13 ) : ( n43471 ) ;
assign n43478 =  ( n13630 ) ? ( VREG_25_13 ) : ( n43476 ) ;
assign n43479 =  ( n3034 ) ? ( n43478 ) : ( VREG_25_13 ) ;
assign n43480 =  ( n2965 ) ? ( n43477 ) : ( n43479 ) ;
assign n43481 =  ( n1930 ) ? ( n43476 ) : ( n43480 ) ;
assign n43482 =  ( n879 ) ? ( n43471 ) : ( n43481 ) ;
assign n43483 =  ( n172 ) ? ( n13641 ) : ( VREG_25_13 ) ;
assign n43484 =  ( n170 ) ? ( n13640 ) : ( n43483 ) ;
assign n43485 =  ( n168 ) ? ( n13639 ) : ( n43484 ) ;
assign n43486 =  ( n166 ) ? ( n13638 ) : ( n43485 ) ;
assign n43487 =  ( n162 ) ? ( n13637 ) : ( n43486 ) ;
assign n43488 =  ( n172 ) ? ( n13651 ) : ( VREG_25_13 ) ;
assign n43489 =  ( n170 ) ? ( n13650 ) : ( n43488 ) ;
assign n43490 =  ( n168 ) ? ( n13649 ) : ( n43489 ) ;
assign n43491 =  ( n166 ) ? ( n13648 ) : ( n43490 ) ;
assign n43492 =  ( n162 ) ? ( n13647 ) : ( n43491 ) ;
assign n43493 =  ( n13630 ) ? ( VREG_25_13 ) : ( n43492 ) ;
assign n43494 =  ( n3051 ) ? ( n43493 ) : ( VREG_25_13 ) ;
assign n43495 =  ( n3040 ) ? ( n43487 ) : ( n43494 ) ;
assign n43496 =  ( n192 ) ? ( VREG_25_13 ) : ( VREG_25_13 ) ;
assign n43497 =  ( n157 ) ? ( n43495 ) : ( n43496 ) ;
assign n43498 =  ( n6 ) ? ( n43482 ) : ( n43497 ) ;
assign n43499 =  ( n571 ) ? ( n43498 ) : ( VREG_25_13 ) ;
assign n43500 =  ( n148 ) ? ( n14708 ) : ( VREG_25_14 ) ;
assign n43501 =  ( n146 ) ? ( n14707 ) : ( n43500 ) ;
assign n43502 =  ( n144 ) ? ( n14706 ) : ( n43501 ) ;
assign n43503 =  ( n142 ) ? ( n14705 ) : ( n43502 ) ;
assign n43504 =  ( n10 ) ? ( n14704 ) : ( n43503 ) ;
assign n43505 =  ( n148 ) ? ( n15742 ) : ( VREG_25_14 ) ;
assign n43506 =  ( n146 ) ? ( n15741 ) : ( n43505 ) ;
assign n43507 =  ( n144 ) ? ( n15740 ) : ( n43506 ) ;
assign n43508 =  ( n142 ) ? ( n15739 ) : ( n43507 ) ;
assign n43509 =  ( n10 ) ? ( n15738 ) : ( n43508 ) ;
assign n43510 =  ( n15749 ) ? ( VREG_25_14 ) : ( n43504 ) ;
assign n43511 =  ( n15749 ) ? ( VREG_25_14 ) : ( n43509 ) ;
assign n43512 =  ( n3034 ) ? ( n43511 ) : ( VREG_25_14 ) ;
assign n43513 =  ( n2965 ) ? ( n43510 ) : ( n43512 ) ;
assign n43514 =  ( n1930 ) ? ( n43509 ) : ( n43513 ) ;
assign n43515 =  ( n879 ) ? ( n43504 ) : ( n43514 ) ;
assign n43516 =  ( n172 ) ? ( n15760 ) : ( VREG_25_14 ) ;
assign n43517 =  ( n170 ) ? ( n15759 ) : ( n43516 ) ;
assign n43518 =  ( n168 ) ? ( n15758 ) : ( n43517 ) ;
assign n43519 =  ( n166 ) ? ( n15757 ) : ( n43518 ) ;
assign n43520 =  ( n162 ) ? ( n15756 ) : ( n43519 ) ;
assign n43521 =  ( n172 ) ? ( n15770 ) : ( VREG_25_14 ) ;
assign n43522 =  ( n170 ) ? ( n15769 ) : ( n43521 ) ;
assign n43523 =  ( n168 ) ? ( n15768 ) : ( n43522 ) ;
assign n43524 =  ( n166 ) ? ( n15767 ) : ( n43523 ) ;
assign n43525 =  ( n162 ) ? ( n15766 ) : ( n43524 ) ;
assign n43526 =  ( n15749 ) ? ( VREG_25_14 ) : ( n43525 ) ;
assign n43527 =  ( n3051 ) ? ( n43526 ) : ( VREG_25_14 ) ;
assign n43528 =  ( n3040 ) ? ( n43520 ) : ( n43527 ) ;
assign n43529 =  ( n192 ) ? ( VREG_25_14 ) : ( VREG_25_14 ) ;
assign n43530 =  ( n157 ) ? ( n43528 ) : ( n43529 ) ;
assign n43531 =  ( n6 ) ? ( n43515 ) : ( n43530 ) ;
assign n43532 =  ( n571 ) ? ( n43531 ) : ( VREG_25_14 ) ;
assign n43533 =  ( n148 ) ? ( n16827 ) : ( VREG_25_15 ) ;
assign n43534 =  ( n146 ) ? ( n16826 ) : ( n43533 ) ;
assign n43535 =  ( n144 ) ? ( n16825 ) : ( n43534 ) ;
assign n43536 =  ( n142 ) ? ( n16824 ) : ( n43535 ) ;
assign n43537 =  ( n10 ) ? ( n16823 ) : ( n43536 ) ;
assign n43538 =  ( n148 ) ? ( n17861 ) : ( VREG_25_15 ) ;
assign n43539 =  ( n146 ) ? ( n17860 ) : ( n43538 ) ;
assign n43540 =  ( n144 ) ? ( n17859 ) : ( n43539 ) ;
assign n43541 =  ( n142 ) ? ( n17858 ) : ( n43540 ) ;
assign n43542 =  ( n10 ) ? ( n17857 ) : ( n43541 ) ;
assign n43543 =  ( n17868 ) ? ( VREG_25_15 ) : ( n43537 ) ;
assign n43544 =  ( n17868 ) ? ( VREG_25_15 ) : ( n43542 ) ;
assign n43545 =  ( n3034 ) ? ( n43544 ) : ( VREG_25_15 ) ;
assign n43546 =  ( n2965 ) ? ( n43543 ) : ( n43545 ) ;
assign n43547 =  ( n1930 ) ? ( n43542 ) : ( n43546 ) ;
assign n43548 =  ( n879 ) ? ( n43537 ) : ( n43547 ) ;
assign n43549 =  ( n172 ) ? ( n17879 ) : ( VREG_25_15 ) ;
assign n43550 =  ( n170 ) ? ( n17878 ) : ( n43549 ) ;
assign n43551 =  ( n168 ) ? ( n17877 ) : ( n43550 ) ;
assign n43552 =  ( n166 ) ? ( n17876 ) : ( n43551 ) ;
assign n43553 =  ( n162 ) ? ( n17875 ) : ( n43552 ) ;
assign n43554 =  ( n172 ) ? ( n17889 ) : ( VREG_25_15 ) ;
assign n43555 =  ( n170 ) ? ( n17888 ) : ( n43554 ) ;
assign n43556 =  ( n168 ) ? ( n17887 ) : ( n43555 ) ;
assign n43557 =  ( n166 ) ? ( n17886 ) : ( n43556 ) ;
assign n43558 =  ( n162 ) ? ( n17885 ) : ( n43557 ) ;
assign n43559 =  ( n17868 ) ? ( VREG_25_15 ) : ( n43558 ) ;
assign n43560 =  ( n3051 ) ? ( n43559 ) : ( VREG_25_15 ) ;
assign n43561 =  ( n3040 ) ? ( n43553 ) : ( n43560 ) ;
assign n43562 =  ( n192 ) ? ( VREG_25_15 ) : ( VREG_25_15 ) ;
assign n43563 =  ( n157 ) ? ( n43561 ) : ( n43562 ) ;
assign n43564 =  ( n6 ) ? ( n43548 ) : ( n43563 ) ;
assign n43565 =  ( n571 ) ? ( n43564 ) : ( VREG_25_15 ) ;
assign n43566 =  ( n148 ) ? ( n18946 ) : ( VREG_25_2 ) ;
assign n43567 =  ( n146 ) ? ( n18945 ) : ( n43566 ) ;
assign n43568 =  ( n144 ) ? ( n18944 ) : ( n43567 ) ;
assign n43569 =  ( n142 ) ? ( n18943 ) : ( n43568 ) ;
assign n43570 =  ( n10 ) ? ( n18942 ) : ( n43569 ) ;
assign n43571 =  ( n148 ) ? ( n19980 ) : ( VREG_25_2 ) ;
assign n43572 =  ( n146 ) ? ( n19979 ) : ( n43571 ) ;
assign n43573 =  ( n144 ) ? ( n19978 ) : ( n43572 ) ;
assign n43574 =  ( n142 ) ? ( n19977 ) : ( n43573 ) ;
assign n43575 =  ( n10 ) ? ( n19976 ) : ( n43574 ) ;
assign n43576 =  ( n19987 ) ? ( VREG_25_2 ) : ( n43570 ) ;
assign n43577 =  ( n19987 ) ? ( VREG_25_2 ) : ( n43575 ) ;
assign n43578 =  ( n3034 ) ? ( n43577 ) : ( VREG_25_2 ) ;
assign n43579 =  ( n2965 ) ? ( n43576 ) : ( n43578 ) ;
assign n43580 =  ( n1930 ) ? ( n43575 ) : ( n43579 ) ;
assign n43581 =  ( n879 ) ? ( n43570 ) : ( n43580 ) ;
assign n43582 =  ( n172 ) ? ( n19998 ) : ( VREG_25_2 ) ;
assign n43583 =  ( n170 ) ? ( n19997 ) : ( n43582 ) ;
assign n43584 =  ( n168 ) ? ( n19996 ) : ( n43583 ) ;
assign n43585 =  ( n166 ) ? ( n19995 ) : ( n43584 ) ;
assign n43586 =  ( n162 ) ? ( n19994 ) : ( n43585 ) ;
assign n43587 =  ( n172 ) ? ( n20008 ) : ( VREG_25_2 ) ;
assign n43588 =  ( n170 ) ? ( n20007 ) : ( n43587 ) ;
assign n43589 =  ( n168 ) ? ( n20006 ) : ( n43588 ) ;
assign n43590 =  ( n166 ) ? ( n20005 ) : ( n43589 ) ;
assign n43591 =  ( n162 ) ? ( n20004 ) : ( n43590 ) ;
assign n43592 =  ( n19987 ) ? ( VREG_25_2 ) : ( n43591 ) ;
assign n43593 =  ( n3051 ) ? ( n43592 ) : ( VREG_25_2 ) ;
assign n43594 =  ( n3040 ) ? ( n43586 ) : ( n43593 ) ;
assign n43595 =  ( n192 ) ? ( VREG_25_2 ) : ( VREG_25_2 ) ;
assign n43596 =  ( n157 ) ? ( n43594 ) : ( n43595 ) ;
assign n43597 =  ( n6 ) ? ( n43581 ) : ( n43596 ) ;
assign n43598 =  ( n571 ) ? ( n43597 ) : ( VREG_25_2 ) ;
assign n43599 =  ( n148 ) ? ( n21065 ) : ( VREG_25_3 ) ;
assign n43600 =  ( n146 ) ? ( n21064 ) : ( n43599 ) ;
assign n43601 =  ( n144 ) ? ( n21063 ) : ( n43600 ) ;
assign n43602 =  ( n142 ) ? ( n21062 ) : ( n43601 ) ;
assign n43603 =  ( n10 ) ? ( n21061 ) : ( n43602 ) ;
assign n43604 =  ( n148 ) ? ( n22099 ) : ( VREG_25_3 ) ;
assign n43605 =  ( n146 ) ? ( n22098 ) : ( n43604 ) ;
assign n43606 =  ( n144 ) ? ( n22097 ) : ( n43605 ) ;
assign n43607 =  ( n142 ) ? ( n22096 ) : ( n43606 ) ;
assign n43608 =  ( n10 ) ? ( n22095 ) : ( n43607 ) ;
assign n43609 =  ( n22106 ) ? ( VREG_25_3 ) : ( n43603 ) ;
assign n43610 =  ( n22106 ) ? ( VREG_25_3 ) : ( n43608 ) ;
assign n43611 =  ( n3034 ) ? ( n43610 ) : ( VREG_25_3 ) ;
assign n43612 =  ( n2965 ) ? ( n43609 ) : ( n43611 ) ;
assign n43613 =  ( n1930 ) ? ( n43608 ) : ( n43612 ) ;
assign n43614 =  ( n879 ) ? ( n43603 ) : ( n43613 ) ;
assign n43615 =  ( n172 ) ? ( n22117 ) : ( VREG_25_3 ) ;
assign n43616 =  ( n170 ) ? ( n22116 ) : ( n43615 ) ;
assign n43617 =  ( n168 ) ? ( n22115 ) : ( n43616 ) ;
assign n43618 =  ( n166 ) ? ( n22114 ) : ( n43617 ) ;
assign n43619 =  ( n162 ) ? ( n22113 ) : ( n43618 ) ;
assign n43620 =  ( n172 ) ? ( n22127 ) : ( VREG_25_3 ) ;
assign n43621 =  ( n170 ) ? ( n22126 ) : ( n43620 ) ;
assign n43622 =  ( n168 ) ? ( n22125 ) : ( n43621 ) ;
assign n43623 =  ( n166 ) ? ( n22124 ) : ( n43622 ) ;
assign n43624 =  ( n162 ) ? ( n22123 ) : ( n43623 ) ;
assign n43625 =  ( n22106 ) ? ( VREG_25_3 ) : ( n43624 ) ;
assign n43626 =  ( n3051 ) ? ( n43625 ) : ( VREG_25_3 ) ;
assign n43627 =  ( n3040 ) ? ( n43619 ) : ( n43626 ) ;
assign n43628 =  ( n192 ) ? ( VREG_25_3 ) : ( VREG_25_3 ) ;
assign n43629 =  ( n157 ) ? ( n43627 ) : ( n43628 ) ;
assign n43630 =  ( n6 ) ? ( n43614 ) : ( n43629 ) ;
assign n43631 =  ( n571 ) ? ( n43630 ) : ( VREG_25_3 ) ;
assign n43632 =  ( n148 ) ? ( n23184 ) : ( VREG_25_4 ) ;
assign n43633 =  ( n146 ) ? ( n23183 ) : ( n43632 ) ;
assign n43634 =  ( n144 ) ? ( n23182 ) : ( n43633 ) ;
assign n43635 =  ( n142 ) ? ( n23181 ) : ( n43634 ) ;
assign n43636 =  ( n10 ) ? ( n23180 ) : ( n43635 ) ;
assign n43637 =  ( n148 ) ? ( n24218 ) : ( VREG_25_4 ) ;
assign n43638 =  ( n146 ) ? ( n24217 ) : ( n43637 ) ;
assign n43639 =  ( n144 ) ? ( n24216 ) : ( n43638 ) ;
assign n43640 =  ( n142 ) ? ( n24215 ) : ( n43639 ) ;
assign n43641 =  ( n10 ) ? ( n24214 ) : ( n43640 ) ;
assign n43642 =  ( n24225 ) ? ( VREG_25_4 ) : ( n43636 ) ;
assign n43643 =  ( n24225 ) ? ( VREG_25_4 ) : ( n43641 ) ;
assign n43644 =  ( n3034 ) ? ( n43643 ) : ( VREG_25_4 ) ;
assign n43645 =  ( n2965 ) ? ( n43642 ) : ( n43644 ) ;
assign n43646 =  ( n1930 ) ? ( n43641 ) : ( n43645 ) ;
assign n43647 =  ( n879 ) ? ( n43636 ) : ( n43646 ) ;
assign n43648 =  ( n172 ) ? ( n24236 ) : ( VREG_25_4 ) ;
assign n43649 =  ( n170 ) ? ( n24235 ) : ( n43648 ) ;
assign n43650 =  ( n168 ) ? ( n24234 ) : ( n43649 ) ;
assign n43651 =  ( n166 ) ? ( n24233 ) : ( n43650 ) ;
assign n43652 =  ( n162 ) ? ( n24232 ) : ( n43651 ) ;
assign n43653 =  ( n172 ) ? ( n24246 ) : ( VREG_25_4 ) ;
assign n43654 =  ( n170 ) ? ( n24245 ) : ( n43653 ) ;
assign n43655 =  ( n168 ) ? ( n24244 ) : ( n43654 ) ;
assign n43656 =  ( n166 ) ? ( n24243 ) : ( n43655 ) ;
assign n43657 =  ( n162 ) ? ( n24242 ) : ( n43656 ) ;
assign n43658 =  ( n24225 ) ? ( VREG_25_4 ) : ( n43657 ) ;
assign n43659 =  ( n3051 ) ? ( n43658 ) : ( VREG_25_4 ) ;
assign n43660 =  ( n3040 ) ? ( n43652 ) : ( n43659 ) ;
assign n43661 =  ( n192 ) ? ( VREG_25_4 ) : ( VREG_25_4 ) ;
assign n43662 =  ( n157 ) ? ( n43660 ) : ( n43661 ) ;
assign n43663 =  ( n6 ) ? ( n43647 ) : ( n43662 ) ;
assign n43664 =  ( n571 ) ? ( n43663 ) : ( VREG_25_4 ) ;
assign n43665 =  ( n148 ) ? ( n25303 ) : ( VREG_25_5 ) ;
assign n43666 =  ( n146 ) ? ( n25302 ) : ( n43665 ) ;
assign n43667 =  ( n144 ) ? ( n25301 ) : ( n43666 ) ;
assign n43668 =  ( n142 ) ? ( n25300 ) : ( n43667 ) ;
assign n43669 =  ( n10 ) ? ( n25299 ) : ( n43668 ) ;
assign n43670 =  ( n148 ) ? ( n26337 ) : ( VREG_25_5 ) ;
assign n43671 =  ( n146 ) ? ( n26336 ) : ( n43670 ) ;
assign n43672 =  ( n144 ) ? ( n26335 ) : ( n43671 ) ;
assign n43673 =  ( n142 ) ? ( n26334 ) : ( n43672 ) ;
assign n43674 =  ( n10 ) ? ( n26333 ) : ( n43673 ) ;
assign n43675 =  ( n26344 ) ? ( VREG_25_5 ) : ( n43669 ) ;
assign n43676 =  ( n26344 ) ? ( VREG_25_5 ) : ( n43674 ) ;
assign n43677 =  ( n3034 ) ? ( n43676 ) : ( VREG_25_5 ) ;
assign n43678 =  ( n2965 ) ? ( n43675 ) : ( n43677 ) ;
assign n43679 =  ( n1930 ) ? ( n43674 ) : ( n43678 ) ;
assign n43680 =  ( n879 ) ? ( n43669 ) : ( n43679 ) ;
assign n43681 =  ( n172 ) ? ( n26355 ) : ( VREG_25_5 ) ;
assign n43682 =  ( n170 ) ? ( n26354 ) : ( n43681 ) ;
assign n43683 =  ( n168 ) ? ( n26353 ) : ( n43682 ) ;
assign n43684 =  ( n166 ) ? ( n26352 ) : ( n43683 ) ;
assign n43685 =  ( n162 ) ? ( n26351 ) : ( n43684 ) ;
assign n43686 =  ( n172 ) ? ( n26365 ) : ( VREG_25_5 ) ;
assign n43687 =  ( n170 ) ? ( n26364 ) : ( n43686 ) ;
assign n43688 =  ( n168 ) ? ( n26363 ) : ( n43687 ) ;
assign n43689 =  ( n166 ) ? ( n26362 ) : ( n43688 ) ;
assign n43690 =  ( n162 ) ? ( n26361 ) : ( n43689 ) ;
assign n43691 =  ( n26344 ) ? ( VREG_25_5 ) : ( n43690 ) ;
assign n43692 =  ( n3051 ) ? ( n43691 ) : ( VREG_25_5 ) ;
assign n43693 =  ( n3040 ) ? ( n43685 ) : ( n43692 ) ;
assign n43694 =  ( n192 ) ? ( VREG_25_5 ) : ( VREG_25_5 ) ;
assign n43695 =  ( n157 ) ? ( n43693 ) : ( n43694 ) ;
assign n43696 =  ( n6 ) ? ( n43680 ) : ( n43695 ) ;
assign n43697 =  ( n571 ) ? ( n43696 ) : ( VREG_25_5 ) ;
assign n43698 =  ( n148 ) ? ( n27422 ) : ( VREG_25_6 ) ;
assign n43699 =  ( n146 ) ? ( n27421 ) : ( n43698 ) ;
assign n43700 =  ( n144 ) ? ( n27420 ) : ( n43699 ) ;
assign n43701 =  ( n142 ) ? ( n27419 ) : ( n43700 ) ;
assign n43702 =  ( n10 ) ? ( n27418 ) : ( n43701 ) ;
assign n43703 =  ( n148 ) ? ( n28456 ) : ( VREG_25_6 ) ;
assign n43704 =  ( n146 ) ? ( n28455 ) : ( n43703 ) ;
assign n43705 =  ( n144 ) ? ( n28454 ) : ( n43704 ) ;
assign n43706 =  ( n142 ) ? ( n28453 ) : ( n43705 ) ;
assign n43707 =  ( n10 ) ? ( n28452 ) : ( n43706 ) ;
assign n43708 =  ( n28463 ) ? ( VREG_25_6 ) : ( n43702 ) ;
assign n43709 =  ( n28463 ) ? ( VREG_25_6 ) : ( n43707 ) ;
assign n43710 =  ( n3034 ) ? ( n43709 ) : ( VREG_25_6 ) ;
assign n43711 =  ( n2965 ) ? ( n43708 ) : ( n43710 ) ;
assign n43712 =  ( n1930 ) ? ( n43707 ) : ( n43711 ) ;
assign n43713 =  ( n879 ) ? ( n43702 ) : ( n43712 ) ;
assign n43714 =  ( n172 ) ? ( n28474 ) : ( VREG_25_6 ) ;
assign n43715 =  ( n170 ) ? ( n28473 ) : ( n43714 ) ;
assign n43716 =  ( n168 ) ? ( n28472 ) : ( n43715 ) ;
assign n43717 =  ( n166 ) ? ( n28471 ) : ( n43716 ) ;
assign n43718 =  ( n162 ) ? ( n28470 ) : ( n43717 ) ;
assign n43719 =  ( n172 ) ? ( n28484 ) : ( VREG_25_6 ) ;
assign n43720 =  ( n170 ) ? ( n28483 ) : ( n43719 ) ;
assign n43721 =  ( n168 ) ? ( n28482 ) : ( n43720 ) ;
assign n43722 =  ( n166 ) ? ( n28481 ) : ( n43721 ) ;
assign n43723 =  ( n162 ) ? ( n28480 ) : ( n43722 ) ;
assign n43724 =  ( n28463 ) ? ( VREG_25_6 ) : ( n43723 ) ;
assign n43725 =  ( n3051 ) ? ( n43724 ) : ( VREG_25_6 ) ;
assign n43726 =  ( n3040 ) ? ( n43718 ) : ( n43725 ) ;
assign n43727 =  ( n192 ) ? ( VREG_25_6 ) : ( VREG_25_6 ) ;
assign n43728 =  ( n157 ) ? ( n43726 ) : ( n43727 ) ;
assign n43729 =  ( n6 ) ? ( n43713 ) : ( n43728 ) ;
assign n43730 =  ( n571 ) ? ( n43729 ) : ( VREG_25_6 ) ;
assign n43731 =  ( n148 ) ? ( n29541 ) : ( VREG_25_7 ) ;
assign n43732 =  ( n146 ) ? ( n29540 ) : ( n43731 ) ;
assign n43733 =  ( n144 ) ? ( n29539 ) : ( n43732 ) ;
assign n43734 =  ( n142 ) ? ( n29538 ) : ( n43733 ) ;
assign n43735 =  ( n10 ) ? ( n29537 ) : ( n43734 ) ;
assign n43736 =  ( n148 ) ? ( n30575 ) : ( VREG_25_7 ) ;
assign n43737 =  ( n146 ) ? ( n30574 ) : ( n43736 ) ;
assign n43738 =  ( n144 ) ? ( n30573 ) : ( n43737 ) ;
assign n43739 =  ( n142 ) ? ( n30572 ) : ( n43738 ) ;
assign n43740 =  ( n10 ) ? ( n30571 ) : ( n43739 ) ;
assign n43741 =  ( n30582 ) ? ( VREG_25_7 ) : ( n43735 ) ;
assign n43742 =  ( n30582 ) ? ( VREG_25_7 ) : ( n43740 ) ;
assign n43743 =  ( n3034 ) ? ( n43742 ) : ( VREG_25_7 ) ;
assign n43744 =  ( n2965 ) ? ( n43741 ) : ( n43743 ) ;
assign n43745 =  ( n1930 ) ? ( n43740 ) : ( n43744 ) ;
assign n43746 =  ( n879 ) ? ( n43735 ) : ( n43745 ) ;
assign n43747 =  ( n172 ) ? ( n30593 ) : ( VREG_25_7 ) ;
assign n43748 =  ( n170 ) ? ( n30592 ) : ( n43747 ) ;
assign n43749 =  ( n168 ) ? ( n30591 ) : ( n43748 ) ;
assign n43750 =  ( n166 ) ? ( n30590 ) : ( n43749 ) ;
assign n43751 =  ( n162 ) ? ( n30589 ) : ( n43750 ) ;
assign n43752 =  ( n172 ) ? ( n30603 ) : ( VREG_25_7 ) ;
assign n43753 =  ( n170 ) ? ( n30602 ) : ( n43752 ) ;
assign n43754 =  ( n168 ) ? ( n30601 ) : ( n43753 ) ;
assign n43755 =  ( n166 ) ? ( n30600 ) : ( n43754 ) ;
assign n43756 =  ( n162 ) ? ( n30599 ) : ( n43755 ) ;
assign n43757 =  ( n30582 ) ? ( VREG_25_7 ) : ( n43756 ) ;
assign n43758 =  ( n3051 ) ? ( n43757 ) : ( VREG_25_7 ) ;
assign n43759 =  ( n3040 ) ? ( n43751 ) : ( n43758 ) ;
assign n43760 =  ( n192 ) ? ( VREG_25_7 ) : ( VREG_25_7 ) ;
assign n43761 =  ( n157 ) ? ( n43759 ) : ( n43760 ) ;
assign n43762 =  ( n6 ) ? ( n43746 ) : ( n43761 ) ;
assign n43763 =  ( n571 ) ? ( n43762 ) : ( VREG_25_7 ) ;
assign n43764 =  ( n148 ) ? ( n31660 ) : ( VREG_25_8 ) ;
assign n43765 =  ( n146 ) ? ( n31659 ) : ( n43764 ) ;
assign n43766 =  ( n144 ) ? ( n31658 ) : ( n43765 ) ;
assign n43767 =  ( n142 ) ? ( n31657 ) : ( n43766 ) ;
assign n43768 =  ( n10 ) ? ( n31656 ) : ( n43767 ) ;
assign n43769 =  ( n148 ) ? ( n32694 ) : ( VREG_25_8 ) ;
assign n43770 =  ( n146 ) ? ( n32693 ) : ( n43769 ) ;
assign n43771 =  ( n144 ) ? ( n32692 ) : ( n43770 ) ;
assign n43772 =  ( n142 ) ? ( n32691 ) : ( n43771 ) ;
assign n43773 =  ( n10 ) ? ( n32690 ) : ( n43772 ) ;
assign n43774 =  ( n32701 ) ? ( VREG_25_8 ) : ( n43768 ) ;
assign n43775 =  ( n32701 ) ? ( VREG_25_8 ) : ( n43773 ) ;
assign n43776 =  ( n3034 ) ? ( n43775 ) : ( VREG_25_8 ) ;
assign n43777 =  ( n2965 ) ? ( n43774 ) : ( n43776 ) ;
assign n43778 =  ( n1930 ) ? ( n43773 ) : ( n43777 ) ;
assign n43779 =  ( n879 ) ? ( n43768 ) : ( n43778 ) ;
assign n43780 =  ( n172 ) ? ( n32712 ) : ( VREG_25_8 ) ;
assign n43781 =  ( n170 ) ? ( n32711 ) : ( n43780 ) ;
assign n43782 =  ( n168 ) ? ( n32710 ) : ( n43781 ) ;
assign n43783 =  ( n166 ) ? ( n32709 ) : ( n43782 ) ;
assign n43784 =  ( n162 ) ? ( n32708 ) : ( n43783 ) ;
assign n43785 =  ( n172 ) ? ( n32722 ) : ( VREG_25_8 ) ;
assign n43786 =  ( n170 ) ? ( n32721 ) : ( n43785 ) ;
assign n43787 =  ( n168 ) ? ( n32720 ) : ( n43786 ) ;
assign n43788 =  ( n166 ) ? ( n32719 ) : ( n43787 ) ;
assign n43789 =  ( n162 ) ? ( n32718 ) : ( n43788 ) ;
assign n43790 =  ( n32701 ) ? ( VREG_25_8 ) : ( n43789 ) ;
assign n43791 =  ( n3051 ) ? ( n43790 ) : ( VREG_25_8 ) ;
assign n43792 =  ( n3040 ) ? ( n43784 ) : ( n43791 ) ;
assign n43793 =  ( n192 ) ? ( VREG_25_8 ) : ( VREG_25_8 ) ;
assign n43794 =  ( n157 ) ? ( n43792 ) : ( n43793 ) ;
assign n43795 =  ( n6 ) ? ( n43779 ) : ( n43794 ) ;
assign n43796 =  ( n571 ) ? ( n43795 ) : ( VREG_25_8 ) ;
assign n43797 =  ( n148 ) ? ( n33779 ) : ( VREG_25_9 ) ;
assign n43798 =  ( n146 ) ? ( n33778 ) : ( n43797 ) ;
assign n43799 =  ( n144 ) ? ( n33777 ) : ( n43798 ) ;
assign n43800 =  ( n142 ) ? ( n33776 ) : ( n43799 ) ;
assign n43801 =  ( n10 ) ? ( n33775 ) : ( n43800 ) ;
assign n43802 =  ( n148 ) ? ( n34813 ) : ( VREG_25_9 ) ;
assign n43803 =  ( n146 ) ? ( n34812 ) : ( n43802 ) ;
assign n43804 =  ( n144 ) ? ( n34811 ) : ( n43803 ) ;
assign n43805 =  ( n142 ) ? ( n34810 ) : ( n43804 ) ;
assign n43806 =  ( n10 ) ? ( n34809 ) : ( n43805 ) ;
assign n43807 =  ( n34820 ) ? ( VREG_25_9 ) : ( n43801 ) ;
assign n43808 =  ( n34820 ) ? ( VREG_25_9 ) : ( n43806 ) ;
assign n43809 =  ( n3034 ) ? ( n43808 ) : ( VREG_25_9 ) ;
assign n43810 =  ( n2965 ) ? ( n43807 ) : ( n43809 ) ;
assign n43811 =  ( n1930 ) ? ( n43806 ) : ( n43810 ) ;
assign n43812 =  ( n879 ) ? ( n43801 ) : ( n43811 ) ;
assign n43813 =  ( n172 ) ? ( n34831 ) : ( VREG_25_9 ) ;
assign n43814 =  ( n170 ) ? ( n34830 ) : ( n43813 ) ;
assign n43815 =  ( n168 ) ? ( n34829 ) : ( n43814 ) ;
assign n43816 =  ( n166 ) ? ( n34828 ) : ( n43815 ) ;
assign n43817 =  ( n162 ) ? ( n34827 ) : ( n43816 ) ;
assign n43818 =  ( n172 ) ? ( n34841 ) : ( VREG_25_9 ) ;
assign n43819 =  ( n170 ) ? ( n34840 ) : ( n43818 ) ;
assign n43820 =  ( n168 ) ? ( n34839 ) : ( n43819 ) ;
assign n43821 =  ( n166 ) ? ( n34838 ) : ( n43820 ) ;
assign n43822 =  ( n162 ) ? ( n34837 ) : ( n43821 ) ;
assign n43823 =  ( n34820 ) ? ( VREG_25_9 ) : ( n43822 ) ;
assign n43824 =  ( n3051 ) ? ( n43823 ) : ( VREG_25_9 ) ;
assign n43825 =  ( n3040 ) ? ( n43817 ) : ( n43824 ) ;
assign n43826 =  ( n192 ) ? ( VREG_25_9 ) : ( VREG_25_9 ) ;
assign n43827 =  ( n157 ) ? ( n43825 ) : ( n43826 ) ;
assign n43828 =  ( n6 ) ? ( n43812 ) : ( n43827 ) ;
assign n43829 =  ( n571 ) ? ( n43828 ) : ( VREG_25_9 ) ;
assign n43830 =  ( n148 ) ? ( n1924 ) : ( VREG_26_0 ) ;
assign n43831 =  ( n146 ) ? ( n1923 ) : ( n43830 ) ;
assign n43832 =  ( n144 ) ? ( n1922 ) : ( n43831 ) ;
assign n43833 =  ( n142 ) ? ( n1921 ) : ( n43832 ) ;
assign n43834 =  ( n10 ) ? ( n1920 ) : ( n43833 ) ;
assign n43835 =  ( n148 ) ? ( n2959 ) : ( VREG_26_0 ) ;
assign n43836 =  ( n146 ) ? ( n2958 ) : ( n43835 ) ;
assign n43837 =  ( n144 ) ? ( n2957 ) : ( n43836 ) ;
assign n43838 =  ( n142 ) ? ( n2956 ) : ( n43837 ) ;
assign n43839 =  ( n10 ) ? ( n2955 ) : ( n43838 ) ;
assign n43840 =  ( n3032 ) ? ( VREG_26_0 ) : ( n43834 ) ;
assign n43841 =  ( n3032 ) ? ( VREG_26_0 ) : ( n43839 ) ;
assign n43842 =  ( n3034 ) ? ( n43841 ) : ( VREG_26_0 ) ;
assign n43843 =  ( n2965 ) ? ( n43840 ) : ( n43842 ) ;
assign n43844 =  ( n1930 ) ? ( n43839 ) : ( n43843 ) ;
assign n43845 =  ( n879 ) ? ( n43834 ) : ( n43844 ) ;
assign n43846 =  ( n172 ) ? ( n3045 ) : ( VREG_26_0 ) ;
assign n43847 =  ( n170 ) ? ( n3044 ) : ( n43846 ) ;
assign n43848 =  ( n168 ) ? ( n3043 ) : ( n43847 ) ;
assign n43849 =  ( n166 ) ? ( n3042 ) : ( n43848 ) ;
assign n43850 =  ( n162 ) ? ( n3041 ) : ( n43849 ) ;
assign n43851 =  ( n172 ) ? ( n3056 ) : ( VREG_26_0 ) ;
assign n43852 =  ( n170 ) ? ( n3055 ) : ( n43851 ) ;
assign n43853 =  ( n168 ) ? ( n3054 ) : ( n43852 ) ;
assign n43854 =  ( n166 ) ? ( n3053 ) : ( n43853 ) ;
assign n43855 =  ( n162 ) ? ( n3052 ) : ( n43854 ) ;
assign n43856 =  ( n3032 ) ? ( VREG_26_0 ) : ( n43855 ) ;
assign n43857 =  ( n3051 ) ? ( n43856 ) : ( VREG_26_0 ) ;
assign n43858 =  ( n3040 ) ? ( n43850 ) : ( n43857 ) ;
assign n43859 =  ( n192 ) ? ( VREG_26_0 ) : ( VREG_26_0 ) ;
assign n43860 =  ( n157 ) ? ( n43858 ) : ( n43859 ) ;
assign n43861 =  ( n6 ) ? ( n43845 ) : ( n43860 ) ;
assign n43862 =  ( n593 ) ? ( n43861 ) : ( VREG_26_0 ) ;
assign n43863 =  ( n148 ) ? ( n4113 ) : ( VREG_26_1 ) ;
assign n43864 =  ( n146 ) ? ( n4112 ) : ( n43863 ) ;
assign n43865 =  ( n144 ) ? ( n4111 ) : ( n43864 ) ;
assign n43866 =  ( n142 ) ? ( n4110 ) : ( n43865 ) ;
assign n43867 =  ( n10 ) ? ( n4109 ) : ( n43866 ) ;
assign n43868 =  ( n148 ) ? ( n5147 ) : ( VREG_26_1 ) ;
assign n43869 =  ( n146 ) ? ( n5146 ) : ( n43868 ) ;
assign n43870 =  ( n144 ) ? ( n5145 ) : ( n43869 ) ;
assign n43871 =  ( n142 ) ? ( n5144 ) : ( n43870 ) ;
assign n43872 =  ( n10 ) ? ( n5143 ) : ( n43871 ) ;
assign n43873 =  ( n5154 ) ? ( VREG_26_1 ) : ( n43867 ) ;
assign n43874 =  ( n5154 ) ? ( VREG_26_1 ) : ( n43872 ) ;
assign n43875 =  ( n3034 ) ? ( n43874 ) : ( VREG_26_1 ) ;
assign n43876 =  ( n2965 ) ? ( n43873 ) : ( n43875 ) ;
assign n43877 =  ( n1930 ) ? ( n43872 ) : ( n43876 ) ;
assign n43878 =  ( n879 ) ? ( n43867 ) : ( n43877 ) ;
assign n43879 =  ( n172 ) ? ( n5165 ) : ( VREG_26_1 ) ;
assign n43880 =  ( n170 ) ? ( n5164 ) : ( n43879 ) ;
assign n43881 =  ( n168 ) ? ( n5163 ) : ( n43880 ) ;
assign n43882 =  ( n166 ) ? ( n5162 ) : ( n43881 ) ;
assign n43883 =  ( n162 ) ? ( n5161 ) : ( n43882 ) ;
assign n43884 =  ( n172 ) ? ( n5175 ) : ( VREG_26_1 ) ;
assign n43885 =  ( n170 ) ? ( n5174 ) : ( n43884 ) ;
assign n43886 =  ( n168 ) ? ( n5173 ) : ( n43885 ) ;
assign n43887 =  ( n166 ) ? ( n5172 ) : ( n43886 ) ;
assign n43888 =  ( n162 ) ? ( n5171 ) : ( n43887 ) ;
assign n43889 =  ( n5154 ) ? ( VREG_26_1 ) : ( n43888 ) ;
assign n43890 =  ( n3051 ) ? ( n43889 ) : ( VREG_26_1 ) ;
assign n43891 =  ( n3040 ) ? ( n43883 ) : ( n43890 ) ;
assign n43892 =  ( n192 ) ? ( VREG_26_1 ) : ( VREG_26_1 ) ;
assign n43893 =  ( n157 ) ? ( n43891 ) : ( n43892 ) ;
assign n43894 =  ( n6 ) ? ( n43878 ) : ( n43893 ) ;
assign n43895 =  ( n593 ) ? ( n43894 ) : ( VREG_26_1 ) ;
assign n43896 =  ( n148 ) ? ( n6232 ) : ( VREG_26_10 ) ;
assign n43897 =  ( n146 ) ? ( n6231 ) : ( n43896 ) ;
assign n43898 =  ( n144 ) ? ( n6230 ) : ( n43897 ) ;
assign n43899 =  ( n142 ) ? ( n6229 ) : ( n43898 ) ;
assign n43900 =  ( n10 ) ? ( n6228 ) : ( n43899 ) ;
assign n43901 =  ( n148 ) ? ( n7266 ) : ( VREG_26_10 ) ;
assign n43902 =  ( n146 ) ? ( n7265 ) : ( n43901 ) ;
assign n43903 =  ( n144 ) ? ( n7264 ) : ( n43902 ) ;
assign n43904 =  ( n142 ) ? ( n7263 ) : ( n43903 ) ;
assign n43905 =  ( n10 ) ? ( n7262 ) : ( n43904 ) ;
assign n43906 =  ( n7273 ) ? ( VREG_26_10 ) : ( n43900 ) ;
assign n43907 =  ( n7273 ) ? ( VREG_26_10 ) : ( n43905 ) ;
assign n43908 =  ( n3034 ) ? ( n43907 ) : ( VREG_26_10 ) ;
assign n43909 =  ( n2965 ) ? ( n43906 ) : ( n43908 ) ;
assign n43910 =  ( n1930 ) ? ( n43905 ) : ( n43909 ) ;
assign n43911 =  ( n879 ) ? ( n43900 ) : ( n43910 ) ;
assign n43912 =  ( n172 ) ? ( n7284 ) : ( VREG_26_10 ) ;
assign n43913 =  ( n170 ) ? ( n7283 ) : ( n43912 ) ;
assign n43914 =  ( n168 ) ? ( n7282 ) : ( n43913 ) ;
assign n43915 =  ( n166 ) ? ( n7281 ) : ( n43914 ) ;
assign n43916 =  ( n162 ) ? ( n7280 ) : ( n43915 ) ;
assign n43917 =  ( n172 ) ? ( n7294 ) : ( VREG_26_10 ) ;
assign n43918 =  ( n170 ) ? ( n7293 ) : ( n43917 ) ;
assign n43919 =  ( n168 ) ? ( n7292 ) : ( n43918 ) ;
assign n43920 =  ( n166 ) ? ( n7291 ) : ( n43919 ) ;
assign n43921 =  ( n162 ) ? ( n7290 ) : ( n43920 ) ;
assign n43922 =  ( n7273 ) ? ( VREG_26_10 ) : ( n43921 ) ;
assign n43923 =  ( n3051 ) ? ( n43922 ) : ( VREG_26_10 ) ;
assign n43924 =  ( n3040 ) ? ( n43916 ) : ( n43923 ) ;
assign n43925 =  ( n192 ) ? ( VREG_26_10 ) : ( VREG_26_10 ) ;
assign n43926 =  ( n157 ) ? ( n43924 ) : ( n43925 ) ;
assign n43927 =  ( n6 ) ? ( n43911 ) : ( n43926 ) ;
assign n43928 =  ( n593 ) ? ( n43927 ) : ( VREG_26_10 ) ;
assign n43929 =  ( n148 ) ? ( n8351 ) : ( VREG_26_11 ) ;
assign n43930 =  ( n146 ) ? ( n8350 ) : ( n43929 ) ;
assign n43931 =  ( n144 ) ? ( n8349 ) : ( n43930 ) ;
assign n43932 =  ( n142 ) ? ( n8348 ) : ( n43931 ) ;
assign n43933 =  ( n10 ) ? ( n8347 ) : ( n43932 ) ;
assign n43934 =  ( n148 ) ? ( n9385 ) : ( VREG_26_11 ) ;
assign n43935 =  ( n146 ) ? ( n9384 ) : ( n43934 ) ;
assign n43936 =  ( n144 ) ? ( n9383 ) : ( n43935 ) ;
assign n43937 =  ( n142 ) ? ( n9382 ) : ( n43936 ) ;
assign n43938 =  ( n10 ) ? ( n9381 ) : ( n43937 ) ;
assign n43939 =  ( n9392 ) ? ( VREG_26_11 ) : ( n43933 ) ;
assign n43940 =  ( n9392 ) ? ( VREG_26_11 ) : ( n43938 ) ;
assign n43941 =  ( n3034 ) ? ( n43940 ) : ( VREG_26_11 ) ;
assign n43942 =  ( n2965 ) ? ( n43939 ) : ( n43941 ) ;
assign n43943 =  ( n1930 ) ? ( n43938 ) : ( n43942 ) ;
assign n43944 =  ( n879 ) ? ( n43933 ) : ( n43943 ) ;
assign n43945 =  ( n172 ) ? ( n9403 ) : ( VREG_26_11 ) ;
assign n43946 =  ( n170 ) ? ( n9402 ) : ( n43945 ) ;
assign n43947 =  ( n168 ) ? ( n9401 ) : ( n43946 ) ;
assign n43948 =  ( n166 ) ? ( n9400 ) : ( n43947 ) ;
assign n43949 =  ( n162 ) ? ( n9399 ) : ( n43948 ) ;
assign n43950 =  ( n172 ) ? ( n9413 ) : ( VREG_26_11 ) ;
assign n43951 =  ( n170 ) ? ( n9412 ) : ( n43950 ) ;
assign n43952 =  ( n168 ) ? ( n9411 ) : ( n43951 ) ;
assign n43953 =  ( n166 ) ? ( n9410 ) : ( n43952 ) ;
assign n43954 =  ( n162 ) ? ( n9409 ) : ( n43953 ) ;
assign n43955 =  ( n9392 ) ? ( VREG_26_11 ) : ( n43954 ) ;
assign n43956 =  ( n3051 ) ? ( n43955 ) : ( VREG_26_11 ) ;
assign n43957 =  ( n3040 ) ? ( n43949 ) : ( n43956 ) ;
assign n43958 =  ( n192 ) ? ( VREG_26_11 ) : ( VREG_26_11 ) ;
assign n43959 =  ( n157 ) ? ( n43957 ) : ( n43958 ) ;
assign n43960 =  ( n6 ) ? ( n43944 ) : ( n43959 ) ;
assign n43961 =  ( n593 ) ? ( n43960 ) : ( VREG_26_11 ) ;
assign n43962 =  ( n148 ) ? ( n10470 ) : ( VREG_26_12 ) ;
assign n43963 =  ( n146 ) ? ( n10469 ) : ( n43962 ) ;
assign n43964 =  ( n144 ) ? ( n10468 ) : ( n43963 ) ;
assign n43965 =  ( n142 ) ? ( n10467 ) : ( n43964 ) ;
assign n43966 =  ( n10 ) ? ( n10466 ) : ( n43965 ) ;
assign n43967 =  ( n148 ) ? ( n11504 ) : ( VREG_26_12 ) ;
assign n43968 =  ( n146 ) ? ( n11503 ) : ( n43967 ) ;
assign n43969 =  ( n144 ) ? ( n11502 ) : ( n43968 ) ;
assign n43970 =  ( n142 ) ? ( n11501 ) : ( n43969 ) ;
assign n43971 =  ( n10 ) ? ( n11500 ) : ( n43970 ) ;
assign n43972 =  ( n11511 ) ? ( VREG_26_12 ) : ( n43966 ) ;
assign n43973 =  ( n11511 ) ? ( VREG_26_12 ) : ( n43971 ) ;
assign n43974 =  ( n3034 ) ? ( n43973 ) : ( VREG_26_12 ) ;
assign n43975 =  ( n2965 ) ? ( n43972 ) : ( n43974 ) ;
assign n43976 =  ( n1930 ) ? ( n43971 ) : ( n43975 ) ;
assign n43977 =  ( n879 ) ? ( n43966 ) : ( n43976 ) ;
assign n43978 =  ( n172 ) ? ( n11522 ) : ( VREG_26_12 ) ;
assign n43979 =  ( n170 ) ? ( n11521 ) : ( n43978 ) ;
assign n43980 =  ( n168 ) ? ( n11520 ) : ( n43979 ) ;
assign n43981 =  ( n166 ) ? ( n11519 ) : ( n43980 ) ;
assign n43982 =  ( n162 ) ? ( n11518 ) : ( n43981 ) ;
assign n43983 =  ( n172 ) ? ( n11532 ) : ( VREG_26_12 ) ;
assign n43984 =  ( n170 ) ? ( n11531 ) : ( n43983 ) ;
assign n43985 =  ( n168 ) ? ( n11530 ) : ( n43984 ) ;
assign n43986 =  ( n166 ) ? ( n11529 ) : ( n43985 ) ;
assign n43987 =  ( n162 ) ? ( n11528 ) : ( n43986 ) ;
assign n43988 =  ( n11511 ) ? ( VREG_26_12 ) : ( n43987 ) ;
assign n43989 =  ( n3051 ) ? ( n43988 ) : ( VREG_26_12 ) ;
assign n43990 =  ( n3040 ) ? ( n43982 ) : ( n43989 ) ;
assign n43991 =  ( n192 ) ? ( VREG_26_12 ) : ( VREG_26_12 ) ;
assign n43992 =  ( n157 ) ? ( n43990 ) : ( n43991 ) ;
assign n43993 =  ( n6 ) ? ( n43977 ) : ( n43992 ) ;
assign n43994 =  ( n593 ) ? ( n43993 ) : ( VREG_26_12 ) ;
assign n43995 =  ( n148 ) ? ( n12589 ) : ( VREG_26_13 ) ;
assign n43996 =  ( n146 ) ? ( n12588 ) : ( n43995 ) ;
assign n43997 =  ( n144 ) ? ( n12587 ) : ( n43996 ) ;
assign n43998 =  ( n142 ) ? ( n12586 ) : ( n43997 ) ;
assign n43999 =  ( n10 ) ? ( n12585 ) : ( n43998 ) ;
assign n44000 =  ( n148 ) ? ( n13623 ) : ( VREG_26_13 ) ;
assign n44001 =  ( n146 ) ? ( n13622 ) : ( n44000 ) ;
assign n44002 =  ( n144 ) ? ( n13621 ) : ( n44001 ) ;
assign n44003 =  ( n142 ) ? ( n13620 ) : ( n44002 ) ;
assign n44004 =  ( n10 ) ? ( n13619 ) : ( n44003 ) ;
assign n44005 =  ( n13630 ) ? ( VREG_26_13 ) : ( n43999 ) ;
assign n44006 =  ( n13630 ) ? ( VREG_26_13 ) : ( n44004 ) ;
assign n44007 =  ( n3034 ) ? ( n44006 ) : ( VREG_26_13 ) ;
assign n44008 =  ( n2965 ) ? ( n44005 ) : ( n44007 ) ;
assign n44009 =  ( n1930 ) ? ( n44004 ) : ( n44008 ) ;
assign n44010 =  ( n879 ) ? ( n43999 ) : ( n44009 ) ;
assign n44011 =  ( n172 ) ? ( n13641 ) : ( VREG_26_13 ) ;
assign n44012 =  ( n170 ) ? ( n13640 ) : ( n44011 ) ;
assign n44013 =  ( n168 ) ? ( n13639 ) : ( n44012 ) ;
assign n44014 =  ( n166 ) ? ( n13638 ) : ( n44013 ) ;
assign n44015 =  ( n162 ) ? ( n13637 ) : ( n44014 ) ;
assign n44016 =  ( n172 ) ? ( n13651 ) : ( VREG_26_13 ) ;
assign n44017 =  ( n170 ) ? ( n13650 ) : ( n44016 ) ;
assign n44018 =  ( n168 ) ? ( n13649 ) : ( n44017 ) ;
assign n44019 =  ( n166 ) ? ( n13648 ) : ( n44018 ) ;
assign n44020 =  ( n162 ) ? ( n13647 ) : ( n44019 ) ;
assign n44021 =  ( n13630 ) ? ( VREG_26_13 ) : ( n44020 ) ;
assign n44022 =  ( n3051 ) ? ( n44021 ) : ( VREG_26_13 ) ;
assign n44023 =  ( n3040 ) ? ( n44015 ) : ( n44022 ) ;
assign n44024 =  ( n192 ) ? ( VREG_26_13 ) : ( VREG_26_13 ) ;
assign n44025 =  ( n157 ) ? ( n44023 ) : ( n44024 ) ;
assign n44026 =  ( n6 ) ? ( n44010 ) : ( n44025 ) ;
assign n44027 =  ( n593 ) ? ( n44026 ) : ( VREG_26_13 ) ;
assign n44028 =  ( n148 ) ? ( n14708 ) : ( VREG_26_14 ) ;
assign n44029 =  ( n146 ) ? ( n14707 ) : ( n44028 ) ;
assign n44030 =  ( n144 ) ? ( n14706 ) : ( n44029 ) ;
assign n44031 =  ( n142 ) ? ( n14705 ) : ( n44030 ) ;
assign n44032 =  ( n10 ) ? ( n14704 ) : ( n44031 ) ;
assign n44033 =  ( n148 ) ? ( n15742 ) : ( VREG_26_14 ) ;
assign n44034 =  ( n146 ) ? ( n15741 ) : ( n44033 ) ;
assign n44035 =  ( n144 ) ? ( n15740 ) : ( n44034 ) ;
assign n44036 =  ( n142 ) ? ( n15739 ) : ( n44035 ) ;
assign n44037 =  ( n10 ) ? ( n15738 ) : ( n44036 ) ;
assign n44038 =  ( n15749 ) ? ( VREG_26_14 ) : ( n44032 ) ;
assign n44039 =  ( n15749 ) ? ( VREG_26_14 ) : ( n44037 ) ;
assign n44040 =  ( n3034 ) ? ( n44039 ) : ( VREG_26_14 ) ;
assign n44041 =  ( n2965 ) ? ( n44038 ) : ( n44040 ) ;
assign n44042 =  ( n1930 ) ? ( n44037 ) : ( n44041 ) ;
assign n44043 =  ( n879 ) ? ( n44032 ) : ( n44042 ) ;
assign n44044 =  ( n172 ) ? ( n15760 ) : ( VREG_26_14 ) ;
assign n44045 =  ( n170 ) ? ( n15759 ) : ( n44044 ) ;
assign n44046 =  ( n168 ) ? ( n15758 ) : ( n44045 ) ;
assign n44047 =  ( n166 ) ? ( n15757 ) : ( n44046 ) ;
assign n44048 =  ( n162 ) ? ( n15756 ) : ( n44047 ) ;
assign n44049 =  ( n172 ) ? ( n15770 ) : ( VREG_26_14 ) ;
assign n44050 =  ( n170 ) ? ( n15769 ) : ( n44049 ) ;
assign n44051 =  ( n168 ) ? ( n15768 ) : ( n44050 ) ;
assign n44052 =  ( n166 ) ? ( n15767 ) : ( n44051 ) ;
assign n44053 =  ( n162 ) ? ( n15766 ) : ( n44052 ) ;
assign n44054 =  ( n15749 ) ? ( VREG_26_14 ) : ( n44053 ) ;
assign n44055 =  ( n3051 ) ? ( n44054 ) : ( VREG_26_14 ) ;
assign n44056 =  ( n3040 ) ? ( n44048 ) : ( n44055 ) ;
assign n44057 =  ( n192 ) ? ( VREG_26_14 ) : ( VREG_26_14 ) ;
assign n44058 =  ( n157 ) ? ( n44056 ) : ( n44057 ) ;
assign n44059 =  ( n6 ) ? ( n44043 ) : ( n44058 ) ;
assign n44060 =  ( n593 ) ? ( n44059 ) : ( VREG_26_14 ) ;
assign n44061 =  ( n148 ) ? ( n16827 ) : ( VREG_26_15 ) ;
assign n44062 =  ( n146 ) ? ( n16826 ) : ( n44061 ) ;
assign n44063 =  ( n144 ) ? ( n16825 ) : ( n44062 ) ;
assign n44064 =  ( n142 ) ? ( n16824 ) : ( n44063 ) ;
assign n44065 =  ( n10 ) ? ( n16823 ) : ( n44064 ) ;
assign n44066 =  ( n148 ) ? ( n17861 ) : ( VREG_26_15 ) ;
assign n44067 =  ( n146 ) ? ( n17860 ) : ( n44066 ) ;
assign n44068 =  ( n144 ) ? ( n17859 ) : ( n44067 ) ;
assign n44069 =  ( n142 ) ? ( n17858 ) : ( n44068 ) ;
assign n44070 =  ( n10 ) ? ( n17857 ) : ( n44069 ) ;
assign n44071 =  ( n17868 ) ? ( VREG_26_15 ) : ( n44065 ) ;
assign n44072 =  ( n17868 ) ? ( VREG_26_15 ) : ( n44070 ) ;
assign n44073 =  ( n3034 ) ? ( n44072 ) : ( VREG_26_15 ) ;
assign n44074 =  ( n2965 ) ? ( n44071 ) : ( n44073 ) ;
assign n44075 =  ( n1930 ) ? ( n44070 ) : ( n44074 ) ;
assign n44076 =  ( n879 ) ? ( n44065 ) : ( n44075 ) ;
assign n44077 =  ( n172 ) ? ( n17879 ) : ( VREG_26_15 ) ;
assign n44078 =  ( n170 ) ? ( n17878 ) : ( n44077 ) ;
assign n44079 =  ( n168 ) ? ( n17877 ) : ( n44078 ) ;
assign n44080 =  ( n166 ) ? ( n17876 ) : ( n44079 ) ;
assign n44081 =  ( n162 ) ? ( n17875 ) : ( n44080 ) ;
assign n44082 =  ( n172 ) ? ( n17889 ) : ( VREG_26_15 ) ;
assign n44083 =  ( n170 ) ? ( n17888 ) : ( n44082 ) ;
assign n44084 =  ( n168 ) ? ( n17887 ) : ( n44083 ) ;
assign n44085 =  ( n166 ) ? ( n17886 ) : ( n44084 ) ;
assign n44086 =  ( n162 ) ? ( n17885 ) : ( n44085 ) ;
assign n44087 =  ( n17868 ) ? ( VREG_26_15 ) : ( n44086 ) ;
assign n44088 =  ( n3051 ) ? ( n44087 ) : ( VREG_26_15 ) ;
assign n44089 =  ( n3040 ) ? ( n44081 ) : ( n44088 ) ;
assign n44090 =  ( n192 ) ? ( VREG_26_15 ) : ( VREG_26_15 ) ;
assign n44091 =  ( n157 ) ? ( n44089 ) : ( n44090 ) ;
assign n44092 =  ( n6 ) ? ( n44076 ) : ( n44091 ) ;
assign n44093 =  ( n593 ) ? ( n44092 ) : ( VREG_26_15 ) ;
assign n44094 =  ( n148 ) ? ( n18946 ) : ( VREG_26_2 ) ;
assign n44095 =  ( n146 ) ? ( n18945 ) : ( n44094 ) ;
assign n44096 =  ( n144 ) ? ( n18944 ) : ( n44095 ) ;
assign n44097 =  ( n142 ) ? ( n18943 ) : ( n44096 ) ;
assign n44098 =  ( n10 ) ? ( n18942 ) : ( n44097 ) ;
assign n44099 =  ( n148 ) ? ( n19980 ) : ( VREG_26_2 ) ;
assign n44100 =  ( n146 ) ? ( n19979 ) : ( n44099 ) ;
assign n44101 =  ( n144 ) ? ( n19978 ) : ( n44100 ) ;
assign n44102 =  ( n142 ) ? ( n19977 ) : ( n44101 ) ;
assign n44103 =  ( n10 ) ? ( n19976 ) : ( n44102 ) ;
assign n44104 =  ( n19987 ) ? ( VREG_26_2 ) : ( n44098 ) ;
assign n44105 =  ( n19987 ) ? ( VREG_26_2 ) : ( n44103 ) ;
assign n44106 =  ( n3034 ) ? ( n44105 ) : ( VREG_26_2 ) ;
assign n44107 =  ( n2965 ) ? ( n44104 ) : ( n44106 ) ;
assign n44108 =  ( n1930 ) ? ( n44103 ) : ( n44107 ) ;
assign n44109 =  ( n879 ) ? ( n44098 ) : ( n44108 ) ;
assign n44110 =  ( n172 ) ? ( n19998 ) : ( VREG_26_2 ) ;
assign n44111 =  ( n170 ) ? ( n19997 ) : ( n44110 ) ;
assign n44112 =  ( n168 ) ? ( n19996 ) : ( n44111 ) ;
assign n44113 =  ( n166 ) ? ( n19995 ) : ( n44112 ) ;
assign n44114 =  ( n162 ) ? ( n19994 ) : ( n44113 ) ;
assign n44115 =  ( n172 ) ? ( n20008 ) : ( VREG_26_2 ) ;
assign n44116 =  ( n170 ) ? ( n20007 ) : ( n44115 ) ;
assign n44117 =  ( n168 ) ? ( n20006 ) : ( n44116 ) ;
assign n44118 =  ( n166 ) ? ( n20005 ) : ( n44117 ) ;
assign n44119 =  ( n162 ) ? ( n20004 ) : ( n44118 ) ;
assign n44120 =  ( n19987 ) ? ( VREG_26_2 ) : ( n44119 ) ;
assign n44121 =  ( n3051 ) ? ( n44120 ) : ( VREG_26_2 ) ;
assign n44122 =  ( n3040 ) ? ( n44114 ) : ( n44121 ) ;
assign n44123 =  ( n192 ) ? ( VREG_26_2 ) : ( VREG_26_2 ) ;
assign n44124 =  ( n157 ) ? ( n44122 ) : ( n44123 ) ;
assign n44125 =  ( n6 ) ? ( n44109 ) : ( n44124 ) ;
assign n44126 =  ( n593 ) ? ( n44125 ) : ( VREG_26_2 ) ;
assign n44127 =  ( n148 ) ? ( n21065 ) : ( VREG_26_3 ) ;
assign n44128 =  ( n146 ) ? ( n21064 ) : ( n44127 ) ;
assign n44129 =  ( n144 ) ? ( n21063 ) : ( n44128 ) ;
assign n44130 =  ( n142 ) ? ( n21062 ) : ( n44129 ) ;
assign n44131 =  ( n10 ) ? ( n21061 ) : ( n44130 ) ;
assign n44132 =  ( n148 ) ? ( n22099 ) : ( VREG_26_3 ) ;
assign n44133 =  ( n146 ) ? ( n22098 ) : ( n44132 ) ;
assign n44134 =  ( n144 ) ? ( n22097 ) : ( n44133 ) ;
assign n44135 =  ( n142 ) ? ( n22096 ) : ( n44134 ) ;
assign n44136 =  ( n10 ) ? ( n22095 ) : ( n44135 ) ;
assign n44137 =  ( n22106 ) ? ( VREG_26_3 ) : ( n44131 ) ;
assign n44138 =  ( n22106 ) ? ( VREG_26_3 ) : ( n44136 ) ;
assign n44139 =  ( n3034 ) ? ( n44138 ) : ( VREG_26_3 ) ;
assign n44140 =  ( n2965 ) ? ( n44137 ) : ( n44139 ) ;
assign n44141 =  ( n1930 ) ? ( n44136 ) : ( n44140 ) ;
assign n44142 =  ( n879 ) ? ( n44131 ) : ( n44141 ) ;
assign n44143 =  ( n172 ) ? ( n22117 ) : ( VREG_26_3 ) ;
assign n44144 =  ( n170 ) ? ( n22116 ) : ( n44143 ) ;
assign n44145 =  ( n168 ) ? ( n22115 ) : ( n44144 ) ;
assign n44146 =  ( n166 ) ? ( n22114 ) : ( n44145 ) ;
assign n44147 =  ( n162 ) ? ( n22113 ) : ( n44146 ) ;
assign n44148 =  ( n172 ) ? ( n22127 ) : ( VREG_26_3 ) ;
assign n44149 =  ( n170 ) ? ( n22126 ) : ( n44148 ) ;
assign n44150 =  ( n168 ) ? ( n22125 ) : ( n44149 ) ;
assign n44151 =  ( n166 ) ? ( n22124 ) : ( n44150 ) ;
assign n44152 =  ( n162 ) ? ( n22123 ) : ( n44151 ) ;
assign n44153 =  ( n22106 ) ? ( VREG_26_3 ) : ( n44152 ) ;
assign n44154 =  ( n3051 ) ? ( n44153 ) : ( VREG_26_3 ) ;
assign n44155 =  ( n3040 ) ? ( n44147 ) : ( n44154 ) ;
assign n44156 =  ( n192 ) ? ( VREG_26_3 ) : ( VREG_26_3 ) ;
assign n44157 =  ( n157 ) ? ( n44155 ) : ( n44156 ) ;
assign n44158 =  ( n6 ) ? ( n44142 ) : ( n44157 ) ;
assign n44159 =  ( n593 ) ? ( n44158 ) : ( VREG_26_3 ) ;
assign n44160 =  ( n148 ) ? ( n23184 ) : ( VREG_26_4 ) ;
assign n44161 =  ( n146 ) ? ( n23183 ) : ( n44160 ) ;
assign n44162 =  ( n144 ) ? ( n23182 ) : ( n44161 ) ;
assign n44163 =  ( n142 ) ? ( n23181 ) : ( n44162 ) ;
assign n44164 =  ( n10 ) ? ( n23180 ) : ( n44163 ) ;
assign n44165 =  ( n148 ) ? ( n24218 ) : ( VREG_26_4 ) ;
assign n44166 =  ( n146 ) ? ( n24217 ) : ( n44165 ) ;
assign n44167 =  ( n144 ) ? ( n24216 ) : ( n44166 ) ;
assign n44168 =  ( n142 ) ? ( n24215 ) : ( n44167 ) ;
assign n44169 =  ( n10 ) ? ( n24214 ) : ( n44168 ) ;
assign n44170 =  ( n24225 ) ? ( VREG_26_4 ) : ( n44164 ) ;
assign n44171 =  ( n24225 ) ? ( VREG_26_4 ) : ( n44169 ) ;
assign n44172 =  ( n3034 ) ? ( n44171 ) : ( VREG_26_4 ) ;
assign n44173 =  ( n2965 ) ? ( n44170 ) : ( n44172 ) ;
assign n44174 =  ( n1930 ) ? ( n44169 ) : ( n44173 ) ;
assign n44175 =  ( n879 ) ? ( n44164 ) : ( n44174 ) ;
assign n44176 =  ( n172 ) ? ( n24236 ) : ( VREG_26_4 ) ;
assign n44177 =  ( n170 ) ? ( n24235 ) : ( n44176 ) ;
assign n44178 =  ( n168 ) ? ( n24234 ) : ( n44177 ) ;
assign n44179 =  ( n166 ) ? ( n24233 ) : ( n44178 ) ;
assign n44180 =  ( n162 ) ? ( n24232 ) : ( n44179 ) ;
assign n44181 =  ( n172 ) ? ( n24246 ) : ( VREG_26_4 ) ;
assign n44182 =  ( n170 ) ? ( n24245 ) : ( n44181 ) ;
assign n44183 =  ( n168 ) ? ( n24244 ) : ( n44182 ) ;
assign n44184 =  ( n166 ) ? ( n24243 ) : ( n44183 ) ;
assign n44185 =  ( n162 ) ? ( n24242 ) : ( n44184 ) ;
assign n44186 =  ( n24225 ) ? ( VREG_26_4 ) : ( n44185 ) ;
assign n44187 =  ( n3051 ) ? ( n44186 ) : ( VREG_26_4 ) ;
assign n44188 =  ( n3040 ) ? ( n44180 ) : ( n44187 ) ;
assign n44189 =  ( n192 ) ? ( VREG_26_4 ) : ( VREG_26_4 ) ;
assign n44190 =  ( n157 ) ? ( n44188 ) : ( n44189 ) ;
assign n44191 =  ( n6 ) ? ( n44175 ) : ( n44190 ) ;
assign n44192 =  ( n593 ) ? ( n44191 ) : ( VREG_26_4 ) ;
assign n44193 =  ( n148 ) ? ( n25303 ) : ( VREG_26_5 ) ;
assign n44194 =  ( n146 ) ? ( n25302 ) : ( n44193 ) ;
assign n44195 =  ( n144 ) ? ( n25301 ) : ( n44194 ) ;
assign n44196 =  ( n142 ) ? ( n25300 ) : ( n44195 ) ;
assign n44197 =  ( n10 ) ? ( n25299 ) : ( n44196 ) ;
assign n44198 =  ( n148 ) ? ( n26337 ) : ( VREG_26_5 ) ;
assign n44199 =  ( n146 ) ? ( n26336 ) : ( n44198 ) ;
assign n44200 =  ( n144 ) ? ( n26335 ) : ( n44199 ) ;
assign n44201 =  ( n142 ) ? ( n26334 ) : ( n44200 ) ;
assign n44202 =  ( n10 ) ? ( n26333 ) : ( n44201 ) ;
assign n44203 =  ( n26344 ) ? ( VREG_26_5 ) : ( n44197 ) ;
assign n44204 =  ( n26344 ) ? ( VREG_26_5 ) : ( n44202 ) ;
assign n44205 =  ( n3034 ) ? ( n44204 ) : ( VREG_26_5 ) ;
assign n44206 =  ( n2965 ) ? ( n44203 ) : ( n44205 ) ;
assign n44207 =  ( n1930 ) ? ( n44202 ) : ( n44206 ) ;
assign n44208 =  ( n879 ) ? ( n44197 ) : ( n44207 ) ;
assign n44209 =  ( n172 ) ? ( n26355 ) : ( VREG_26_5 ) ;
assign n44210 =  ( n170 ) ? ( n26354 ) : ( n44209 ) ;
assign n44211 =  ( n168 ) ? ( n26353 ) : ( n44210 ) ;
assign n44212 =  ( n166 ) ? ( n26352 ) : ( n44211 ) ;
assign n44213 =  ( n162 ) ? ( n26351 ) : ( n44212 ) ;
assign n44214 =  ( n172 ) ? ( n26365 ) : ( VREG_26_5 ) ;
assign n44215 =  ( n170 ) ? ( n26364 ) : ( n44214 ) ;
assign n44216 =  ( n168 ) ? ( n26363 ) : ( n44215 ) ;
assign n44217 =  ( n166 ) ? ( n26362 ) : ( n44216 ) ;
assign n44218 =  ( n162 ) ? ( n26361 ) : ( n44217 ) ;
assign n44219 =  ( n26344 ) ? ( VREG_26_5 ) : ( n44218 ) ;
assign n44220 =  ( n3051 ) ? ( n44219 ) : ( VREG_26_5 ) ;
assign n44221 =  ( n3040 ) ? ( n44213 ) : ( n44220 ) ;
assign n44222 =  ( n192 ) ? ( VREG_26_5 ) : ( VREG_26_5 ) ;
assign n44223 =  ( n157 ) ? ( n44221 ) : ( n44222 ) ;
assign n44224 =  ( n6 ) ? ( n44208 ) : ( n44223 ) ;
assign n44225 =  ( n593 ) ? ( n44224 ) : ( VREG_26_5 ) ;
assign n44226 =  ( n148 ) ? ( n27422 ) : ( VREG_26_6 ) ;
assign n44227 =  ( n146 ) ? ( n27421 ) : ( n44226 ) ;
assign n44228 =  ( n144 ) ? ( n27420 ) : ( n44227 ) ;
assign n44229 =  ( n142 ) ? ( n27419 ) : ( n44228 ) ;
assign n44230 =  ( n10 ) ? ( n27418 ) : ( n44229 ) ;
assign n44231 =  ( n148 ) ? ( n28456 ) : ( VREG_26_6 ) ;
assign n44232 =  ( n146 ) ? ( n28455 ) : ( n44231 ) ;
assign n44233 =  ( n144 ) ? ( n28454 ) : ( n44232 ) ;
assign n44234 =  ( n142 ) ? ( n28453 ) : ( n44233 ) ;
assign n44235 =  ( n10 ) ? ( n28452 ) : ( n44234 ) ;
assign n44236 =  ( n28463 ) ? ( VREG_26_6 ) : ( n44230 ) ;
assign n44237 =  ( n28463 ) ? ( VREG_26_6 ) : ( n44235 ) ;
assign n44238 =  ( n3034 ) ? ( n44237 ) : ( VREG_26_6 ) ;
assign n44239 =  ( n2965 ) ? ( n44236 ) : ( n44238 ) ;
assign n44240 =  ( n1930 ) ? ( n44235 ) : ( n44239 ) ;
assign n44241 =  ( n879 ) ? ( n44230 ) : ( n44240 ) ;
assign n44242 =  ( n172 ) ? ( n28474 ) : ( VREG_26_6 ) ;
assign n44243 =  ( n170 ) ? ( n28473 ) : ( n44242 ) ;
assign n44244 =  ( n168 ) ? ( n28472 ) : ( n44243 ) ;
assign n44245 =  ( n166 ) ? ( n28471 ) : ( n44244 ) ;
assign n44246 =  ( n162 ) ? ( n28470 ) : ( n44245 ) ;
assign n44247 =  ( n172 ) ? ( n28484 ) : ( VREG_26_6 ) ;
assign n44248 =  ( n170 ) ? ( n28483 ) : ( n44247 ) ;
assign n44249 =  ( n168 ) ? ( n28482 ) : ( n44248 ) ;
assign n44250 =  ( n166 ) ? ( n28481 ) : ( n44249 ) ;
assign n44251 =  ( n162 ) ? ( n28480 ) : ( n44250 ) ;
assign n44252 =  ( n28463 ) ? ( VREG_26_6 ) : ( n44251 ) ;
assign n44253 =  ( n3051 ) ? ( n44252 ) : ( VREG_26_6 ) ;
assign n44254 =  ( n3040 ) ? ( n44246 ) : ( n44253 ) ;
assign n44255 =  ( n192 ) ? ( VREG_26_6 ) : ( VREG_26_6 ) ;
assign n44256 =  ( n157 ) ? ( n44254 ) : ( n44255 ) ;
assign n44257 =  ( n6 ) ? ( n44241 ) : ( n44256 ) ;
assign n44258 =  ( n593 ) ? ( n44257 ) : ( VREG_26_6 ) ;
assign n44259 =  ( n148 ) ? ( n29541 ) : ( VREG_26_7 ) ;
assign n44260 =  ( n146 ) ? ( n29540 ) : ( n44259 ) ;
assign n44261 =  ( n144 ) ? ( n29539 ) : ( n44260 ) ;
assign n44262 =  ( n142 ) ? ( n29538 ) : ( n44261 ) ;
assign n44263 =  ( n10 ) ? ( n29537 ) : ( n44262 ) ;
assign n44264 =  ( n148 ) ? ( n30575 ) : ( VREG_26_7 ) ;
assign n44265 =  ( n146 ) ? ( n30574 ) : ( n44264 ) ;
assign n44266 =  ( n144 ) ? ( n30573 ) : ( n44265 ) ;
assign n44267 =  ( n142 ) ? ( n30572 ) : ( n44266 ) ;
assign n44268 =  ( n10 ) ? ( n30571 ) : ( n44267 ) ;
assign n44269 =  ( n30582 ) ? ( VREG_26_7 ) : ( n44263 ) ;
assign n44270 =  ( n30582 ) ? ( VREG_26_7 ) : ( n44268 ) ;
assign n44271 =  ( n3034 ) ? ( n44270 ) : ( VREG_26_7 ) ;
assign n44272 =  ( n2965 ) ? ( n44269 ) : ( n44271 ) ;
assign n44273 =  ( n1930 ) ? ( n44268 ) : ( n44272 ) ;
assign n44274 =  ( n879 ) ? ( n44263 ) : ( n44273 ) ;
assign n44275 =  ( n172 ) ? ( n30593 ) : ( VREG_26_7 ) ;
assign n44276 =  ( n170 ) ? ( n30592 ) : ( n44275 ) ;
assign n44277 =  ( n168 ) ? ( n30591 ) : ( n44276 ) ;
assign n44278 =  ( n166 ) ? ( n30590 ) : ( n44277 ) ;
assign n44279 =  ( n162 ) ? ( n30589 ) : ( n44278 ) ;
assign n44280 =  ( n172 ) ? ( n30603 ) : ( VREG_26_7 ) ;
assign n44281 =  ( n170 ) ? ( n30602 ) : ( n44280 ) ;
assign n44282 =  ( n168 ) ? ( n30601 ) : ( n44281 ) ;
assign n44283 =  ( n166 ) ? ( n30600 ) : ( n44282 ) ;
assign n44284 =  ( n162 ) ? ( n30599 ) : ( n44283 ) ;
assign n44285 =  ( n30582 ) ? ( VREG_26_7 ) : ( n44284 ) ;
assign n44286 =  ( n3051 ) ? ( n44285 ) : ( VREG_26_7 ) ;
assign n44287 =  ( n3040 ) ? ( n44279 ) : ( n44286 ) ;
assign n44288 =  ( n192 ) ? ( VREG_26_7 ) : ( VREG_26_7 ) ;
assign n44289 =  ( n157 ) ? ( n44287 ) : ( n44288 ) ;
assign n44290 =  ( n6 ) ? ( n44274 ) : ( n44289 ) ;
assign n44291 =  ( n593 ) ? ( n44290 ) : ( VREG_26_7 ) ;
assign n44292 =  ( n148 ) ? ( n31660 ) : ( VREG_26_8 ) ;
assign n44293 =  ( n146 ) ? ( n31659 ) : ( n44292 ) ;
assign n44294 =  ( n144 ) ? ( n31658 ) : ( n44293 ) ;
assign n44295 =  ( n142 ) ? ( n31657 ) : ( n44294 ) ;
assign n44296 =  ( n10 ) ? ( n31656 ) : ( n44295 ) ;
assign n44297 =  ( n148 ) ? ( n32694 ) : ( VREG_26_8 ) ;
assign n44298 =  ( n146 ) ? ( n32693 ) : ( n44297 ) ;
assign n44299 =  ( n144 ) ? ( n32692 ) : ( n44298 ) ;
assign n44300 =  ( n142 ) ? ( n32691 ) : ( n44299 ) ;
assign n44301 =  ( n10 ) ? ( n32690 ) : ( n44300 ) ;
assign n44302 =  ( n32701 ) ? ( VREG_26_8 ) : ( n44296 ) ;
assign n44303 =  ( n32701 ) ? ( VREG_26_8 ) : ( n44301 ) ;
assign n44304 =  ( n3034 ) ? ( n44303 ) : ( VREG_26_8 ) ;
assign n44305 =  ( n2965 ) ? ( n44302 ) : ( n44304 ) ;
assign n44306 =  ( n1930 ) ? ( n44301 ) : ( n44305 ) ;
assign n44307 =  ( n879 ) ? ( n44296 ) : ( n44306 ) ;
assign n44308 =  ( n172 ) ? ( n32712 ) : ( VREG_26_8 ) ;
assign n44309 =  ( n170 ) ? ( n32711 ) : ( n44308 ) ;
assign n44310 =  ( n168 ) ? ( n32710 ) : ( n44309 ) ;
assign n44311 =  ( n166 ) ? ( n32709 ) : ( n44310 ) ;
assign n44312 =  ( n162 ) ? ( n32708 ) : ( n44311 ) ;
assign n44313 =  ( n172 ) ? ( n32722 ) : ( VREG_26_8 ) ;
assign n44314 =  ( n170 ) ? ( n32721 ) : ( n44313 ) ;
assign n44315 =  ( n168 ) ? ( n32720 ) : ( n44314 ) ;
assign n44316 =  ( n166 ) ? ( n32719 ) : ( n44315 ) ;
assign n44317 =  ( n162 ) ? ( n32718 ) : ( n44316 ) ;
assign n44318 =  ( n32701 ) ? ( VREG_26_8 ) : ( n44317 ) ;
assign n44319 =  ( n3051 ) ? ( n44318 ) : ( VREG_26_8 ) ;
assign n44320 =  ( n3040 ) ? ( n44312 ) : ( n44319 ) ;
assign n44321 =  ( n192 ) ? ( VREG_26_8 ) : ( VREG_26_8 ) ;
assign n44322 =  ( n157 ) ? ( n44320 ) : ( n44321 ) ;
assign n44323 =  ( n6 ) ? ( n44307 ) : ( n44322 ) ;
assign n44324 =  ( n593 ) ? ( n44323 ) : ( VREG_26_8 ) ;
assign n44325 =  ( n148 ) ? ( n33779 ) : ( VREG_26_9 ) ;
assign n44326 =  ( n146 ) ? ( n33778 ) : ( n44325 ) ;
assign n44327 =  ( n144 ) ? ( n33777 ) : ( n44326 ) ;
assign n44328 =  ( n142 ) ? ( n33776 ) : ( n44327 ) ;
assign n44329 =  ( n10 ) ? ( n33775 ) : ( n44328 ) ;
assign n44330 =  ( n148 ) ? ( n34813 ) : ( VREG_26_9 ) ;
assign n44331 =  ( n146 ) ? ( n34812 ) : ( n44330 ) ;
assign n44332 =  ( n144 ) ? ( n34811 ) : ( n44331 ) ;
assign n44333 =  ( n142 ) ? ( n34810 ) : ( n44332 ) ;
assign n44334 =  ( n10 ) ? ( n34809 ) : ( n44333 ) ;
assign n44335 =  ( n34820 ) ? ( VREG_26_9 ) : ( n44329 ) ;
assign n44336 =  ( n34820 ) ? ( VREG_26_9 ) : ( n44334 ) ;
assign n44337 =  ( n3034 ) ? ( n44336 ) : ( VREG_26_9 ) ;
assign n44338 =  ( n2965 ) ? ( n44335 ) : ( n44337 ) ;
assign n44339 =  ( n1930 ) ? ( n44334 ) : ( n44338 ) ;
assign n44340 =  ( n879 ) ? ( n44329 ) : ( n44339 ) ;
assign n44341 =  ( n172 ) ? ( n34831 ) : ( VREG_26_9 ) ;
assign n44342 =  ( n170 ) ? ( n34830 ) : ( n44341 ) ;
assign n44343 =  ( n168 ) ? ( n34829 ) : ( n44342 ) ;
assign n44344 =  ( n166 ) ? ( n34828 ) : ( n44343 ) ;
assign n44345 =  ( n162 ) ? ( n34827 ) : ( n44344 ) ;
assign n44346 =  ( n172 ) ? ( n34841 ) : ( VREG_26_9 ) ;
assign n44347 =  ( n170 ) ? ( n34840 ) : ( n44346 ) ;
assign n44348 =  ( n168 ) ? ( n34839 ) : ( n44347 ) ;
assign n44349 =  ( n166 ) ? ( n34838 ) : ( n44348 ) ;
assign n44350 =  ( n162 ) ? ( n34837 ) : ( n44349 ) ;
assign n44351 =  ( n34820 ) ? ( VREG_26_9 ) : ( n44350 ) ;
assign n44352 =  ( n3051 ) ? ( n44351 ) : ( VREG_26_9 ) ;
assign n44353 =  ( n3040 ) ? ( n44345 ) : ( n44352 ) ;
assign n44354 =  ( n192 ) ? ( VREG_26_9 ) : ( VREG_26_9 ) ;
assign n44355 =  ( n157 ) ? ( n44353 ) : ( n44354 ) ;
assign n44356 =  ( n6 ) ? ( n44340 ) : ( n44355 ) ;
assign n44357 =  ( n593 ) ? ( n44356 ) : ( VREG_26_9 ) ;
assign n44358 =  ( n148 ) ? ( n1924 ) : ( VREG_27_0 ) ;
assign n44359 =  ( n146 ) ? ( n1923 ) : ( n44358 ) ;
assign n44360 =  ( n144 ) ? ( n1922 ) : ( n44359 ) ;
assign n44361 =  ( n142 ) ? ( n1921 ) : ( n44360 ) ;
assign n44362 =  ( n10 ) ? ( n1920 ) : ( n44361 ) ;
assign n44363 =  ( n148 ) ? ( n2959 ) : ( VREG_27_0 ) ;
assign n44364 =  ( n146 ) ? ( n2958 ) : ( n44363 ) ;
assign n44365 =  ( n144 ) ? ( n2957 ) : ( n44364 ) ;
assign n44366 =  ( n142 ) ? ( n2956 ) : ( n44365 ) ;
assign n44367 =  ( n10 ) ? ( n2955 ) : ( n44366 ) ;
assign n44368 =  ( n3032 ) ? ( VREG_27_0 ) : ( n44362 ) ;
assign n44369 =  ( n3032 ) ? ( VREG_27_0 ) : ( n44367 ) ;
assign n44370 =  ( n3034 ) ? ( n44369 ) : ( VREG_27_0 ) ;
assign n44371 =  ( n2965 ) ? ( n44368 ) : ( n44370 ) ;
assign n44372 =  ( n1930 ) ? ( n44367 ) : ( n44371 ) ;
assign n44373 =  ( n879 ) ? ( n44362 ) : ( n44372 ) ;
assign n44374 =  ( n172 ) ? ( n3045 ) : ( VREG_27_0 ) ;
assign n44375 =  ( n170 ) ? ( n3044 ) : ( n44374 ) ;
assign n44376 =  ( n168 ) ? ( n3043 ) : ( n44375 ) ;
assign n44377 =  ( n166 ) ? ( n3042 ) : ( n44376 ) ;
assign n44378 =  ( n162 ) ? ( n3041 ) : ( n44377 ) ;
assign n44379 =  ( n172 ) ? ( n3056 ) : ( VREG_27_0 ) ;
assign n44380 =  ( n170 ) ? ( n3055 ) : ( n44379 ) ;
assign n44381 =  ( n168 ) ? ( n3054 ) : ( n44380 ) ;
assign n44382 =  ( n166 ) ? ( n3053 ) : ( n44381 ) ;
assign n44383 =  ( n162 ) ? ( n3052 ) : ( n44382 ) ;
assign n44384 =  ( n3032 ) ? ( VREG_27_0 ) : ( n44383 ) ;
assign n44385 =  ( n3051 ) ? ( n44384 ) : ( VREG_27_0 ) ;
assign n44386 =  ( n3040 ) ? ( n44378 ) : ( n44385 ) ;
assign n44387 =  ( n192 ) ? ( VREG_27_0 ) : ( VREG_27_0 ) ;
assign n44388 =  ( n157 ) ? ( n44386 ) : ( n44387 ) ;
assign n44389 =  ( n6 ) ? ( n44373 ) : ( n44388 ) ;
assign n44390 =  ( n615 ) ? ( n44389 ) : ( VREG_27_0 ) ;
assign n44391 =  ( n148 ) ? ( n4113 ) : ( VREG_27_1 ) ;
assign n44392 =  ( n146 ) ? ( n4112 ) : ( n44391 ) ;
assign n44393 =  ( n144 ) ? ( n4111 ) : ( n44392 ) ;
assign n44394 =  ( n142 ) ? ( n4110 ) : ( n44393 ) ;
assign n44395 =  ( n10 ) ? ( n4109 ) : ( n44394 ) ;
assign n44396 =  ( n148 ) ? ( n5147 ) : ( VREG_27_1 ) ;
assign n44397 =  ( n146 ) ? ( n5146 ) : ( n44396 ) ;
assign n44398 =  ( n144 ) ? ( n5145 ) : ( n44397 ) ;
assign n44399 =  ( n142 ) ? ( n5144 ) : ( n44398 ) ;
assign n44400 =  ( n10 ) ? ( n5143 ) : ( n44399 ) ;
assign n44401 =  ( n5154 ) ? ( VREG_27_1 ) : ( n44395 ) ;
assign n44402 =  ( n5154 ) ? ( VREG_27_1 ) : ( n44400 ) ;
assign n44403 =  ( n3034 ) ? ( n44402 ) : ( VREG_27_1 ) ;
assign n44404 =  ( n2965 ) ? ( n44401 ) : ( n44403 ) ;
assign n44405 =  ( n1930 ) ? ( n44400 ) : ( n44404 ) ;
assign n44406 =  ( n879 ) ? ( n44395 ) : ( n44405 ) ;
assign n44407 =  ( n172 ) ? ( n5165 ) : ( VREG_27_1 ) ;
assign n44408 =  ( n170 ) ? ( n5164 ) : ( n44407 ) ;
assign n44409 =  ( n168 ) ? ( n5163 ) : ( n44408 ) ;
assign n44410 =  ( n166 ) ? ( n5162 ) : ( n44409 ) ;
assign n44411 =  ( n162 ) ? ( n5161 ) : ( n44410 ) ;
assign n44412 =  ( n172 ) ? ( n5175 ) : ( VREG_27_1 ) ;
assign n44413 =  ( n170 ) ? ( n5174 ) : ( n44412 ) ;
assign n44414 =  ( n168 ) ? ( n5173 ) : ( n44413 ) ;
assign n44415 =  ( n166 ) ? ( n5172 ) : ( n44414 ) ;
assign n44416 =  ( n162 ) ? ( n5171 ) : ( n44415 ) ;
assign n44417 =  ( n5154 ) ? ( VREG_27_1 ) : ( n44416 ) ;
assign n44418 =  ( n3051 ) ? ( n44417 ) : ( VREG_27_1 ) ;
assign n44419 =  ( n3040 ) ? ( n44411 ) : ( n44418 ) ;
assign n44420 =  ( n192 ) ? ( VREG_27_1 ) : ( VREG_27_1 ) ;
assign n44421 =  ( n157 ) ? ( n44419 ) : ( n44420 ) ;
assign n44422 =  ( n6 ) ? ( n44406 ) : ( n44421 ) ;
assign n44423 =  ( n615 ) ? ( n44422 ) : ( VREG_27_1 ) ;
assign n44424 =  ( n148 ) ? ( n6232 ) : ( VREG_27_10 ) ;
assign n44425 =  ( n146 ) ? ( n6231 ) : ( n44424 ) ;
assign n44426 =  ( n144 ) ? ( n6230 ) : ( n44425 ) ;
assign n44427 =  ( n142 ) ? ( n6229 ) : ( n44426 ) ;
assign n44428 =  ( n10 ) ? ( n6228 ) : ( n44427 ) ;
assign n44429 =  ( n148 ) ? ( n7266 ) : ( VREG_27_10 ) ;
assign n44430 =  ( n146 ) ? ( n7265 ) : ( n44429 ) ;
assign n44431 =  ( n144 ) ? ( n7264 ) : ( n44430 ) ;
assign n44432 =  ( n142 ) ? ( n7263 ) : ( n44431 ) ;
assign n44433 =  ( n10 ) ? ( n7262 ) : ( n44432 ) ;
assign n44434 =  ( n7273 ) ? ( VREG_27_10 ) : ( n44428 ) ;
assign n44435 =  ( n7273 ) ? ( VREG_27_10 ) : ( n44433 ) ;
assign n44436 =  ( n3034 ) ? ( n44435 ) : ( VREG_27_10 ) ;
assign n44437 =  ( n2965 ) ? ( n44434 ) : ( n44436 ) ;
assign n44438 =  ( n1930 ) ? ( n44433 ) : ( n44437 ) ;
assign n44439 =  ( n879 ) ? ( n44428 ) : ( n44438 ) ;
assign n44440 =  ( n172 ) ? ( n7284 ) : ( VREG_27_10 ) ;
assign n44441 =  ( n170 ) ? ( n7283 ) : ( n44440 ) ;
assign n44442 =  ( n168 ) ? ( n7282 ) : ( n44441 ) ;
assign n44443 =  ( n166 ) ? ( n7281 ) : ( n44442 ) ;
assign n44444 =  ( n162 ) ? ( n7280 ) : ( n44443 ) ;
assign n44445 =  ( n172 ) ? ( n7294 ) : ( VREG_27_10 ) ;
assign n44446 =  ( n170 ) ? ( n7293 ) : ( n44445 ) ;
assign n44447 =  ( n168 ) ? ( n7292 ) : ( n44446 ) ;
assign n44448 =  ( n166 ) ? ( n7291 ) : ( n44447 ) ;
assign n44449 =  ( n162 ) ? ( n7290 ) : ( n44448 ) ;
assign n44450 =  ( n7273 ) ? ( VREG_27_10 ) : ( n44449 ) ;
assign n44451 =  ( n3051 ) ? ( n44450 ) : ( VREG_27_10 ) ;
assign n44452 =  ( n3040 ) ? ( n44444 ) : ( n44451 ) ;
assign n44453 =  ( n192 ) ? ( VREG_27_10 ) : ( VREG_27_10 ) ;
assign n44454 =  ( n157 ) ? ( n44452 ) : ( n44453 ) ;
assign n44455 =  ( n6 ) ? ( n44439 ) : ( n44454 ) ;
assign n44456 =  ( n615 ) ? ( n44455 ) : ( VREG_27_10 ) ;
assign n44457 =  ( n148 ) ? ( n8351 ) : ( VREG_27_11 ) ;
assign n44458 =  ( n146 ) ? ( n8350 ) : ( n44457 ) ;
assign n44459 =  ( n144 ) ? ( n8349 ) : ( n44458 ) ;
assign n44460 =  ( n142 ) ? ( n8348 ) : ( n44459 ) ;
assign n44461 =  ( n10 ) ? ( n8347 ) : ( n44460 ) ;
assign n44462 =  ( n148 ) ? ( n9385 ) : ( VREG_27_11 ) ;
assign n44463 =  ( n146 ) ? ( n9384 ) : ( n44462 ) ;
assign n44464 =  ( n144 ) ? ( n9383 ) : ( n44463 ) ;
assign n44465 =  ( n142 ) ? ( n9382 ) : ( n44464 ) ;
assign n44466 =  ( n10 ) ? ( n9381 ) : ( n44465 ) ;
assign n44467 =  ( n9392 ) ? ( VREG_27_11 ) : ( n44461 ) ;
assign n44468 =  ( n9392 ) ? ( VREG_27_11 ) : ( n44466 ) ;
assign n44469 =  ( n3034 ) ? ( n44468 ) : ( VREG_27_11 ) ;
assign n44470 =  ( n2965 ) ? ( n44467 ) : ( n44469 ) ;
assign n44471 =  ( n1930 ) ? ( n44466 ) : ( n44470 ) ;
assign n44472 =  ( n879 ) ? ( n44461 ) : ( n44471 ) ;
assign n44473 =  ( n172 ) ? ( n9403 ) : ( VREG_27_11 ) ;
assign n44474 =  ( n170 ) ? ( n9402 ) : ( n44473 ) ;
assign n44475 =  ( n168 ) ? ( n9401 ) : ( n44474 ) ;
assign n44476 =  ( n166 ) ? ( n9400 ) : ( n44475 ) ;
assign n44477 =  ( n162 ) ? ( n9399 ) : ( n44476 ) ;
assign n44478 =  ( n172 ) ? ( n9413 ) : ( VREG_27_11 ) ;
assign n44479 =  ( n170 ) ? ( n9412 ) : ( n44478 ) ;
assign n44480 =  ( n168 ) ? ( n9411 ) : ( n44479 ) ;
assign n44481 =  ( n166 ) ? ( n9410 ) : ( n44480 ) ;
assign n44482 =  ( n162 ) ? ( n9409 ) : ( n44481 ) ;
assign n44483 =  ( n9392 ) ? ( VREG_27_11 ) : ( n44482 ) ;
assign n44484 =  ( n3051 ) ? ( n44483 ) : ( VREG_27_11 ) ;
assign n44485 =  ( n3040 ) ? ( n44477 ) : ( n44484 ) ;
assign n44486 =  ( n192 ) ? ( VREG_27_11 ) : ( VREG_27_11 ) ;
assign n44487 =  ( n157 ) ? ( n44485 ) : ( n44486 ) ;
assign n44488 =  ( n6 ) ? ( n44472 ) : ( n44487 ) ;
assign n44489 =  ( n615 ) ? ( n44488 ) : ( VREG_27_11 ) ;
assign n44490 =  ( n148 ) ? ( n10470 ) : ( VREG_27_12 ) ;
assign n44491 =  ( n146 ) ? ( n10469 ) : ( n44490 ) ;
assign n44492 =  ( n144 ) ? ( n10468 ) : ( n44491 ) ;
assign n44493 =  ( n142 ) ? ( n10467 ) : ( n44492 ) ;
assign n44494 =  ( n10 ) ? ( n10466 ) : ( n44493 ) ;
assign n44495 =  ( n148 ) ? ( n11504 ) : ( VREG_27_12 ) ;
assign n44496 =  ( n146 ) ? ( n11503 ) : ( n44495 ) ;
assign n44497 =  ( n144 ) ? ( n11502 ) : ( n44496 ) ;
assign n44498 =  ( n142 ) ? ( n11501 ) : ( n44497 ) ;
assign n44499 =  ( n10 ) ? ( n11500 ) : ( n44498 ) ;
assign n44500 =  ( n11511 ) ? ( VREG_27_12 ) : ( n44494 ) ;
assign n44501 =  ( n11511 ) ? ( VREG_27_12 ) : ( n44499 ) ;
assign n44502 =  ( n3034 ) ? ( n44501 ) : ( VREG_27_12 ) ;
assign n44503 =  ( n2965 ) ? ( n44500 ) : ( n44502 ) ;
assign n44504 =  ( n1930 ) ? ( n44499 ) : ( n44503 ) ;
assign n44505 =  ( n879 ) ? ( n44494 ) : ( n44504 ) ;
assign n44506 =  ( n172 ) ? ( n11522 ) : ( VREG_27_12 ) ;
assign n44507 =  ( n170 ) ? ( n11521 ) : ( n44506 ) ;
assign n44508 =  ( n168 ) ? ( n11520 ) : ( n44507 ) ;
assign n44509 =  ( n166 ) ? ( n11519 ) : ( n44508 ) ;
assign n44510 =  ( n162 ) ? ( n11518 ) : ( n44509 ) ;
assign n44511 =  ( n172 ) ? ( n11532 ) : ( VREG_27_12 ) ;
assign n44512 =  ( n170 ) ? ( n11531 ) : ( n44511 ) ;
assign n44513 =  ( n168 ) ? ( n11530 ) : ( n44512 ) ;
assign n44514 =  ( n166 ) ? ( n11529 ) : ( n44513 ) ;
assign n44515 =  ( n162 ) ? ( n11528 ) : ( n44514 ) ;
assign n44516 =  ( n11511 ) ? ( VREG_27_12 ) : ( n44515 ) ;
assign n44517 =  ( n3051 ) ? ( n44516 ) : ( VREG_27_12 ) ;
assign n44518 =  ( n3040 ) ? ( n44510 ) : ( n44517 ) ;
assign n44519 =  ( n192 ) ? ( VREG_27_12 ) : ( VREG_27_12 ) ;
assign n44520 =  ( n157 ) ? ( n44518 ) : ( n44519 ) ;
assign n44521 =  ( n6 ) ? ( n44505 ) : ( n44520 ) ;
assign n44522 =  ( n615 ) ? ( n44521 ) : ( VREG_27_12 ) ;
assign n44523 =  ( n148 ) ? ( n12589 ) : ( VREG_27_13 ) ;
assign n44524 =  ( n146 ) ? ( n12588 ) : ( n44523 ) ;
assign n44525 =  ( n144 ) ? ( n12587 ) : ( n44524 ) ;
assign n44526 =  ( n142 ) ? ( n12586 ) : ( n44525 ) ;
assign n44527 =  ( n10 ) ? ( n12585 ) : ( n44526 ) ;
assign n44528 =  ( n148 ) ? ( n13623 ) : ( VREG_27_13 ) ;
assign n44529 =  ( n146 ) ? ( n13622 ) : ( n44528 ) ;
assign n44530 =  ( n144 ) ? ( n13621 ) : ( n44529 ) ;
assign n44531 =  ( n142 ) ? ( n13620 ) : ( n44530 ) ;
assign n44532 =  ( n10 ) ? ( n13619 ) : ( n44531 ) ;
assign n44533 =  ( n13630 ) ? ( VREG_27_13 ) : ( n44527 ) ;
assign n44534 =  ( n13630 ) ? ( VREG_27_13 ) : ( n44532 ) ;
assign n44535 =  ( n3034 ) ? ( n44534 ) : ( VREG_27_13 ) ;
assign n44536 =  ( n2965 ) ? ( n44533 ) : ( n44535 ) ;
assign n44537 =  ( n1930 ) ? ( n44532 ) : ( n44536 ) ;
assign n44538 =  ( n879 ) ? ( n44527 ) : ( n44537 ) ;
assign n44539 =  ( n172 ) ? ( n13641 ) : ( VREG_27_13 ) ;
assign n44540 =  ( n170 ) ? ( n13640 ) : ( n44539 ) ;
assign n44541 =  ( n168 ) ? ( n13639 ) : ( n44540 ) ;
assign n44542 =  ( n166 ) ? ( n13638 ) : ( n44541 ) ;
assign n44543 =  ( n162 ) ? ( n13637 ) : ( n44542 ) ;
assign n44544 =  ( n172 ) ? ( n13651 ) : ( VREG_27_13 ) ;
assign n44545 =  ( n170 ) ? ( n13650 ) : ( n44544 ) ;
assign n44546 =  ( n168 ) ? ( n13649 ) : ( n44545 ) ;
assign n44547 =  ( n166 ) ? ( n13648 ) : ( n44546 ) ;
assign n44548 =  ( n162 ) ? ( n13647 ) : ( n44547 ) ;
assign n44549 =  ( n13630 ) ? ( VREG_27_13 ) : ( n44548 ) ;
assign n44550 =  ( n3051 ) ? ( n44549 ) : ( VREG_27_13 ) ;
assign n44551 =  ( n3040 ) ? ( n44543 ) : ( n44550 ) ;
assign n44552 =  ( n192 ) ? ( VREG_27_13 ) : ( VREG_27_13 ) ;
assign n44553 =  ( n157 ) ? ( n44551 ) : ( n44552 ) ;
assign n44554 =  ( n6 ) ? ( n44538 ) : ( n44553 ) ;
assign n44555 =  ( n615 ) ? ( n44554 ) : ( VREG_27_13 ) ;
assign n44556 =  ( n148 ) ? ( n14708 ) : ( VREG_27_14 ) ;
assign n44557 =  ( n146 ) ? ( n14707 ) : ( n44556 ) ;
assign n44558 =  ( n144 ) ? ( n14706 ) : ( n44557 ) ;
assign n44559 =  ( n142 ) ? ( n14705 ) : ( n44558 ) ;
assign n44560 =  ( n10 ) ? ( n14704 ) : ( n44559 ) ;
assign n44561 =  ( n148 ) ? ( n15742 ) : ( VREG_27_14 ) ;
assign n44562 =  ( n146 ) ? ( n15741 ) : ( n44561 ) ;
assign n44563 =  ( n144 ) ? ( n15740 ) : ( n44562 ) ;
assign n44564 =  ( n142 ) ? ( n15739 ) : ( n44563 ) ;
assign n44565 =  ( n10 ) ? ( n15738 ) : ( n44564 ) ;
assign n44566 =  ( n15749 ) ? ( VREG_27_14 ) : ( n44560 ) ;
assign n44567 =  ( n15749 ) ? ( VREG_27_14 ) : ( n44565 ) ;
assign n44568 =  ( n3034 ) ? ( n44567 ) : ( VREG_27_14 ) ;
assign n44569 =  ( n2965 ) ? ( n44566 ) : ( n44568 ) ;
assign n44570 =  ( n1930 ) ? ( n44565 ) : ( n44569 ) ;
assign n44571 =  ( n879 ) ? ( n44560 ) : ( n44570 ) ;
assign n44572 =  ( n172 ) ? ( n15760 ) : ( VREG_27_14 ) ;
assign n44573 =  ( n170 ) ? ( n15759 ) : ( n44572 ) ;
assign n44574 =  ( n168 ) ? ( n15758 ) : ( n44573 ) ;
assign n44575 =  ( n166 ) ? ( n15757 ) : ( n44574 ) ;
assign n44576 =  ( n162 ) ? ( n15756 ) : ( n44575 ) ;
assign n44577 =  ( n172 ) ? ( n15770 ) : ( VREG_27_14 ) ;
assign n44578 =  ( n170 ) ? ( n15769 ) : ( n44577 ) ;
assign n44579 =  ( n168 ) ? ( n15768 ) : ( n44578 ) ;
assign n44580 =  ( n166 ) ? ( n15767 ) : ( n44579 ) ;
assign n44581 =  ( n162 ) ? ( n15766 ) : ( n44580 ) ;
assign n44582 =  ( n15749 ) ? ( VREG_27_14 ) : ( n44581 ) ;
assign n44583 =  ( n3051 ) ? ( n44582 ) : ( VREG_27_14 ) ;
assign n44584 =  ( n3040 ) ? ( n44576 ) : ( n44583 ) ;
assign n44585 =  ( n192 ) ? ( VREG_27_14 ) : ( VREG_27_14 ) ;
assign n44586 =  ( n157 ) ? ( n44584 ) : ( n44585 ) ;
assign n44587 =  ( n6 ) ? ( n44571 ) : ( n44586 ) ;
assign n44588 =  ( n615 ) ? ( n44587 ) : ( VREG_27_14 ) ;
assign n44589 =  ( n148 ) ? ( n16827 ) : ( VREG_27_15 ) ;
assign n44590 =  ( n146 ) ? ( n16826 ) : ( n44589 ) ;
assign n44591 =  ( n144 ) ? ( n16825 ) : ( n44590 ) ;
assign n44592 =  ( n142 ) ? ( n16824 ) : ( n44591 ) ;
assign n44593 =  ( n10 ) ? ( n16823 ) : ( n44592 ) ;
assign n44594 =  ( n148 ) ? ( n17861 ) : ( VREG_27_15 ) ;
assign n44595 =  ( n146 ) ? ( n17860 ) : ( n44594 ) ;
assign n44596 =  ( n144 ) ? ( n17859 ) : ( n44595 ) ;
assign n44597 =  ( n142 ) ? ( n17858 ) : ( n44596 ) ;
assign n44598 =  ( n10 ) ? ( n17857 ) : ( n44597 ) ;
assign n44599 =  ( n17868 ) ? ( VREG_27_15 ) : ( n44593 ) ;
assign n44600 =  ( n17868 ) ? ( VREG_27_15 ) : ( n44598 ) ;
assign n44601 =  ( n3034 ) ? ( n44600 ) : ( VREG_27_15 ) ;
assign n44602 =  ( n2965 ) ? ( n44599 ) : ( n44601 ) ;
assign n44603 =  ( n1930 ) ? ( n44598 ) : ( n44602 ) ;
assign n44604 =  ( n879 ) ? ( n44593 ) : ( n44603 ) ;
assign n44605 =  ( n172 ) ? ( n17879 ) : ( VREG_27_15 ) ;
assign n44606 =  ( n170 ) ? ( n17878 ) : ( n44605 ) ;
assign n44607 =  ( n168 ) ? ( n17877 ) : ( n44606 ) ;
assign n44608 =  ( n166 ) ? ( n17876 ) : ( n44607 ) ;
assign n44609 =  ( n162 ) ? ( n17875 ) : ( n44608 ) ;
assign n44610 =  ( n172 ) ? ( n17889 ) : ( VREG_27_15 ) ;
assign n44611 =  ( n170 ) ? ( n17888 ) : ( n44610 ) ;
assign n44612 =  ( n168 ) ? ( n17887 ) : ( n44611 ) ;
assign n44613 =  ( n166 ) ? ( n17886 ) : ( n44612 ) ;
assign n44614 =  ( n162 ) ? ( n17885 ) : ( n44613 ) ;
assign n44615 =  ( n17868 ) ? ( VREG_27_15 ) : ( n44614 ) ;
assign n44616 =  ( n3051 ) ? ( n44615 ) : ( VREG_27_15 ) ;
assign n44617 =  ( n3040 ) ? ( n44609 ) : ( n44616 ) ;
assign n44618 =  ( n192 ) ? ( VREG_27_15 ) : ( VREG_27_15 ) ;
assign n44619 =  ( n157 ) ? ( n44617 ) : ( n44618 ) ;
assign n44620 =  ( n6 ) ? ( n44604 ) : ( n44619 ) ;
assign n44621 =  ( n615 ) ? ( n44620 ) : ( VREG_27_15 ) ;
assign n44622 =  ( n148 ) ? ( n18946 ) : ( VREG_27_2 ) ;
assign n44623 =  ( n146 ) ? ( n18945 ) : ( n44622 ) ;
assign n44624 =  ( n144 ) ? ( n18944 ) : ( n44623 ) ;
assign n44625 =  ( n142 ) ? ( n18943 ) : ( n44624 ) ;
assign n44626 =  ( n10 ) ? ( n18942 ) : ( n44625 ) ;
assign n44627 =  ( n148 ) ? ( n19980 ) : ( VREG_27_2 ) ;
assign n44628 =  ( n146 ) ? ( n19979 ) : ( n44627 ) ;
assign n44629 =  ( n144 ) ? ( n19978 ) : ( n44628 ) ;
assign n44630 =  ( n142 ) ? ( n19977 ) : ( n44629 ) ;
assign n44631 =  ( n10 ) ? ( n19976 ) : ( n44630 ) ;
assign n44632 =  ( n19987 ) ? ( VREG_27_2 ) : ( n44626 ) ;
assign n44633 =  ( n19987 ) ? ( VREG_27_2 ) : ( n44631 ) ;
assign n44634 =  ( n3034 ) ? ( n44633 ) : ( VREG_27_2 ) ;
assign n44635 =  ( n2965 ) ? ( n44632 ) : ( n44634 ) ;
assign n44636 =  ( n1930 ) ? ( n44631 ) : ( n44635 ) ;
assign n44637 =  ( n879 ) ? ( n44626 ) : ( n44636 ) ;
assign n44638 =  ( n172 ) ? ( n19998 ) : ( VREG_27_2 ) ;
assign n44639 =  ( n170 ) ? ( n19997 ) : ( n44638 ) ;
assign n44640 =  ( n168 ) ? ( n19996 ) : ( n44639 ) ;
assign n44641 =  ( n166 ) ? ( n19995 ) : ( n44640 ) ;
assign n44642 =  ( n162 ) ? ( n19994 ) : ( n44641 ) ;
assign n44643 =  ( n172 ) ? ( n20008 ) : ( VREG_27_2 ) ;
assign n44644 =  ( n170 ) ? ( n20007 ) : ( n44643 ) ;
assign n44645 =  ( n168 ) ? ( n20006 ) : ( n44644 ) ;
assign n44646 =  ( n166 ) ? ( n20005 ) : ( n44645 ) ;
assign n44647 =  ( n162 ) ? ( n20004 ) : ( n44646 ) ;
assign n44648 =  ( n19987 ) ? ( VREG_27_2 ) : ( n44647 ) ;
assign n44649 =  ( n3051 ) ? ( n44648 ) : ( VREG_27_2 ) ;
assign n44650 =  ( n3040 ) ? ( n44642 ) : ( n44649 ) ;
assign n44651 =  ( n192 ) ? ( VREG_27_2 ) : ( VREG_27_2 ) ;
assign n44652 =  ( n157 ) ? ( n44650 ) : ( n44651 ) ;
assign n44653 =  ( n6 ) ? ( n44637 ) : ( n44652 ) ;
assign n44654 =  ( n615 ) ? ( n44653 ) : ( VREG_27_2 ) ;
assign n44655 =  ( n148 ) ? ( n21065 ) : ( VREG_27_3 ) ;
assign n44656 =  ( n146 ) ? ( n21064 ) : ( n44655 ) ;
assign n44657 =  ( n144 ) ? ( n21063 ) : ( n44656 ) ;
assign n44658 =  ( n142 ) ? ( n21062 ) : ( n44657 ) ;
assign n44659 =  ( n10 ) ? ( n21061 ) : ( n44658 ) ;
assign n44660 =  ( n148 ) ? ( n22099 ) : ( VREG_27_3 ) ;
assign n44661 =  ( n146 ) ? ( n22098 ) : ( n44660 ) ;
assign n44662 =  ( n144 ) ? ( n22097 ) : ( n44661 ) ;
assign n44663 =  ( n142 ) ? ( n22096 ) : ( n44662 ) ;
assign n44664 =  ( n10 ) ? ( n22095 ) : ( n44663 ) ;
assign n44665 =  ( n22106 ) ? ( VREG_27_3 ) : ( n44659 ) ;
assign n44666 =  ( n22106 ) ? ( VREG_27_3 ) : ( n44664 ) ;
assign n44667 =  ( n3034 ) ? ( n44666 ) : ( VREG_27_3 ) ;
assign n44668 =  ( n2965 ) ? ( n44665 ) : ( n44667 ) ;
assign n44669 =  ( n1930 ) ? ( n44664 ) : ( n44668 ) ;
assign n44670 =  ( n879 ) ? ( n44659 ) : ( n44669 ) ;
assign n44671 =  ( n172 ) ? ( n22117 ) : ( VREG_27_3 ) ;
assign n44672 =  ( n170 ) ? ( n22116 ) : ( n44671 ) ;
assign n44673 =  ( n168 ) ? ( n22115 ) : ( n44672 ) ;
assign n44674 =  ( n166 ) ? ( n22114 ) : ( n44673 ) ;
assign n44675 =  ( n162 ) ? ( n22113 ) : ( n44674 ) ;
assign n44676 =  ( n172 ) ? ( n22127 ) : ( VREG_27_3 ) ;
assign n44677 =  ( n170 ) ? ( n22126 ) : ( n44676 ) ;
assign n44678 =  ( n168 ) ? ( n22125 ) : ( n44677 ) ;
assign n44679 =  ( n166 ) ? ( n22124 ) : ( n44678 ) ;
assign n44680 =  ( n162 ) ? ( n22123 ) : ( n44679 ) ;
assign n44681 =  ( n22106 ) ? ( VREG_27_3 ) : ( n44680 ) ;
assign n44682 =  ( n3051 ) ? ( n44681 ) : ( VREG_27_3 ) ;
assign n44683 =  ( n3040 ) ? ( n44675 ) : ( n44682 ) ;
assign n44684 =  ( n192 ) ? ( VREG_27_3 ) : ( VREG_27_3 ) ;
assign n44685 =  ( n157 ) ? ( n44683 ) : ( n44684 ) ;
assign n44686 =  ( n6 ) ? ( n44670 ) : ( n44685 ) ;
assign n44687 =  ( n615 ) ? ( n44686 ) : ( VREG_27_3 ) ;
assign n44688 =  ( n148 ) ? ( n23184 ) : ( VREG_27_4 ) ;
assign n44689 =  ( n146 ) ? ( n23183 ) : ( n44688 ) ;
assign n44690 =  ( n144 ) ? ( n23182 ) : ( n44689 ) ;
assign n44691 =  ( n142 ) ? ( n23181 ) : ( n44690 ) ;
assign n44692 =  ( n10 ) ? ( n23180 ) : ( n44691 ) ;
assign n44693 =  ( n148 ) ? ( n24218 ) : ( VREG_27_4 ) ;
assign n44694 =  ( n146 ) ? ( n24217 ) : ( n44693 ) ;
assign n44695 =  ( n144 ) ? ( n24216 ) : ( n44694 ) ;
assign n44696 =  ( n142 ) ? ( n24215 ) : ( n44695 ) ;
assign n44697 =  ( n10 ) ? ( n24214 ) : ( n44696 ) ;
assign n44698 =  ( n24225 ) ? ( VREG_27_4 ) : ( n44692 ) ;
assign n44699 =  ( n24225 ) ? ( VREG_27_4 ) : ( n44697 ) ;
assign n44700 =  ( n3034 ) ? ( n44699 ) : ( VREG_27_4 ) ;
assign n44701 =  ( n2965 ) ? ( n44698 ) : ( n44700 ) ;
assign n44702 =  ( n1930 ) ? ( n44697 ) : ( n44701 ) ;
assign n44703 =  ( n879 ) ? ( n44692 ) : ( n44702 ) ;
assign n44704 =  ( n172 ) ? ( n24236 ) : ( VREG_27_4 ) ;
assign n44705 =  ( n170 ) ? ( n24235 ) : ( n44704 ) ;
assign n44706 =  ( n168 ) ? ( n24234 ) : ( n44705 ) ;
assign n44707 =  ( n166 ) ? ( n24233 ) : ( n44706 ) ;
assign n44708 =  ( n162 ) ? ( n24232 ) : ( n44707 ) ;
assign n44709 =  ( n172 ) ? ( n24246 ) : ( VREG_27_4 ) ;
assign n44710 =  ( n170 ) ? ( n24245 ) : ( n44709 ) ;
assign n44711 =  ( n168 ) ? ( n24244 ) : ( n44710 ) ;
assign n44712 =  ( n166 ) ? ( n24243 ) : ( n44711 ) ;
assign n44713 =  ( n162 ) ? ( n24242 ) : ( n44712 ) ;
assign n44714 =  ( n24225 ) ? ( VREG_27_4 ) : ( n44713 ) ;
assign n44715 =  ( n3051 ) ? ( n44714 ) : ( VREG_27_4 ) ;
assign n44716 =  ( n3040 ) ? ( n44708 ) : ( n44715 ) ;
assign n44717 =  ( n192 ) ? ( VREG_27_4 ) : ( VREG_27_4 ) ;
assign n44718 =  ( n157 ) ? ( n44716 ) : ( n44717 ) ;
assign n44719 =  ( n6 ) ? ( n44703 ) : ( n44718 ) ;
assign n44720 =  ( n615 ) ? ( n44719 ) : ( VREG_27_4 ) ;
assign n44721 =  ( n148 ) ? ( n25303 ) : ( VREG_27_5 ) ;
assign n44722 =  ( n146 ) ? ( n25302 ) : ( n44721 ) ;
assign n44723 =  ( n144 ) ? ( n25301 ) : ( n44722 ) ;
assign n44724 =  ( n142 ) ? ( n25300 ) : ( n44723 ) ;
assign n44725 =  ( n10 ) ? ( n25299 ) : ( n44724 ) ;
assign n44726 =  ( n148 ) ? ( n26337 ) : ( VREG_27_5 ) ;
assign n44727 =  ( n146 ) ? ( n26336 ) : ( n44726 ) ;
assign n44728 =  ( n144 ) ? ( n26335 ) : ( n44727 ) ;
assign n44729 =  ( n142 ) ? ( n26334 ) : ( n44728 ) ;
assign n44730 =  ( n10 ) ? ( n26333 ) : ( n44729 ) ;
assign n44731 =  ( n26344 ) ? ( VREG_27_5 ) : ( n44725 ) ;
assign n44732 =  ( n26344 ) ? ( VREG_27_5 ) : ( n44730 ) ;
assign n44733 =  ( n3034 ) ? ( n44732 ) : ( VREG_27_5 ) ;
assign n44734 =  ( n2965 ) ? ( n44731 ) : ( n44733 ) ;
assign n44735 =  ( n1930 ) ? ( n44730 ) : ( n44734 ) ;
assign n44736 =  ( n879 ) ? ( n44725 ) : ( n44735 ) ;
assign n44737 =  ( n172 ) ? ( n26355 ) : ( VREG_27_5 ) ;
assign n44738 =  ( n170 ) ? ( n26354 ) : ( n44737 ) ;
assign n44739 =  ( n168 ) ? ( n26353 ) : ( n44738 ) ;
assign n44740 =  ( n166 ) ? ( n26352 ) : ( n44739 ) ;
assign n44741 =  ( n162 ) ? ( n26351 ) : ( n44740 ) ;
assign n44742 =  ( n172 ) ? ( n26365 ) : ( VREG_27_5 ) ;
assign n44743 =  ( n170 ) ? ( n26364 ) : ( n44742 ) ;
assign n44744 =  ( n168 ) ? ( n26363 ) : ( n44743 ) ;
assign n44745 =  ( n166 ) ? ( n26362 ) : ( n44744 ) ;
assign n44746 =  ( n162 ) ? ( n26361 ) : ( n44745 ) ;
assign n44747 =  ( n26344 ) ? ( VREG_27_5 ) : ( n44746 ) ;
assign n44748 =  ( n3051 ) ? ( n44747 ) : ( VREG_27_5 ) ;
assign n44749 =  ( n3040 ) ? ( n44741 ) : ( n44748 ) ;
assign n44750 =  ( n192 ) ? ( VREG_27_5 ) : ( VREG_27_5 ) ;
assign n44751 =  ( n157 ) ? ( n44749 ) : ( n44750 ) ;
assign n44752 =  ( n6 ) ? ( n44736 ) : ( n44751 ) ;
assign n44753 =  ( n615 ) ? ( n44752 ) : ( VREG_27_5 ) ;
assign n44754 =  ( n148 ) ? ( n27422 ) : ( VREG_27_6 ) ;
assign n44755 =  ( n146 ) ? ( n27421 ) : ( n44754 ) ;
assign n44756 =  ( n144 ) ? ( n27420 ) : ( n44755 ) ;
assign n44757 =  ( n142 ) ? ( n27419 ) : ( n44756 ) ;
assign n44758 =  ( n10 ) ? ( n27418 ) : ( n44757 ) ;
assign n44759 =  ( n148 ) ? ( n28456 ) : ( VREG_27_6 ) ;
assign n44760 =  ( n146 ) ? ( n28455 ) : ( n44759 ) ;
assign n44761 =  ( n144 ) ? ( n28454 ) : ( n44760 ) ;
assign n44762 =  ( n142 ) ? ( n28453 ) : ( n44761 ) ;
assign n44763 =  ( n10 ) ? ( n28452 ) : ( n44762 ) ;
assign n44764 =  ( n28463 ) ? ( VREG_27_6 ) : ( n44758 ) ;
assign n44765 =  ( n28463 ) ? ( VREG_27_6 ) : ( n44763 ) ;
assign n44766 =  ( n3034 ) ? ( n44765 ) : ( VREG_27_6 ) ;
assign n44767 =  ( n2965 ) ? ( n44764 ) : ( n44766 ) ;
assign n44768 =  ( n1930 ) ? ( n44763 ) : ( n44767 ) ;
assign n44769 =  ( n879 ) ? ( n44758 ) : ( n44768 ) ;
assign n44770 =  ( n172 ) ? ( n28474 ) : ( VREG_27_6 ) ;
assign n44771 =  ( n170 ) ? ( n28473 ) : ( n44770 ) ;
assign n44772 =  ( n168 ) ? ( n28472 ) : ( n44771 ) ;
assign n44773 =  ( n166 ) ? ( n28471 ) : ( n44772 ) ;
assign n44774 =  ( n162 ) ? ( n28470 ) : ( n44773 ) ;
assign n44775 =  ( n172 ) ? ( n28484 ) : ( VREG_27_6 ) ;
assign n44776 =  ( n170 ) ? ( n28483 ) : ( n44775 ) ;
assign n44777 =  ( n168 ) ? ( n28482 ) : ( n44776 ) ;
assign n44778 =  ( n166 ) ? ( n28481 ) : ( n44777 ) ;
assign n44779 =  ( n162 ) ? ( n28480 ) : ( n44778 ) ;
assign n44780 =  ( n28463 ) ? ( VREG_27_6 ) : ( n44779 ) ;
assign n44781 =  ( n3051 ) ? ( n44780 ) : ( VREG_27_6 ) ;
assign n44782 =  ( n3040 ) ? ( n44774 ) : ( n44781 ) ;
assign n44783 =  ( n192 ) ? ( VREG_27_6 ) : ( VREG_27_6 ) ;
assign n44784 =  ( n157 ) ? ( n44782 ) : ( n44783 ) ;
assign n44785 =  ( n6 ) ? ( n44769 ) : ( n44784 ) ;
assign n44786 =  ( n615 ) ? ( n44785 ) : ( VREG_27_6 ) ;
assign n44787 =  ( n148 ) ? ( n29541 ) : ( VREG_27_7 ) ;
assign n44788 =  ( n146 ) ? ( n29540 ) : ( n44787 ) ;
assign n44789 =  ( n144 ) ? ( n29539 ) : ( n44788 ) ;
assign n44790 =  ( n142 ) ? ( n29538 ) : ( n44789 ) ;
assign n44791 =  ( n10 ) ? ( n29537 ) : ( n44790 ) ;
assign n44792 =  ( n148 ) ? ( n30575 ) : ( VREG_27_7 ) ;
assign n44793 =  ( n146 ) ? ( n30574 ) : ( n44792 ) ;
assign n44794 =  ( n144 ) ? ( n30573 ) : ( n44793 ) ;
assign n44795 =  ( n142 ) ? ( n30572 ) : ( n44794 ) ;
assign n44796 =  ( n10 ) ? ( n30571 ) : ( n44795 ) ;
assign n44797 =  ( n30582 ) ? ( VREG_27_7 ) : ( n44791 ) ;
assign n44798 =  ( n30582 ) ? ( VREG_27_7 ) : ( n44796 ) ;
assign n44799 =  ( n3034 ) ? ( n44798 ) : ( VREG_27_7 ) ;
assign n44800 =  ( n2965 ) ? ( n44797 ) : ( n44799 ) ;
assign n44801 =  ( n1930 ) ? ( n44796 ) : ( n44800 ) ;
assign n44802 =  ( n879 ) ? ( n44791 ) : ( n44801 ) ;
assign n44803 =  ( n172 ) ? ( n30593 ) : ( VREG_27_7 ) ;
assign n44804 =  ( n170 ) ? ( n30592 ) : ( n44803 ) ;
assign n44805 =  ( n168 ) ? ( n30591 ) : ( n44804 ) ;
assign n44806 =  ( n166 ) ? ( n30590 ) : ( n44805 ) ;
assign n44807 =  ( n162 ) ? ( n30589 ) : ( n44806 ) ;
assign n44808 =  ( n172 ) ? ( n30603 ) : ( VREG_27_7 ) ;
assign n44809 =  ( n170 ) ? ( n30602 ) : ( n44808 ) ;
assign n44810 =  ( n168 ) ? ( n30601 ) : ( n44809 ) ;
assign n44811 =  ( n166 ) ? ( n30600 ) : ( n44810 ) ;
assign n44812 =  ( n162 ) ? ( n30599 ) : ( n44811 ) ;
assign n44813 =  ( n30582 ) ? ( VREG_27_7 ) : ( n44812 ) ;
assign n44814 =  ( n3051 ) ? ( n44813 ) : ( VREG_27_7 ) ;
assign n44815 =  ( n3040 ) ? ( n44807 ) : ( n44814 ) ;
assign n44816 =  ( n192 ) ? ( VREG_27_7 ) : ( VREG_27_7 ) ;
assign n44817 =  ( n157 ) ? ( n44815 ) : ( n44816 ) ;
assign n44818 =  ( n6 ) ? ( n44802 ) : ( n44817 ) ;
assign n44819 =  ( n615 ) ? ( n44818 ) : ( VREG_27_7 ) ;
assign n44820 =  ( n148 ) ? ( n31660 ) : ( VREG_27_8 ) ;
assign n44821 =  ( n146 ) ? ( n31659 ) : ( n44820 ) ;
assign n44822 =  ( n144 ) ? ( n31658 ) : ( n44821 ) ;
assign n44823 =  ( n142 ) ? ( n31657 ) : ( n44822 ) ;
assign n44824 =  ( n10 ) ? ( n31656 ) : ( n44823 ) ;
assign n44825 =  ( n148 ) ? ( n32694 ) : ( VREG_27_8 ) ;
assign n44826 =  ( n146 ) ? ( n32693 ) : ( n44825 ) ;
assign n44827 =  ( n144 ) ? ( n32692 ) : ( n44826 ) ;
assign n44828 =  ( n142 ) ? ( n32691 ) : ( n44827 ) ;
assign n44829 =  ( n10 ) ? ( n32690 ) : ( n44828 ) ;
assign n44830 =  ( n32701 ) ? ( VREG_27_8 ) : ( n44824 ) ;
assign n44831 =  ( n32701 ) ? ( VREG_27_8 ) : ( n44829 ) ;
assign n44832 =  ( n3034 ) ? ( n44831 ) : ( VREG_27_8 ) ;
assign n44833 =  ( n2965 ) ? ( n44830 ) : ( n44832 ) ;
assign n44834 =  ( n1930 ) ? ( n44829 ) : ( n44833 ) ;
assign n44835 =  ( n879 ) ? ( n44824 ) : ( n44834 ) ;
assign n44836 =  ( n172 ) ? ( n32712 ) : ( VREG_27_8 ) ;
assign n44837 =  ( n170 ) ? ( n32711 ) : ( n44836 ) ;
assign n44838 =  ( n168 ) ? ( n32710 ) : ( n44837 ) ;
assign n44839 =  ( n166 ) ? ( n32709 ) : ( n44838 ) ;
assign n44840 =  ( n162 ) ? ( n32708 ) : ( n44839 ) ;
assign n44841 =  ( n172 ) ? ( n32722 ) : ( VREG_27_8 ) ;
assign n44842 =  ( n170 ) ? ( n32721 ) : ( n44841 ) ;
assign n44843 =  ( n168 ) ? ( n32720 ) : ( n44842 ) ;
assign n44844 =  ( n166 ) ? ( n32719 ) : ( n44843 ) ;
assign n44845 =  ( n162 ) ? ( n32718 ) : ( n44844 ) ;
assign n44846 =  ( n32701 ) ? ( VREG_27_8 ) : ( n44845 ) ;
assign n44847 =  ( n3051 ) ? ( n44846 ) : ( VREG_27_8 ) ;
assign n44848 =  ( n3040 ) ? ( n44840 ) : ( n44847 ) ;
assign n44849 =  ( n192 ) ? ( VREG_27_8 ) : ( VREG_27_8 ) ;
assign n44850 =  ( n157 ) ? ( n44848 ) : ( n44849 ) ;
assign n44851 =  ( n6 ) ? ( n44835 ) : ( n44850 ) ;
assign n44852 =  ( n615 ) ? ( n44851 ) : ( VREG_27_8 ) ;
assign n44853 =  ( n148 ) ? ( n33779 ) : ( VREG_27_9 ) ;
assign n44854 =  ( n146 ) ? ( n33778 ) : ( n44853 ) ;
assign n44855 =  ( n144 ) ? ( n33777 ) : ( n44854 ) ;
assign n44856 =  ( n142 ) ? ( n33776 ) : ( n44855 ) ;
assign n44857 =  ( n10 ) ? ( n33775 ) : ( n44856 ) ;
assign n44858 =  ( n148 ) ? ( n34813 ) : ( VREG_27_9 ) ;
assign n44859 =  ( n146 ) ? ( n34812 ) : ( n44858 ) ;
assign n44860 =  ( n144 ) ? ( n34811 ) : ( n44859 ) ;
assign n44861 =  ( n142 ) ? ( n34810 ) : ( n44860 ) ;
assign n44862 =  ( n10 ) ? ( n34809 ) : ( n44861 ) ;
assign n44863 =  ( n34820 ) ? ( VREG_27_9 ) : ( n44857 ) ;
assign n44864 =  ( n34820 ) ? ( VREG_27_9 ) : ( n44862 ) ;
assign n44865 =  ( n3034 ) ? ( n44864 ) : ( VREG_27_9 ) ;
assign n44866 =  ( n2965 ) ? ( n44863 ) : ( n44865 ) ;
assign n44867 =  ( n1930 ) ? ( n44862 ) : ( n44866 ) ;
assign n44868 =  ( n879 ) ? ( n44857 ) : ( n44867 ) ;
assign n44869 =  ( n172 ) ? ( n34831 ) : ( VREG_27_9 ) ;
assign n44870 =  ( n170 ) ? ( n34830 ) : ( n44869 ) ;
assign n44871 =  ( n168 ) ? ( n34829 ) : ( n44870 ) ;
assign n44872 =  ( n166 ) ? ( n34828 ) : ( n44871 ) ;
assign n44873 =  ( n162 ) ? ( n34827 ) : ( n44872 ) ;
assign n44874 =  ( n172 ) ? ( n34841 ) : ( VREG_27_9 ) ;
assign n44875 =  ( n170 ) ? ( n34840 ) : ( n44874 ) ;
assign n44876 =  ( n168 ) ? ( n34839 ) : ( n44875 ) ;
assign n44877 =  ( n166 ) ? ( n34838 ) : ( n44876 ) ;
assign n44878 =  ( n162 ) ? ( n34837 ) : ( n44877 ) ;
assign n44879 =  ( n34820 ) ? ( VREG_27_9 ) : ( n44878 ) ;
assign n44880 =  ( n3051 ) ? ( n44879 ) : ( VREG_27_9 ) ;
assign n44881 =  ( n3040 ) ? ( n44873 ) : ( n44880 ) ;
assign n44882 =  ( n192 ) ? ( VREG_27_9 ) : ( VREG_27_9 ) ;
assign n44883 =  ( n157 ) ? ( n44881 ) : ( n44882 ) ;
assign n44884 =  ( n6 ) ? ( n44868 ) : ( n44883 ) ;
assign n44885 =  ( n615 ) ? ( n44884 ) : ( VREG_27_9 ) ;
assign n44886 =  ( n148 ) ? ( n1924 ) : ( VREG_28_0 ) ;
assign n44887 =  ( n146 ) ? ( n1923 ) : ( n44886 ) ;
assign n44888 =  ( n144 ) ? ( n1922 ) : ( n44887 ) ;
assign n44889 =  ( n142 ) ? ( n1921 ) : ( n44888 ) ;
assign n44890 =  ( n10 ) ? ( n1920 ) : ( n44889 ) ;
assign n44891 =  ( n148 ) ? ( n2959 ) : ( VREG_28_0 ) ;
assign n44892 =  ( n146 ) ? ( n2958 ) : ( n44891 ) ;
assign n44893 =  ( n144 ) ? ( n2957 ) : ( n44892 ) ;
assign n44894 =  ( n142 ) ? ( n2956 ) : ( n44893 ) ;
assign n44895 =  ( n10 ) ? ( n2955 ) : ( n44894 ) ;
assign n44896 =  ( n3032 ) ? ( VREG_28_0 ) : ( n44890 ) ;
assign n44897 =  ( n3032 ) ? ( VREG_28_0 ) : ( n44895 ) ;
assign n44898 =  ( n3034 ) ? ( n44897 ) : ( VREG_28_0 ) ;
assign n44899 =  ( n2965 ) ? ( n44896 ) : ( n44898 ) ;
assign n44900 =  ( n1930 ) ? ( n44895 ) : ( n44899 ) ;
assign n44901 =  ( n879 ) ? ( n44890 ) : ( n44900 ) ;
assign n44902 =  ( n172 ) ? ( n3045 ) : ( VREG_28_0 ) ;
assign n44903 =  ( n170 ) ? ( n3044 ) : ( n44902 ) ;
assign n44904 =  ( n168 ) ? ( n3043 ) : ( n44903 ) ;
assign n44905 =  ( n166 ) ? ( n3042 ) : ( n44904 ) ;
assign n44906 =  ( n162 ) ? ( n3041 ) : ( n44905 ) ;
assign n44907 =  ( n172 ) ? ( n3056 ) : ( VREG_28_0 ) ;
assign n44908 =  ( n170 ) ? ( n3055 ) : ( n44907 ) ;
assign n44909 =  ( n168 ) ? ( n3054 ) : ( n44908 ) ;
assign n44910 =  ( n166 ) ? ( n3053 ) : ( n44909 ) ;
assign n44911 =  ( n162 ) ? ( n3052 ) : ( n44910 ) ;
assign n44912 =  ( n3032 ) ? ( VREG_28_0 ) : ( n44911 ) ;
assign n44913 =  ( n3051 ) ? ( n44912 ) : ( VREG_28_0 ) ;
assign n44914 =  ( n3040 ) ? ( n44906 ) : ( n44913 ) ;
assign n44915 =  ( n192 ) ? ( VREG_28_0 ) : ( VREG_28_0 ) ;
assign n44916 =  ( n157 ) ? ( n44914 ) : ( n44915 ) ;
assign n44917 =  ( n6 ) ? ( n44901 ) : ( n44916 ) ;
assign n44918 =  ( n637 ) ? ( n44917 ) : ( VREG_28_0 ) ;
assign n44919 =  ( n148 ) ? ( n4113 ) : ( VREG_28_1 ) ;
assign n44920 =  ( n146 ) ? ( n4112 ) : ( n44919 ) ;
assign n44921 =  ( n144 ) ? ( n4111 ) : ( n44920 ) ;
assign n44922 =  ( n142 ) ? ( n4110 ) : ( n44921 ) ;
assign n44923 =  ( n10 ) ? ( n4109 ) : ( n44922 ) ;
assign n44924 =  ( n148 ) ? ( n5147 ) : ( VREG_28_1 ) ;
assign n44925 =  ( n146 ) ? ( n5146 ) : ( n44924 ) ;
assign n44926 =  ( n144 ) ? ( n5145 ) : ( n44925 ) ;
assign n44927 =  ( n142 ) ? ( n5144 ) : ( n44926 ) ;
assign n44928 =  ( n10 ) ? ( n5143 ) : ( n44927 ) ;
assign n44929 =  ( n5154 ) ? ( VREG_28_1 ) : ( n44923 ) ;
assign n44930 =  ( n5154 ) ? ( VREG_28_1 ) : ( n44928 ) ;
assign n44931 =  ( n3034 ) ? ( n44930 ) : ( VREG_28_1 ) ;
assign n44932 =  ( n2965 ) ? ( n44929 ) : ( n44931 ) ;
assign n44933 =  ( n1930 ) ? ( n44928 ) : ( n44932 ) ;
assign n44934 =  ( n879 ) ? ( n44923 ) : ( n44933 ) ;
assign n44935 =  ( n172 ) ? ( n5165 ) : ( VREG_28_1 ) ;
assign n44936 =  ( n170 ) ? ( n5164 ) : ( n44935 ) ;
assign n44937 =  ( n168 ) ? ( n5163 ) : ( n44936 ) ;
assign n44938 =  ( n166 ) ? ( n5162 ) : ( n44937 ) ;
assign n44939 =  ( n162 ) ? ( n5161 ) : ( n44938 ) ;
assign n44940 =  ( n172 ) ? ( n5175 ) : ( VREG_28_1 ) ;
assign n44941 =  ( n170 ) ? ( n5174 ) : ( n44940 ) ;
assign n44942 =  ( n168 ) ? ( n5173 ) : ( n44941 ) ;
assign n44943 =  ( n166 ) ? ( n5172 ) : ( n44942 ) ;
assign n44944 =  ( n162 ) ? ( n5171 ) : ( n44943 ) ;
assign n44945 =  ( n5154 ) ? ( VREG_28_1 ) : ( n44944 ) ;
assign n44946 =  ( n3051 ) ? ( n44945 ) : ( VREG_28_1 ) ;
assign n44947 =  ( n3040 ) ? ( n44939 ) : ( n44946 ) ;
assign n44948 =  ( n192 ) ? ( VREG_28_1 ) : ( VREG_28_1 ) ;
assign n44949 =  ( n157 ) ? ( n44947 ) : ( n44948 ) ;
assign n44950 =  ( n6 ) ? ( n44934 ) : ( n44949 ) ;
assign n44951 =  ( n637 ) ? ( n44950 ) : ( VREG_28_1 ) ;
assign n44952 =  ( n148 ) ? ( n6232 ) : ( VREG_28_10 ) ;
assign n44953 =  ( n146 ) ? ( n6231 ) : ( n44952 ) ;
assign n44954 =  ( n144 ) ? ( n6230 ) : ( n44953 ) ;
assign n44955 =  ( n142 ) ? ( n6229 ) : ( n44954 ) ;
assign n44956 =  ( n10 ) ? ( n6228 ) : ( n44955 ) ;
assign n44957 =  ( n148 ) ? ( n7266 ) : ( VREG_28_10 ) ;
assign n44958 =  ( n146 ) ? ( n7265 ) : ( n44957 ) ;
assign n44959 =  ( n144 ) ? ( n7264 ) : ( n44958 ) ;
assign n44960 =  ( n142 ) ? ( n7263 ) : ( n44959 ) ;
assign n44961 =  ( n10 ) ? ( n7262 ) : ( n44960 ) ;
assign n44962 =  ( n7273 ) ? ( VREG_28_10 ) : ( n44956 ) ;
assign n44963 =  ( n7273 ) ? ( VREG_28_10 ) : ( n44961 ) ;
assign n44964 =  ( n3034 ) ? ( n44963 ) : ( VREG_28_10 ) ;
assign n44965 =  ( n2965 ) ? ( n44962 ) : ( n44964 ) ;
assign n44966 =  ( n1930 ) ? ( n44961 ) : ( n44965 ) ;
assign n44967 =  ( n879 ) ? ( n44956 ) : ( n44966 ) ;
assign n44968 =  ( n172 ) ? ( n7284 ) : ( VREG_28_10 ) ;
assign n44969 =  ( n170 ) ? ( n7283 ) : ( n44968 ) ;
assign n44970 =  ( n168 ) ? ( n7282 ) : ( n44969 ) ;
assign n44971 =  ( n166 ) ? ( n7281 ) : ( n44970 ) ;
assign n44972 =  ( n162 ) ? ( n7280 ) : ( n44971 ) ;
assign n44973 =  ( n172 ) ? ( n7294 ) : ( VREG_28_10 ) ;
assign n44974 =  ( n170 ) ? ( n7293 ) : ( n44973 ) ;
assign n44975 =  ( n168 ) ? ( n7292 ) : ( n44974 ) ;
assign n44976 =  ( n166 ) ? ( n7291 ) : ( n44975 ) ;
assign n44977 =  ( n162 ) ? ( n7290 ) : ( n44976 ) ;
assign n44978 =  ( n7273 ) ? ( VREG_28_10 ) : ( n44977 ) ;
assign n44979 =  ( n3051 ) ? ( n44978 ) : ( VREG_28_10 ) ;
assign n44980 =  ( n3040 ) ? ( n44972 ) : ( n44979 ) ;
assign n44981 =  ( n192 ) ? ( VREG_28_10 ) : ( VREG_28_10 ) ;
assign n44982 =  ( n157 ) ? ( n44980 ) : ( n44981 ) ;
assign n44983 =  ( n6 ) ? ( n44967 ) : ( n44982 ) ;
assign n44984 =  ( n637 ) ? ( n44983 ) : ( VREG_28_10 ) ;
assign n44985 =  ( n148 ) ? ( n8351 ) : ( VREG_28_11 ) ;
assign n44986 =  ( n146 ) ? ( n8350 ) : ( n44985 ) ;
assign n44987 =  ( n144 ) ? ( n8349 ) : ( n44986 ) ;
assign n44988 =  ( n142 ) ? ( n8348 ) : ( n44987 ) ;
assign n44989 =  ( n10 ) ? ( n8347 ) : ( n44988 ) ;
assign n44990 =  ( n148 ) ? ( n9385 ) : ( VREG_28_11 ) ;
assign n44991 =  ( n146 ) ? ( n9384 ) : ( n44990 ) ;
assign n44992 =  ( n144 ) ? ( n9383 ) : ( n44991 ) ;
assign n44993 =  ( n142 ) ? ( n9382 ) : ( n44992 ) ;
assign n44994 =  ( n10 ) ? ( n9381 ) : ( n44993 ) ;
assign n44995 =  ( n9392 ) ? ( VREG_28_11 ) : ( n44989 ) ;
assign n44996 =  ( n9392 ) ? ( VREG_28_11 ) : ( n44994 ) ;
assign n44997 =  ( n3034 ) ? ( n44996 ) : ( VREG_28_11 ) ;
assign n44998 =  ( n2965 ) ? ( n44995 ) : ( n44997 ) ;
assign n44999 =  ( n1930 ) ? ( n44994 ) : ( n44998 ) ;
assign n45000 =  ( n879 ) ? ( n44989 ) : ( n44999 ) ;
assign n45001 =  ( n172 ) ? ( n9403 ) : ( VREG_28_11 ) ;
assign n45002 =  ( n170 ) ? ( n9402 ) : ( n45001 ) ;
assign n45003 =  ( n168 ) ? ( n9401 ) : ( n45002 ) ;
assign n45004 =  ( n166 ) ? ( n9400 ) : ( n45003 ) ;
assign n45005 =  ( n162 ) ? ( n9399 ) : ( n45004 ) ;
assign n45006 =  ( n172 ) ? ( n9413 ) : ( VREG_28_11 ) ;
assign n45007 =  ( n170 ) ? ( n9412 ) : ( n45006 ) ;
assign n45008 =  ( n168 ) ? ( n9411 ) : ( n45007 ) ;
assign n45009 =  ( n166 ) ? ( n9410 ) : ( n45008 ) ;
assign n45010 =  ( n162 ) ? ( n9409 ) : ( n45009 ) ;
assign n45011 =  ( n9392 ) ? ( VREG_28_11 ) : ( n45010 ) ;
assign n45012 =  ( n3051 ) ? ( n45011 ) : ( VREG_28_11 ) ;
assign n45013 =  ( n3040 ) ? ( n45005 ) : ( n45012 ) ;
assign n45014 =  ( n192 ) ? ( VREG_28_11 ) : ( VREG_28_11 ) ;
assign n45015 =  ( n157 ) ? ( n45013 ) : ( n45014 ) ;
assign n45016 =  ( n6 ) ? ( n45000 ) : ( n45015 ) ;
assign n45017 =  ( n637 ) ? ( n45016 ) : ( VREG_28_11 ) ;
assign n45018 =  ( n148 ) ? ( n10470 ) : ( VREG_28_12 ) ;
assign n45019 =  ( n146 ) ? ( n10469 ) : ( n45018 ) ;
assign n45020 =  ( n144 ) ? ( n10468 ) : ( n45019 ) ;
assign n45021 =  ( n142 ) ? ( n10467 ) : ( n45020 ) ;
assign n45022 =  ( n10 ) ? ( n10466 ) : ( n45021 ) ;
assign n45023 =  ( n148 ) ? ( n11504 ) : ( VREG_28_12 ) ;
assign n45024 =  ( n146 ) ? ( n11503 ) : ( n45023 ) ;
assign n45025 =  ( n144 ) ? ( n11502 ) : ( n45024 ) ;
assign n45026 =  ( n142 ) ? ( n11501 ) : ( n45025 ) ;
assign n45027 =  ( n10 ) ? ( n11500 ) : ( n45026 ) ;
assign n45028 =  ( n11511 ) ? ( VREG_28_12 ) : ( n45022 ) ;
assign n45029 =  ( n11511 ) ? ( VREG_28_12 ) : ( n45027 ) ;
assign n45030 =  ( n3034 ) ? ( n45029 ) : ( VREG_28_12 ) ;
assign n45031 =  ( n2965 ) ? ( n45028 ) : ( n45030 ) ;
assign n45032 =  ( n1930 ) ? ( n45027 ) : ( n45031 ) ;
assign n45033 =  ( n879 ) ? ( n45022 ) : ( n45032 ) ;
assign n45034 =  ( n172 ) ? ( n11522 ) : ( VREG_28_12 ) ;
assign n45035 =  ( n170 ) ? ( n11521 ) : ( n45034 ) ;
assign n45036 =  ( n168 ) ? ( n11520 ) : ( n45035 ) ;
assign n45037 =  ( n166 ) ? ( n11519 ) : ( n45036 ) ;
assign n45038 =  ( n162 ) ? ( n11518 ) : ( n45037 ) ;
assign n45039 =  ( n172 ) ? ( n11532 ) : ( VREG_28_12 ) ;
assign n45040 =  ( n170 ) ? ( n11531 ) : ( n45039 ) ;
assign n45041 =  ( n168 ) ? ( n11530 ) : ( n45040 ) ;
assign n45042 =  ( n166 ) ? ( n11529 ) : ( n45041 ) ;
assign n45043 =  ( n162 ) ? ( n11528 ) : ( n45042 ) ;
assign n45044 =  ( n11511 ) ? ( VREG_28_12 ) : ( n45043 ) ;
assign n45045 =  ( n3051 ) ? ( n45044 ) : ( VREG_28_12 ) ;
assign n45046 =  ( n3040 ) ? ( n45038 ) : ( n45045 ) ;
assign n45047 =  ( n192 ) ? ( VREG_28_12 ) : ( VREG_28_12 ) ;
assign n45048 =  ( n157 ) ? ( n45046 ) : ( n45047 ) ;
assign n45049 =  ( n6 ) ? ( n45033 ) : ( n45048 ) ;
assign n45050 =  ( n637 ) ? ( n45049 ) : ( VREG_28_12 ) ;
assign n45051 =  ( n148 ) ? ( n12589 ) : ( VREG_28_13 ) ;
assign n45052 =  ( n146 ) ? ( n12588 ) : ( n45051 ) ;
assign n45053 =  ( n144 ) ? ( n12587 ) : ( n45052 ) ;
assign n45054 =  ( n142 ) ? ( n12586 ) : ( n45053 ) ;
assign n45055 =  ( n10 ) ? ( n12585 ) : ( n45054 ) ;
assign n45056 =  ( n148 ) ? ( n13623 ) : ( VREG_28_13 ) ;
assign n45057 =  ( n146 ) ? ( n13622 ) : ( n45056 ) ;
assign n45058 =  ( n144 ) ? ( n13621 ) : ( n45057 ) ;
assign n45059 =  ( n142 ) ? ( n13620 ) : ( n45058 ) ;
assign n45060 =  ( n10 ) ? ( n13619 ) : ( n45059 ) ;
assign n45061 =  ( n13630 ) ? ( VREG_28_13 ) : ( n45055 ) ;
assign n45062 =  ( n13630 ) ? ( VREG_28_13 ) : ( n45060 ) ;
assign n45063 =  ( n3034 ) ? ( n45062 ) : ( VREG_28_13 ) ;
assign n45064 =  ( n2965 ) ? ( n45061 ) : ( n45063 ) ;
assign n45065 =  ( n1930 ) ? ( n45060 ) : ( n45064 ) ;
assign n45066 =  ( n879 ) ? ( n45055 ) : ( n45065 ) ;
assign n45067 =  ( n172 ) ? ( n13641 ) : ( VREG_28_13 ) ;
assign n45068 =  ( n170 ) ? ( n13640 ) : ( n45067 ) ;
assign n45069 =  ( n168 ) ? ( n13639 ) : ( n45068 ) ;
assign n45070 =  ( n166 ) ? ( n13638 ) : ( n45069 ) ;
assign n45071 =  ( n162 ) ? ( n13637 ) : ( n45070 ) ;
assign n45072 =  ( n172 ) ? ( n13651 ) : ( VREG_28_13 ) ;
assign n45073 =  ( n170 ) ? ( n13650 ) : ( n45072 ) ;
assign n45074 =  ( n168 ) ? ( n13649 ) : ( n45073 ) ;
assign n45075 =  ( n166 ) ? ( n13648 ) : ( n45074 ) ;
assign n45076 =  ( n162 ) ? ( n13647 ) : ( n45075 ) ;
assign n45077 =  ( n13630 ) ? ( VREG_28_13 ) : ( n45076 ) ;
assign n45078 =  ( n3051 ) ? ( n45077 ) : ( VREG_28_13 ) ;
assign n45079 =  ( n3040 ) ? ( n45071 ) : ( n45078 ) ;
assign n45080 =  ( n192 ) ? ( VREG_28_13 ) : ( VREG_28_13 ) ;
assign n45081 =  ( n157 ) ? ( n45079 ) : ( n45080 ) ;
assign n45082 =  ( n6 ) ? ( n45066 ) : ( n45081 ) ;
assign n45083 =  ( n637 ) ? ( n45082 ) : ( VREG_28_13 ) ;
assign n45084 =  ( n148 ) ? ( n14708 ) : ( VREG_28_14 ) ;
assign n45085 =  ( n146 ) ? ( n14707 ) : ( n45084 ) ;
assign n45086 =  ( n144 ) ? ( n14706 ) : ( n45085 ) ;
assign n45087 =  ( n142 ) ? ( n14705 ) : ( n45086 ) ;
assign n45088 =  ( n10 ) ? ( n14704 ) : ( n45087 ) ;
assign n45089 =  ( n148 ) ? ( n15742 ) : ( VREG_28_14 ) ;
assign n45090 =  ( n146 ) ? ( n15741 ) : ( n45089 ) ;
assign n45091 =  ( n144 ) ? ( n15740 ) : ( n45090 ) ;
assign n45092 =  ( n142 ) ? ( n15739 ) : ( n45091 ) ;
assign n45093 =  ( n10 ) ? ( n15738 ) : ( n45092 ) ;
assign n45094 =  ( n15749 ) ? ( VREG_28_14 ) : ( n45088 ) ;
assign n45095 =  ( n15749 ) ? ( VREG_28_14 ) : ( n45093 ) ;
assign n45096 =  ( n3034 ) ? ( n45095 ) : ( VREG_28_14 ) ;
assign n45097 =  ( n2965 ) ? ( n45094 ) : ( n45096 ) ;
assign n45098 =  ( n1930 ) ? ( n45093 ) : ( n45097 ) ;
assign n45099 =  ( n879 ) ? ( n45088 ) : ( n45098 ) ;
assign n45100 =  ( n172 ) ? ( n15760 ) : ( VREG_28_14 ) ;
assign n45101 =  ( n170 ) ? ( n15759 ) : ( n45100 ) ;
assign n45102 =  ( n168 ) ? ( n15758 ) : ( n45101 ) ;
assign n45103 =  ( n166 ) ? ( n15757 ) : ( n45102 ) ;
assign n45104 =  ( n162 ) ? ( n15756 ) : ( n45103 ) ;
assign n45105 =  ( n172 ) ? ( n15770 ) : ( VREG_28_14 ) ;
assign n45106 =  ( n170 ) ? ( n15769 ) : ( n45105 ) ;
assign n45107 =  ( n168 ) ? ( n15768 ) : ( n45106 ) ;
assign n45108 =  ( n166 ) ? ( n15767 ) : ( n45107 ) ;
assign n45109 =  ( n162 ) ? ( n15766 ) : ( n45108 ) ;
assign n45110 =  ( n15749 ) ? ( VREG_28_14 ) : ( n45109 ) ;
assign n45111 =  ( n3051 ) ? ( n45110 ) : ( VREG_28_14 ) ;
assign n45112 =  ( n3040 ) ? ( n45104 ) : ( n45111 ) ;
assign n45113 =  ( n192 ) ? ( VREG_28_14 ) : ( VREG_28_14 ) ;
assign n45114 =  ( n157 ) ? ( n45112 ) : ( n45113 ) ;
assign n45115 =  ( n6 ) ? ( n45099 ) : ( n45114 ) ;
assign n45116 =  ( n637 ) ? ( n45115 ) : ( VREG_28_14 ) ;
assign n45117 =  ( n148 ) ? ( n16827 ) : ( VREG_28_15 ) ;
assign n45118 =  ( n146 ) ? ( n16826 ) : ( n45117 ) ;
assign n45119 =  ( n144 ) ? ( n16825 ) : ( n45118 ) ;
assign n45120 =  ( n142 ) ? ( n16824 ) : ( n45119 ) ;
assign n45121 =  ( n10 ) ? ( n16823 ) : ( n45120 ) ;
assign n45122 =  ( n148 ) ? ( n17861 ) : ( VREG_28_15 ) ;
assign n45123 =  ( n146 ) ? ( n17860 ) : ( n45122 ) ;
assign n45124 =  ( n144 ) ? ( n17859 ) : ( n45123 ) ;
assign n45125 =  ( n142 ) ? ( n17858 ) : ( n45124 ) ;
assign n45126 =  ( n10 ) ? ( n17857 ) : ( n45125 ) ;
assign n45127 =  ( n17868 ) ? ( VREG_28_15 ) : ( n45121 ) ;
assign n45128 =  ( n17868 ) ? ( VREG_28_15 ) : ( n45126 ) ;
assign n45129 =  ( n3034 ) ? ( n45128 ) : ( VREG_28_15 ) ;
assign n45130 =  ( n2965 ) ? ( n45127 ) : ( n45129 ) ;
assign n45131 =  ( n1930 ) ? ( n45126 ) : ( n45130 ) ;
assign n45132 =  ( n879 ) ? ( n45121 ) : ( n45131 ) ;
assign n45133 =  ( n172 ) ? ( n17879 ) : ( VREG_28_15 ) ;
assign n45134 =  ( n170 ) ? ( n17878 ) : ( n45133 ) ;
assign n45135 =  ( n168 ) ? ( n17877 ) : ( n45134 ) ;
assign n45136 =  ( n166 ) ? ( n17876 ) : ( n45135 ) ;
assign n45137 =  ( n162 ) ? ( n17875 ) : ( n45136 ) ;
assign n45138 =  ( n172 ) ? ( n17889 ) : ( VREG_28_15 ) ;
assign n45139 =  ( n170 ) ? ( n17888 ) : ( n45138 ) ;
assign n45140 =  ( n168 ) ? ( n17887 ) : ( n45139 ) ;
assign n45141 =  ( n166 ) ? ( n17886 ) : ( n45140 ) ;
assign n45142 =  ( n162 ) ? ( n17885 ) : ( n45141 ) ;
assign n45143 =  ( n17868 ) ? ( VREG_28_15 ) : ( n45142 ) ;
assign n45144 =  ( n3051 ) ? ( n45143 ) : ( VREG_28_15 ) ;
assign n45145 =  ( n3040 ) ? ( n45137 ) : ( n45144 ) ;
assign n45146 =  ( n192 ) ? ( VREG_28_15 ) : ( VREG_28_15 ) ;
assign n45147 =  ( n157 ) ? ( n45145 ) : ( n45146 ) ;
assign n45148 =  ( n6 ) ? ( n45132 ) : ( n45147 ) ;
assign n45149 =  ( n637 ) ? ( n45148 ) : ( VREG_28_15 ) ;
assign n45150 =  ( n148 ) ? ( n18946 ) : ( VREG_28_2 ) ;
assign n45151 =  ( n146 ) ? ( n18945 ) : ( n45150 ) ;
assign n45152 =  ( n144 ) ? ( n18944 ) : ( n45151 ) ;
assign n45153 =  ( n142 ) ? ( n18943 ) : ( n45152 ) ;
assign n45154 =  ( n10 ) ? ( n18942 ) : ( n45153 ) ;
assign n45155 =  ( n148 ) ? ( n19980 ) : ( VREG_28_2 ) ;
assign n45156 =  ( n146 ) ? ( n19979 ) : ( n45155 ) ;
assign n45157 =  ( n144 ) ? ( n19978 ) : ( n45156 ) ;
assign n45158 =  ( n142 ) ? ( n19977 ) : ( n45157 ) ;
assign n45159 =  ( n10 ) ? ( n19976 ) : ( n45158 ) ;
assign n45160 =  ( n19987 ) ? ( VREG_28_2 ) : ( n45154 ) ;
assign n45161 =  ( n19987 ) ? ( VREG_28_2 ) : ( n45159 ) ;
assign n45162 =  ( n3034 ) ? ( n45161 ) : ( VREG_28_2 ) ;
assign n45163 =  ( n2965 ) ? ( n45160 ) : ( n45162 ) ;
assign n45164 =  ( n1930 ) ? ( n45159 ) : ( n45163 ) ;
assign n45165 =  ( n879 ) ? ( n45154 ) : ( n45164 ) ;
assign n45166 =  ( n172 ) ? ( n19998 ) : ( VREG_28_2 ) ;
assign n45167 =  ( n170 ) ? ( n19997 ) : ( n45166 ) ;
assign n45168 =  ( n168 ) ? ( n19996 ) : ( n45167 ) ;
assign n45169 =  ( n166 ) ? ( n19995 ) : ( n45168 ) ;
assign n45170 =  ( n162 ) ? ( n19994 ) : ( n45169 ) ;
assign n45171 =  ( n172 ) ? ( n20008 ) : ( VREG_28_2 ) ;
assign n45172 =  ( n170 ) ? ( n20007 ) : ( n45171 ) ;
assign n45173 =  ( n168 ) ? ( n20006 ) : ( n45172 ) ;
assign n45174 =  ( n166 ) ? ( n20005 ) : ( n45173 ) ;
assign n45175 =  ( n162 ) ? ( n20004 ) : ( n45174 ) ;
assign n45176 =  ( n19987 ) ? ( VREG_28_2 ) : ( n45175 ) ;
assign n45177 =  ( n3051 ) ? ( n45176 ) : ( VREG_28_2 ) ;
assign n45178 =  ( n3040 ) ? ( n45170 ) : ( n45177 ) ;
assign n45179 =  ( n192 ) ? ( VREG_28_2 ) : ( VREG_28_2 ) ;
assign n45180 =  ( n157 ) ? ( n45178 ) : ( n45179 ) ;
assign n45181 =  ( n6 ) ? ( n45165 ) : ( n45180 ) ;
assign n45182 =  ( n637 ) ? ( n45181 ) : ( VREG_28_2 ) ;
assign n45183 =  ( n148 ) ? ( n21065 ) : ( VREG_28_3 ) ;
assign n45184 =  ( n146 ) ? ( n21064 ) : ( n45183 ) ;
assign n45185 =  ( n144 ) ? ( n21063 ) : ( n45184 ) ;
assign n45186 =  ( n142 ) ? ( n21062 ) : ( n45185 ) ;
assign n45187 =  ( n10 ) ? ( n21061 ) : ( n45186 ) ;
assign n45188 =  ( n148 ) ? ( n22099 ) : ( VREG_28_3 ) ;
assign n45189 =  ( n146 ) ? ( n22098 ) : ( n45188 ) ;
assign n45190 =  ( n144 ) ? ( n22097 ) : ( n45189 ) ;
assign n45191 =  ( n142 ) ? ( n22096 ) : ( n45190 ) ;
assign n45192 =  ( n10 ) ? ( n22095 ) : ( n45191 ) ;
assign n45193 =  ( n22106 ) ? ( VREG_28_3 ) : ( n45187 ) ;
assign n45194 =  ( n22106 ) ? ( VREG_28_3 ) : ( n45192 ) ;
assign n45195 =  ( n3034 ) ? ( n45194 ) : ( VREG_28_3 ) ;
assign n45196 =  ( n2965 ) ? ( n45193 ) : ( n45195 ) ;
assign n45197 =  ( n1930 ) ? ( n45192 ) : ( n45196 ) ;
assign n45198 =  ( n879 ) ? ( n45187 ) : ( n45197 ) ;
assign n45199 =  ( n172 ) ? ( n22117 ) : ( VREG_28_3 ) ;
assign n45200 =  ( n170 ) ? ( n22116 ) : ( n45199 ) ;
assign n45201 =  ( n168 ) ? ( n22115 ) : ( n45200 ) ;
assign n45202 =  ( n166 ) ? ( n22114 ) : ( n45201 ) ;
assign n45203 =  ( n162 ) ? ( n22113 ) : ( n45202 ) ;
assign n45204 =  ( n172 ) ? ( n22127 ) : ( VREG_28_3 ) ;
assign n45205 =  ( n170 ) ? ( n22126 ) : ( n45204 ) ;
assign n45206 =  ( n168 ) ? ( n22125 ) : ( n45205 ) ;
assign n45207 =  ( n166 ) ? ( n22124 ) : ( n45206 ) ;
assign n45208 =  ( n162 ) ? ( n22123 ) : ( n45207 ) ;
assign n45209 =  ( n22106 ) ? ( VREG_28_3 ) : ( n45208 ) ;
assign n45210 =  ( n3051 ) ? ( n45209 ) : ( VREG_28_3 ) ;
assign n45211 =  ( n3040 ) ? ( n45203 ) : ( n45210 ) ;
assign n45212 =  ( n192 ) ? ( VREG_28_3 ) : ( VREG_28_3 ) ;
assign n45213 =  ( n157 ) ? ( n45211 ) : ( n45212 ) ;
assign n45214 =  ( n6 ) ? ( n45198 ) : ( n45213 ) ;
assign n45215 =  ( n637 ) ? ( n45214 ) : ( VREG_28_3 ) ;
assign n45216 =  ( n148 ) ? ( n23184 ) : ( VREG_28_4 ) ;
assign n45217 =  ( n146 ) ? ( n23183 ) : ( n45216 ) ;
assign n45218 =  ( n144 ) ? ( n23182 ) : ( n45217 ) ;
assign n45219 =  ( n142 ) ? ( n23181 ) : ( n45218 ) ;
assign n45220 =  ( n10 ) ? ( n23180 ) : ( n45219 ) ;
assign n45221 =  ( n148 ) ? ( n24218 ) : ( VREG_28_4 ) ;
assign n45222 =  ( n146 ) ? ( n24217 ) : ( n45221 ) ;
assign n45223 =  ( n144 ) ? ( n24216 ) : ( n45222 ) ;
assign n45224 =  ( n142 ) ? ( n24215 ) : ( n45223 ) ;
assign n45225 =  ( n10 ) ? ( n24214 ) : ( n45224 ) ;
assign n45226 =  ( n24225 ) ? ( VREG_28_4 ) : ( n45220 ) ;
assign n45227 =  ( n24225 ) ? ( VREG_28_4 ) : ( n45225 ) ;
assign n45228 =  ( n3034 ) ? ( n45227 ) : ( VREG_28_4 ) ;
assign n45229 =  ( n2965 ) ? ( n45226 ) : ( n45228 ) ;
assign n45230 =  ( n1930 ) ? ( n45225 ) : ( n45229 ) ;
assign n45231 =  ( n879 ) ? ( n45220 ) : ( n45230 ) ;
assign n45232 =  ( n172 ) ? ( n24236 ) : ( VREG_28_4 ) ;
assign n45233 =  ( n170 ) ? ( n24235 ) : ( n45232 ) ;
assign n45234 =  ( n168 ) ? ( n24234 ) : ( n45233 ) ;
assign n45235 =  ( n166 ) ? ( n24233 ) : ( n45234 ) ;
assign n45236 =  ( n162 ) ? ( n24232 ) : ( n45235 ) ;
assign n45237 =  ( n172 ) ? ( n24246 ) : ( VREG_28_4 ) ;
assign n45238 =  ( n170 ) ? ( n24245 ) : ( n45237 ) ;
assign n45239 =  ( n168 ) ? ( n24244 ) : ( n45238 ) ;
assign n45240 =  ( n166 ) ? ( n24243 ) : ( n45239 ) ;
assign n45241 =  ( n162 ) ? ( n24242 ) : ( n45240 ) ;
assign n45242 =  ( n24225 ) ? ( VREG_28_4 ) : ( n45241 ) ;
assign n45243 =  ( n3051 ) ? ( n45242 ) : ( VREG_28_4 ) ;
assign n45244 =  ( n3040 ) ? ( n45236 ) : ( n45243 ) ;
assign n45245 =  ( n192 ) ? ( VREG_28_4 ) : ( VREG_28_4 ) ;
assign n45246 =  ( n157 ) ? ( n45244 ) : ( n45245 ) ;
assign n45247 =  ( n6 ) ? ( n45231 ) : ( n45246 ) ;
assign n45248 =  ( n637 ) ? ( n45247 ) : ( VREG_28_4 ) ;
assign n45249 =  ( n148 ) ? ( n25303 ) : ( VREG_28_5 ) ;
assign n45250 =  ( n146 ) ? ( n25302 ) : ( n45249 ) ;
assign n45251 =  ( n144 ) ? ( n25301 ) : ( n45250 ) ;
assign n45252 =  ( n142 ) ? ( n25300 ) : ( n45251 ) ;
assign n45253 =  ( n10 ) ? ( n25299 ) : ( n45252 ) ;
assign n45254 =  ( n148 ) ? ( n26337 ) : ( VREG_28_5 ) ;
assign n45255 =  ( n146 ) ? ( n26336 ) : ( n45254 ) ;
assign n45256 =  ( n144 ) ? ( n26335 ) : ( n45255 ) ;
assign n45257 =  ( n142 ) ? ( n26334 ) : ( n45256 ) ;
assign n45258 =  ( n10 ) ? ( n26333 ) : ( n45257 ) ;
assign n45259 =  ( n26344 ) ? ( VREG_28_5 ) : ( n45253 ) ;
assign n45260 =  ( n26344 ) ? ( VREG_28_5 ) : ( n45258 ) ;
assign n45261 =  ( n3034 ) ? ( n45260 ) : ( VREG_28_5 ) ;
assign n45262 =  ( n2965 ) ? ( n45259 ) : ( n45261 ) ;
assign n45263 =  ( n1930 ) ? ( n45258 ) : ( n45262 ) ;
assign n45264 =  ( n879 ) ? ( n45253 ) : ( n45263 ) ;
assign n45265 =  ( n172 ) ? ( n26355 ) : ( VREG_28_5 ) ;
assign n45266 =  ( n170 ) ? ( n26354 ) : ( n45265 ) ;
assign n45267 =  ( n168 ) ? ( n26353 ) : ( n45266 ) ;
assign n45268 =  ( n166 ) ? ( n26352 ) : ( n45267 ) ;
assign n45269 =  ( n162 ) ? ( n26351 ) : ( n45268 ) ;
assign n45270 =  ( n172 ) ? ( n26365 ) : ( VREG_28_5 ) ;
assign n45271 =  ( n170 ) ? ( n26364 ) : ( n45270 ) ;
assign n45272 =  ( n168 ) ? ( n26363 ) : ( n45271 ) ;
assign n45273 =  ( n166 ) ? ( n26362 ) : ( n45272 ) ;
assign n45274 =  ( n162 ) ? ( n26361 ) : ( n45273 ) ;
assign n45275 =  ( n26344 ) ? ( VREG_28_5 ) : ( n45274 ) ;
assign n45276 =  ( n3051 ) ? ( n45275 ) : ( VREG_28_5 ) ;
assign n45277 =  ( n3040 ) ? ( n45269 ) : ( n45276 ) ;
assign n45278 =  ( n192 ) ? ( VREG_28_5 ) : ( VREG_28_5 ) ;
assign n45279 =  ( n157 ) ? ( n45277 ) : ( n45278 ) ;
assign n45280 =  ( n6 ) ? ( n45264 ) : ( n45279 ) ;
assign n45281 =  ( n637 ) ? ( n45280 ) : ( VREG_28_5 ) ;
assign n45282 =  ( n148 ) ? ( n27422 ) : ( VREG_28_6 ) ;
assign n45283 =  ( n146 ) ? ( n27421 ) : ( n45282 ) ;
assign n45284 =  ( n144 ) ? ( n27420 ) : ( n45283 ) ;
assign n45285 =  ( n142 ) ? ( n27419 ) : ( n45284 ) ;
assign n45286 =  ( n10 ) ? ( n27418 ) : ( n45285 ) ;
assign n45287 =  ( n148 ) ? ( n28456 ) : ( VREG_28_6 ) ;
assign n45288 =  ( n146 ) ? ( n28455 ) : ( n45287 ) ;
assign n45289 =  ( n144 ) ? ( n28454 ) : ( n45288 ) ;
assign n45290 =  ( n142 ) ? ( n28453 ) : ( n45289 ) ;
assign n45291 =  ( n10 ) ? ( n28452 ) : ( n45290 ) ;
assign n45292 =  ( n28463 ) ? ( VREG_28_6 ) : ( n45286 ) ;
assign n45293 =  ( n28463 ) ? ( VREG_28_6 ) : ( n45291 ) ;
assign n45294 =  ( n3034 ) ? ( n45293 ) : ( VREG_28_6 ) ;
assign n45295 =  ( n2965 ) ? ( n45292 ) : ( n45294 ) ;
assign n45296 =  ( n1930 ) ? ( n45291 ) : ( n45295 ) ;
assign n45297 =  ( n879 ) ? ( n45286 ) : ( n45296 ) ;
assign n45298 =  ( n172 ) ? ( n28474 ) : ( VREG_28_6 ) ;
assign n45299 =  ( n170 ) ? ( n28473 ) : ( n45298 ) ;
assign n45300 =  ( n168 ) ? ( n28472 ) : ( n45299 ) ;
assign n45301 =  ( n166 ) ? ( n28471 ) : ( n45300 ) ;
assign n45302 =  ( n162 ) ? ( n28470 ) : ( n45301 ) ;
assign n45303 =  ( n172 ) ? ( n28484 ) : ( VREG_28_6 ) ;
assign n45304 =  ( n170 ) ? ( n28483 ) : ( n45303 ) ;
assign n45305 =  ( n168 ) ? ( n28482 ) : ( n45304 ) ;
assign n45306 =  ( n166 ) ? ( n28481 ) : ( n45305 ) ;
assign n45307 =  ( n162 ) ? ( n28480 ) : ( n45306 ) ;
assign n45308 =  ( n28463 ) ? ( VREG_28_6 ) : ( n45307 ) ;
assign n45309 =  ( n3051 ) ? ( n45308 ) : ( VREG_28_6 ) ;
assign n45310 =  ( n3040 ) ? ( n45302 ) : ( n45309 ) ;
assign n45311 =  ( n192 ) ? ( VREG_28_6 ) : ( VREG_28_6 ) ;
assign n45312 =  ( n157 ) ? ( n45310 ) : ( n45311 ) ;
assign n45313 =  ( n6 ) ? ( n45297 ) : ( n45312 ) ;
assign n45314 =  ( n637 ) ? ( n45313 ) : ( VREG_28_6 ) ;
assign n45315 =  ( n148 ) ? ( n29541 ) : ( VREG_28_7 ) ;
assign n45316 =  ( n146 ) ? ( n29540 ) : ( n45315 ) ;
assign n45317 =  ( n144 ) ? ( n29539 ) : ( n45316 ) ;
assign n45318 =  ( n142 ) ? ( n29538 ) : ( n45317 ) ;
assign n45319 =  ( n10 ) ? ( n29537 ) : ( n45318 ) ;
assign n45320 =  ( n148 ) ? ( n30575 ) : ( VREG_28_7 ) ;
assign n45321 =  ( n146 ) ? ( n30574 ) : ( n45320 ) ;
assign n45322 =  ( n144 ) ? ( n30573 ) : ( n45321 ) ;
assign n45323 =  ( n142 ) ? ( n30572 ) : ( n45322 ) ;
assign n45324 =  ( n10 ) ? ( n30571 ) : ( n45323 ) ;
assign n45325 =  ( n30582 ) ? ( VREG_28_7 ) : ( n45319 ) ;
assign n45326 =  ( n30582 ) ? ( VREG_28_7 ) : ( n45324 ) ;
assign n45327 =  ( n3034 ) ? ( n45326 ) : ( VREG_28_7 ) ;
assign n45328 =  ( n2965 ) ? ( n45325 ) : ( n45327 ) ;
assign n45329 =  ( n1930 ) ? ( n45324 ) : ( n45328 ) ;
assign n45330 =  ( n879 ) ? ( n45319 ) : ( n45329 ) ;
assign n45331 =  ( n172 ) ? ( n30593 ) : ( VREG_28_7 ) ;
assign n45332 =  ( n170 ) ? ( n30592 ) : ( n45331 ) ;
assign n45333 =  ( n168 ) ? ( n30591 ) : ( n45332 ) ;
assign n45334 =  ( n166 ) ? ( n30590 ) : ( n45333 ) ;
assign n45335 =  ( n162 ) ? ( n30589 ) : ( n45334 ) ;
assign n45336 =  ( n172 ) ? ( n30603 ) : ( VREG_28_7 ) ;
assign n45337 =  ( n170 ) ? ( n30602 ) : ( n45336 ) ;
assign n45338 =  ( n168 ) ? ( n30601 ) : ( n45337 ) ;
assign n45339 =  ( n166 ) ? ( n30600 ) : ( n45338 ) ;
assign n45340 =  ( n162 ) ? ( n30599 ) : ( n45339 ) ;
assign n45341 =  ( n30582 ) ? ( VREG_28_7 ) : ( n45340 ) ;
assign n45342 =  ( n3051 ) ? ( n45341 ) : ( VREG_28_7 ) ;
assign n45343 =  ( n3040 ) ? ( n45335 ) : ( n45342 ) ;
assign n45344 =  ( n192 ) ? ( VREG_28_7 ) : ( VREG_28_7 ) ;
assign n45345 =  ( n157 ) ? ( n45343 ) : ( n45344 ) ;
assign n45346 =  ( n6 ) ? ( n45330 ) : ( n45345 ) ;
assign n45347 =  ( n637 ) ? ( n45346 ) : ( VREG_28_7 ) ;
assign n45348 =  ( n148 ) ? ( n31660 ) : ( VREG_28_8 ) ;
assign n45349 =  ( n146 ) ? ( n31659 ) : ( n45348 ) ;
assign n45350 =  ( n144 ) ? ( n31658 ) : ( n45349 ) ;
assign n45351 =  ( n142 ) ? ( n31657 ) : ( n45350 ) ;
assign n45352 =  ( n10 ) ? ( n31656 ) : ( n45351 ) ;
assign n45353 =  ( n148 ) ? ( n32694 ) : ( VREG_28_8 ) ;
assign n45354 =  ( n146 ) ? ( n32693 ) : ( n45353 ) ;
assign n45355 =  ( n144 ) ? ( n32692 ) : ( n45354 ) ;
assign n45356 =  ( n142 ) ? ( n32691 ) : ( n45355 ) ;
assign n45357 =  ( n10 ) ? ( n32690 ) : ( n45356 ) ;
assign n45358 =  ( n32701 ) ? ( VREG_28_8 ) : ( n45352 ) ;
assign n45359 =  ( n32701 ) ? ( VREG_28_8 ) : ( n45357 ) ;
assign n45360 =  ( n3034 ) ? ( n45359 ) : ( VREG_28_8 ) ;
assign n45361 =  ( n2965 ) ? ( n45358 ) : ( n45360 ) ;
assign n45362 =  ( n1930 ) ? ( n45357 ) : ( n45361 ) ;
assign n45363 =  ( n879 ) ? ( n45352 ) : ( n45362 ) ;
assign n45364 =  ( n172 ) ? ( n32712 ) : ( VREG_28_8 ) ;
assign n45365 =  ( n170 ) ? ( n32711 ) : ( n45364 ) ;
assign n45366 =  ( n168 ) ? ( n32710 ) : ( n45365 ) ;
assign n45367 =  ( n166 ) ? ( n32709 ) : ( n45366 ) ;
assign n45368 =  ( n162 ) ? ( n32708 ) : ( n45367 ) ;
assign n45369 =  ( n172 ) ? ( n32722 ) : ( VREG_28_8 ) ;
assign n45370 =  ( n170 ) ? ( n32721 ) : ( n45369 ) ;
assign n45371 =  ( n168 ) ? ( n32720 ) : ( n45370 ) ;
assign n45372 =  ( n166 ) ? ( n32719 ) : ( n45371 ) ;
assign n45373 =  ( n162 ) ? ( n32718 ) : ( n45372 ) ;
assign n45374 =  ( n32701 ) ? ( VREG_28_8 ) : ( n45373 ) ;
assign n45375 =  ( n3051 ) ? ( n45374 ) : ( VREG_28_8 ) ;
assign n45376 =  ( n3040 ) ? ( n45368 ) : ( n45375 ) ;
assign n45377 =  ( n192 ) ? ( VREG_28_8 ) : ( VREG_28_8 ) ;
assign n45378 =  ( n157 ) ? ( n45376 ) : ( n45377 ) ;
assign n45379 =  ( n6 ) ? ( n45363 ) : ( n45378 ) ;
assign n45380 =  ( n637 ) ? ( n45379 ) : ( VREG_28_8 ) ;
assign n45381 =  ( n148 ) ? ( n33779 ) : ( VREG_28_9 ) ;
assign n45382 =  ( n146 ) ? ( n33778 ) : ( n45381 ) ;
assign n45383 =  ( n144 ) ? ( n33777 ) : ( n45382 ) ;
assign n45384 =  ( n142 ) ? ( n33776 ) : ( n45383 ) ;
assign n45385 =  ( n10 ) ? ( n33775 ) : ( n45384 ) ;
assign n45386 =  ( n148 ) ? ( n34813 ) : ( VREG_28_9 ) ;
assign n45387 =  ( n146 ) ? ( n34812 ) : ( n45386 ) ;
assign n45388 =  ( n144 ) ? ( n34811 ) : ( n45387 ) ;
assign n45389 =  ( n142 ) ? ( n34810 ) : ( n45388 ) ;
assign n45390 =  ( n10 ) ? ( n34809 ) : ( n45389 ) ;
assign n45391 =  ( n34820 ) ? ( VREG_28_9 ) : ( n45385 ) ;
assign n45392 =  ( n34820 ) ? ( VREG_28_9 ) : ( n45390 ) ;
assign n45393 =  ( n3034 ) ? ( n45392 ) : ( VREG_28_9 ) ;
assign n45394 =  ( n2965 ) ? ( n45391 ) : ( n45393 ) ;
assign n45395 =  ( n1930 ) ? ( n45390 ) : ( n45394 ) ;
assign n45396 =  ( n879 ) ? ( n45385 ) : ( n45395 ) ;
assign n45397 =  ( n172 ) ? ( n34831 ) : ( VREG_28_9 ) ;
assign n45398 =  ( n170 ) ? ( n34830 ) : ( n45397 ) ;
assign n45399 =  ( n168 ) ? ( n34829 ) : ( n45398 ) ;
assign n45400 =  ( n166 ) ? ( n34828 ) : ( n45399 ) ;
assign n45401 =  ( n162 ) ? ( n34827 ) : ( n45400 ) ;
assign n45402 =  ( n172 ) ? ( n34841 ) : ( VREG_28_9 ) ;
assign n45403 =  ( n170 ) ? ( n34840 ) : ( n45402 ) ;
assign n45404 =  ( n168 ) ? ( n34839 ) : ( n45403 ) ;
assign n45405 =  ( n166 ) ? ( n34838 ) : ( n45404 ) ;
assign n45406 =  ( n162 ) ? ( n34837 ) : ( n45405 ) ;
assign n45407 =  ( n34820 ) ? ( VREG_28_9 ) : ( n45406 ) ;
assign n45408 =  ( n3051 ) ? ( n45407 ) : ( VREG_28_9 ) ;
assign n45409 =  ( n3040 ) ? ( n45401 ) : ( n45408 ) ;
assign n45410 =  ( n192 ) ? ( VREG_28_9 ) : ( VREG_28_9 ) ;
assign n45411 =  ( n157 ) ? ( n45409 ) : ( n45410 ) ;
assign n45412 =  ( n6 ) ? ( n45396 ) : ( n45411 ) ;
assign n45413 =  ( n637 ) ? ( n45412 ) : ( VREG_28_9 ) ;
assign n45414 =  ( n148 ) ? ( n1924 ) : ( VREG_29_0 ) ;
assign n45415 =  ( n146 ) ? ( n1923 ) : ( n45414 ) ;
assign n45416 =  ( n144 ) ? ( n1922 ) : ( n45415 ) ;
assign n45417 =  ( n142 ) ? ( n1921 ) : ( n45416 ) ;
assign n45418 =  ( n10 ) ? ( n1920 ) : ( n45417 ) ;
assign n45419 =  ( n148 ) ? ( n2959 ) : ( VREG_29_0 ) ;
assign n45420 =  ( n146 ) ? ( n2958 ) : ( n45419 ) ;
assign n45421 =  ( n144 ) ? ( n2957 ) : ( n45420 ) ;
assign n45422 =  ( n142 ) ? ( n2956 ) : ( n45421 ) ;
assign n45423 =  ( n10 ) ? ( n2955 ) : ( n45422 ) ;
assign n45424 =  ( n3032 ) ? ( VREG_29_0 ) : ( n45418 ) ;
assign n45425 =  ( n3032 ) ? ( VREG_29_0 ) : ( n45423 ) ;
assign n45426 =  ( n3034 ) ? ( n45425 ) : ( VREG_29_0 ) ;
assign n45427 =  ( n2965 ) ? ( n45424 ) : ( n45426 ) ;
assign n45428 =  ( n1930 ) ? ( n45423 ) : ( n45427 ) ;
assign n45429 =  ( n879 ) ? ( n45418 ) : ( n45428 ) ;
assign n45430 =  ( n172 ) ? ( n3045 ) : ( VREG_29_0 ) ;
assign n45431 =  ( n170 ) ? ( n3044 ) : ( n45430 ) ;
assign n45432 =  ( n168 ) ? ( n3043 ) : ( n45431 ) ;
assign n45433 =  ( n166 ) ? ( n3042 ) : ( n45432 ) ;
assign n45434 =  ( n162 ) ? ( n3041 ) : ( n45433 ) ;
assign n45435 =  ( n172 ) ? ( n3056 ) : ( VREG_29_0 ) ;
assign n45436 =  ( n170 ) ? ( n3055 ) : ( n45435 ) ;
assign n45437 =  ( n168 ) ? ( n3054 ) : ( n45436 ) ;
assign n45438 =  ( n166 ) ? ( n3053 ) : ( n45437 ) ;
assign n45439 =  ( n162 ) ? ( n3052 ) : ( n45438 ) ;
assign n45440 =  ( n3032 ) ? ( VREG_29_0 ) : ( n45439 ) ;
assign n45441 =  ( n3051 ) ? ( n45440 ) : ( VREG_29_0 ) ;
assign n45442 =  ( n3040 ) ? ( n45434 ) : ( n45441 ) ;
assign n45443 =  ( n192 ) ? ( VREG_29_0 ) : ( VREG_29_0 ) ;
assign n45444 =  ( n157 ) ? ( n45442 ) : ( n45443 ) ;
assign n45445 =  ( n6 ) ? ( n45429 ) : ( n45444 ) ;
assign n45446 =  ( n659 ) ? ( n45445 ) : ( VREG_29_0 ) ;
assign n45447 =  ( n148 ) ? ( n4113 ) : ( VREG_29_1 ) ;
assign n45448 =  ( n146 ) ? ( n4112 ) : ( n45447 ) ;
assign n45449 =  ( n144 ) ? ( n4111 ) : ( n45448 ) ;
assign n45450 =  ( n142 ) ? ( n4110 ) : ( n45449 ) ;
assign n45451 =  ( n10 ) ? ( n4109 ) : ( n45450 ) ;
assign n45452 =  ( n148 ) ? ( n5147 ) : ( VREG_29_1 ) ;
assign n45453 =  ( n146 ) ? ( n5146 ) : ( n45452 ) ;
assign n45454 =  ( n144 ) ? ( n5145 ) : ( n45453 ) ;
assign n45455 =  ( n142 ) ? ( n5144 ) : ( n45454 ) ;
assign n45456 =  ( n10 ) ? ( n5143 ) : ( n45455 ) ;
assign n45457 =  ( n5154 ) ? ( VREG_29_1 ) : ( n45451 ) ;
assign n45458 =  ( n5154 ) ? ( VREG_29_1 ) : ( n45456 ) ;
assign n45459 =  ( n3034 ) ? ( n45458 ) : ( VREG_29_1 ) ;
assign n45460 =  ( n2965 ) ? ( n45457 ) : ( n45459 ) ;
assign n45461 =  ( n1930 ) ? ( n45456 ) : ( n45460 ) ;
assign n45462 =  ( n879 ) ? ( n45451 ) : ( n45461 ) ;
assign n45463 =  ( n172 ) ? ( n5165 ) : ( VREG_29_1 ) ;
assign n45464 =  ( n170 ) ? ( n5164 ) : ( n45463 ) ;
assign n45465 =  ( n168 ) ? ( n5163 ) : ( n45464 ) ;
assign n45466 =  ( n166 ) ? ( n5162 ) : ( n45465 ) ;
assign n45467 =  ( n162 ) ? ( n5161 ) : ( n45466 ) ;
assign n45468 =  ( n172 ) ? ( n5175 ) : ( VREG_29_1 ) ;
assign n45469 =  ( n170 ) ? ( n5174 ) : ( n45468 ) ;
assign n45470 =  ( n168 ) ? ( n5173 ) : ( n45469 ) ;
assign n45471 =  ( n166 ) ? ( n5172 ) : ( n45470 ) ;
assign n45472 =  ( n162 ) ? ( n5171 ) : ( n45471 ) ;
assign n45473 =  ( n5154 ) ? ( VREG_29_1 ) : ( n45472 ) ;
assign n45474 =  ( n3051 ) ? ( n45473 ) : ( VREG_29_1 ) ;
assign n45475 =  ( n3040 ) ? ( n45467 ) : ( n45474 ) ;
assign n45476 =  ( n192 ) ? ( VREG_29_1 ) : ( VREG_29_1 ) ;
assign n45477 =  ( n157 ) ? ( n45475 ) : ( n45476 ) ;
assign n45478 =  ( n6 ) ? ( n45462 ) : ( n45477 ) ;
assign n45479 =  ( n659 ) ? ( n45478 ) : ( VREG_29_1 ) ;
assign n45480 =  ( n148 ) ? ( n6232 ) : ( VREG_29_10 ) ;
assign n45481 =  ( n146 ) ? ( n6231 ) : ( n45480 ) ;
assign n45482 =  ( n144 ) ? ( n6230 ) : ( n45481 ) ;
assign n45483 =  ( n142 ) ? ( n6229 ) : ( n45482 ) ;
assign n45484 =  ( n10 ) ? ( n6228 ) : ( n45483 ) ;
assign n45485 =  ( n148 ) ? ( n7266 ) : ( VREG_29_10 ) ;
assign n45486 =  ( n146 ) ? ( n7265 ) : ( n45485 ) ;
assign n45487 =  ( n144 ) ? ( n7264 ) : ( n45486 ) ;
assign n45488 =  ( n142 ) ? ( n7263 ) : ( n45487 ) ;
assign n45489 =  ( n10 ) ? ( n7262 ) : ( n45488 ) ;
assign n45490 =  ( n7273 ) ? ( VREG_29_10 ) : ( n45484 ) ;
assign n45491 =  ( n7273 ) ? ( VREG_29_10 ) : ( n45489 ) ;
assign n45492 =  ( n3034 ) ? ( n45491 ) : ( VREG_29_10 ) ;
assign n45493 =  ( n2965 ) ? ( n45490 ) : ( n45492 ) ;
assign n45494 =  ( n1930 ) ? ( n45489 ) : ( n45493 ) ;
assign n45495 =  ( n879 ) ? ( n45484 ) : ( n45494 ) ;
assign n45496 =  ( n172 ) ? ( n7284 ) : ( VREG_29_10 ) ;
assign n45497 =  ( n170 ) ? ( n7283 ) : ( n45496 ) ;
assign n45498 =  ( n168 ) ? ( n7282 ) : ( n45497 ) ;
assign n45499 =  ( n166 ) ? ( n7281 ) : ( n45498 ) ;
assign n45500 =  ( n162 ) ? ( n7280 ) : ( n45499 ) ;
assign n45501 =  ( n172 ) ? ( n7294 ) : ( VREG_29_10 ) ;
assign n45502 =  ( n170 ) ? ( n7293 ) : ( n45501 ) ;
assign n45503 =  ( n168 ) ? ( n7292 ) : ( n45502 ) ;
assign n45504 =  ( n166 ) ? ( n7291 ) : ( n45503 ) ;
assign n45505 =  ( n162 ) ? ( n7290 ) : ( n45504 ) ;
assign n45506 =  ( n7273 ) ? ( VREG_29_10 ) : ( n45505 ) ;
assign n45507 =  ( n3051 ) ? ( n45506 ) : ( VREG_29_10 ) ;
assign n45508 =  ( n3040 ) ? ( n45500 ) : ( n45507 ) ;
assign n45509 =  ( n192 ) ? ( VREG_29_10 ) : ( VREG_29_10 ) ;
assign n45510 =  ( n157 ) ? ( n45508 ) : ( n45509 ) ;
assign n45511 =  ( n6 ) ? ( n45495 ) : ( n45510 ) ;
assign n45512 =  ( n659 ) ? ( n45511 ) : ( VREG_29_10 ) ;
assign n45513 =  ( n148 ) ? ( n8351 ) : ( VREG_29_11 ) ;
assign n45514 =  ( n146 ) ? ( n8350 ) : ( n45513 ) ;
assign n45515 =  ( n144 ) ? ( n8349 ) : ( n45514 ) ;
assign n45516 =  ( n142 ) ? ( n8348 ) : ( n45515 ) ;
assign n45517 =  ( n10 ) ? ( n8347 ) : ( n45516 ) ;
assign n45518 =  ( n148 ) ? ( n9385 ) : ( VREG_29_11 ) ;
assign n45519 =  ( n146 ) ? ( n9384 ) : ( n45518 ) ;
assign n45520 =  ( n144 ) ? ( n9383 ) : ( n45519 ) ;
assign n45521 =  ( n142 ) ? ( n9382 ) : ( n45520 ) ;
assign n45522 =  ( n10 ) ? ( n9381 ) : ( n45521 ) ;
assign n45523 =  ( n9392 ) ? ( VREG_29_11 ) : ( n45517 ) ;
assign n45524 =  ( n9392 ) ? ( VREG_29_11 ) : ( n45522 ) ;
assign n45525 =  ( n3034 ) ? ( n45524 ) : ( VREG_29_11 ) ;
assign n45526 =  ( n2965 ) ? ( n45523 ) : ( n45525 ) ;
assign n45527 =  ( n1930 ) ? ( n45522 ) : ( n45526 ) ;
assign n45528 =  ( n879 ) ? ( n45517 ) : ( n45527 ) ;
assign n45529 =  ( n172 ) ? ( n9403 ) : ( VREG_29_11 ) ;
assign n45530 =  ( n170 ) ? ( n9402 ) : ( n45529 ) ;
assign n45531 =  ( n168 ) ? ( n9401 ) : ( n45530 ) ;
assign n45532 =  ( n166 ) ? ( n9400 ) : ( n45531 ) ;
assign n45533 =  ( n162 ) ? ( n9399 ) : ( n45532 ) ;
assign n45534 =  ( n172 ) ? ( n9413 ) : ( VREG_29_11 ) ;
assign n45535 =  ( n170 ) ? ( n9412 ) : ( n45534 ) ;
assign n45536 =  ( n168 ) ? ( n9411 ) : ( n45535 ) ;
assign n45537 =  ( n166 ) ? ( n9410 ) : ( n45536 ) ;
assign n45538 =  ( n162 ) ? ( n9409 ) : ( n45537 ) ;
assign n45539 =  ( n9392 ) ? ( VREG_29_11 ) : ( n45538 ) ;
assign n45540 =  ( n3051 ) ? ( n45539 ) : ( VREG_29_11 ) ;
assign n45541 =  ( n3040 ) ? ( n45533 ) : ( n45540 ) ;
assign n45542 =  ( n192 ) ? ( VREG_29_11 ) : ( VREG_29_11 ) ;
assign n45543 =  ( n157 ) ? ( n45541 ) : ( n45542 ) ;
assign n45544 =  ( n6 ) ? ( n45528 ) : ( n45543 ) ;
assign n45545 =  ( n659 ) ? ( n45544 ) : ( VREG_29_11 ) ;
assign n45546 =  ( n148 ) ? ( n10470 ) : ( VREG_29_12 ) ;
assign n45547 =  ( n146 ) ? ( n10469 ) : ( n45546 ) ;
assign n45548 =  ( n144 ) ? ( n10468 ) : ( n45547 ) ;
assign n45549 =  ( n142 ) ? ( n10467 ) : ( n45548 ) ;
assign n45550 =  ( n10 ) ? ( n10466 ) : ( n45549 ) ;
assign n45551 =  ( n148 ) ? ( n11504 ) : ( VREG_29_12 ) ;
assign n45552 =  ( n146 ) ? ( n11503 ) : ( n45551 ) ;
assign n45553 =  ( n144 ) ? ( n11502 ) : ( n45552 ) ;
assign n45554 =  ( n142 ) ? ( n11501 ) : ( n45553 ) ;
assign n45555 =  ( n10 ) ? ( n11500 ) : ( n45554 ) ;
assign n45556 =  ( n11511 ) ? ( VREG_29_12 ) : ( n45550 ) ;
assign n45557 =  ( n11511 ) ? ( VREG_29_12 ) : ( n45555 ) ;
assign n45558 =  ( n3034 ) ? ( n45557 ) : ( VREG_29_12 ) ;
assign n45559 =  ( n2965 ) ? ( n45556 ) : ( n45558 ) ;
assign n45560 =  ( n1930 ) ? ( n45555 ) : ( n45559 ) ;
assign n45561 =  ( n879 ) ? ( n45550 ) : ( n45560 ) ;
assign n45562 =  ( n172 ) ? ( n11522 ) : ( VREG_29_12 ) ;
assign n45563 =  ( n170 ) ? ( n11521 ) : ( n45562 ) ;
assign n45564 =  ( n168 ) ? ( n11520 ) : ( n45563 ) ;
assign n45565 =  ( n166 ) ? ( n11519 ) : ( n45564 ) ;
assign n45566 =  ( n162 ) ? ( n11518 ) : ( n45565 ) ;
assign n45567 =  ( n172 ) ? ( n11532 ) : ( VREG_29_12 ) ;
assign n45568 =  ( n170 ) ? ( n11531 ) : ( n45567 ) ;
assign n45569 =  ( n168 ) ? ( n11530 ) : ( n45568 ) ;
assign n45570 =  ( n166 ) ? ( n11529 ) : ( n45569 ) ;
assign n45571 =  ( n162 ) ? ( n11528 ) : ( n45570 ) ;
assign n45572 =  ( n11511 ) ? ( VREG_29_12 ) : ( n45571 ) ;
assign n45573 =  ( n3051 ) ? ( n45572 ) : ( VREG_29_12 ) ;
assign n45574 =  ( n3040 ) ? ( n45566 ) : ( n45573 ) ;
assign n45575 =  ( n192 ) ? ( VREG_29_12 ) : ( VREG_29_12 ) ;
assign n45576 =  ( n157 ) ? ( n45574 ) : ( n45575 ) ;
assign n45577 =  ( n6 ) ? ( n45561 ) : ( n45576 ) ;
assign n45578 =  ( n659 ) ? ( n45577 ) : ( VREG_29_12 ) ;
assign n45579 =  ( n148 ) ? ( n12589 ) : ( VREG_29_13 ) ;
assign n45580 =  ( n146 ) ? ( n12588 ) : ( n45579 ) ;
assign n45581 =  ( n144 ) ? ( n12587 ) : ( n45580 ) ;
assign n45582 =  ( n142 ) ? ( n12586 ) : ( n45581 ) ;
assign n45583 =  ( n10 ) ? ( n12585 ) : ( n45582 ) ;
assign n45584 =  ( n148 ) ? ( n13623 ) : ( VREG_29_13 ) ;
assign n45585 =  ( n146 ) ? ( n13622 ) : ( n45584 ) ;
assign n45586 =  ( n144 ) ? ( n13621 ) : ( n45585 ) ;
assign n45587 =  ( n142 ) ? ( n13620 ) : ( n45586 ) ;
assign n45588 =  ( n10 ) ? ( n13619 ) : ( n45587 ) ;
assign n45589 =  ( n13630 ) ? ( VREG_29_13 ) : ( n45583 ) ;
assign n45590 =  ( n13630 ) ? ( VREG_29_13 ) : ( n45588 ) ;
assign n45591 =  ( n3034 ) ? ( n45590 ) : ( VREG_29_13 ) ;
assign n45592 =  ( n2965 ) ? ( n45589 ) : ( n45591 ) ;
assign n45593 =  ( n1930 ) ? ( n45588 ) : ( n45592 ) ;
assign n45594 =  ( n879 ) ? ( n45583 ) : ( n45593 ) ;
assign n45595 =  ( n172 ) ? ( n13641 ) : ( VREG_29_13 ) ;
assign n45596 =  ( n170 ) ? ( n13640 ) : ( n45595 ) ;
assign n45597 =  ( n168 ) ? ( n13639 ) : ( n45596 ) ;
assign n45598 =  ( n166 ) ? ( n13638 ) : ( n45597 ) ;
assign n45599 =  ( n162 ) ? ( n13637 ) : ( n45598 ) ;
assign n45600 =  ( n172 ) ? ( n13651 ) : ( VREG_29_13 ) ;
assign n45601 =  ( n170 ) ? ( n13650 ) : ( n45600 ) ;
assign n45602 =  ( n168 ) ? ( n13649 ) : ( n45601 ) ;
assign n45603 =  ( n166 ) ? ( n13648 ) : ( n45602 ) ;
assign n45604 =  ( n162 ) ? ( n13647 ) : ( n45603 ) ;
assign n45605 =  ( n13630 ) ? ( VREG_29_13 ) : ( n45604 ) ;
assign n45606 =  ( n3051 ) ? ( n45605 ) : ( VREG_29_13 ) ;
assign n45607 =  ( n3040 ) ? ( n45599 ) : ( n45606 ) ;
assign n45608 =  ( n192 ) ? ( VREG_29_13 ) : ( VREG_29_13 ) ;
assign n45609 =  ( n157 ) ? ( n45607 ) : ( n45608 ) ;
assign n45610 =  ( n6 ) ? ( n45594 ) : ( n45609 ) ;
assign n45611 =  ( n659 ) ? ( n45610 ) : ( VREG_29_13 ) ;
assign n45612 =  ( n148 ) ? ( n14708 ) : ( VREG_29_14 ) ;
assign n45613 =  ( n146 ) ? ( n14707 ) : ( n45612 ) ;
assign n45614 =  ( n144 ) ? ( n14706 ) : ( n45613 ) ;
assign n45615 =  ( n142 ) ? ( n14705 ) : ( n45614 ) ;
assign n45616 =  ( n10 ) ? ( n14704 ) : ( n45615 ) ;
assign n45617 =  ( n148 ) ? ( n15742 ) : ( VREG_29_14 ) ;
assign n45618 =  ( n146 ) ? ( n15741 ) : ( n45617 ) ;
assign n45619 =  ( n144 ) ? ( n15740 ) : ( n45618 ) ;
assign n45620 =  ( n142 ) ? ( n15739 ) : ( n45619 ) ;
assign n45621 =  ( n10 ) ? ( n15738 ) : ( n45620 ) ;
assign n45622 =  ( n15749 ) ? ( VREG_29_14 ) : ( n45616 ) ;
assign n45623 =  ( n15749 ) ? ( VREG_29_14 ) : ( n45621 ) ;
assign n45624 =  ( n3034 ) ? ( n45623 ) : ( VREG_29_14 ) ;
assign n45625 =  ( n2965 ) ? ( n45622 ) : ( n45624 ) ;
assign n45626 =  ( n1930 ) ? ( n45621 ) : ( n45625 ) ;
assign n45627 =  ( n879 ) ? ( n45616 ) : ( n45626 ) ;
assign n45628 =  ( n172 ) ? ( n15760 ) : ( VREG_29_14 ) ;
assign n45629 =  ( n170 ) ? ( n15759 ) : ( n45628 ) ;
assign n45630 =  ( n168 ) ? ( n15758 ) : ( n45629 ) ;
assign n45631 =  ( n166 ) ? ( n15757 ) : ( n45630 ) ;
assign n45632 =  ( n162 ) ? ( n15756 ) : ( n45631 ) ;
assign n45633 =  ( n172 ) ? ( n15770 ) : ( VREG_29_14 ) ;
assign n45634 =  ( n170 ) ? ( n15769 ) : ( n45633 ) ;
assign n45635 =  ( n168 ) ? ( n15768 ) : ( n45634 ) ;
assign n45636 =  ( n166 ) ? ( n15767 ) : ( n45635 ) ;
assign n45637 =  ( n162 ) ? ( n15766 ) : ( n45636 ) ;
assign n45638 =  ( n15749 ) ? ( VREG_29_14 ) : ( n45637 ) ;
assign n45639 =  ( n3051 ) ? ( n45638 ) : ( VREG_29_14 ) ;
assign n45640 =  ( n3040 ) ? ( n45632 ) : ( n45639 ) ;
assign n45641 =  ( n192 ) ? ( VREG_29_14 ) : ( VREG_29_14 ) ;
assign n45642 =  ( n157 ) ? ( n45640 ) : ( n45641 ) ;
assign n45643 =  ( n6 ) ? ( n45627 ) : ( n45642 ) ;
assign n45644 =  ( n659 ) ? ( n45643 ) : ( VREG_29_14 ) ;
assign n45645 =  ( n148 ) ? ( n16827 ) : ( VREG_29_15 ) ;
assign n45646 =  ( n146 ) ? ( n16826 ) : ( n45645 ) ;
assign n45647 =  ( n144 ) ? ( n16825 ) : ( n45646 ) ;
assign n45648 =  ( n142 ) ? ( n16824 ) : ( n45647 ) ;
assign n45649 =  ( n10 ) ? ( n16823 ) : ( n45648 ) ;
assign n45650 =  ( n148 ) ? ( n17861 ) : ( VREG_29_15 ) ;
assign n45651 =  ( n146 ) ? ( n17860 ) : ( n45650 ) ;
assign n45652 =  ( n144 ) ? ( n17859 ) : ( n45651 ) ;
assign n45653 =  ( n142 ) ? ( n17858 ) : ( n45652 ) ;
assign n45654 =  ( n10 ) ? ( n17857 ) : ( n45653 ) ;
assign n45655 =  ( n17868 ) ? ( VREG_29_15 ) : ( n45649 ) ;
assign n45656 =  ( n17868 ) ? ( VREG_29_15 ) : ( n45654 ) ;
assign n45657 =  ( n3034 ) ? ( n45656 ) : ( VREG_29_15 ) ;
assign n45658 =  ( n2965 ) ? ( n45655 ) : ( n45657 ) ;
assign n45659 =  ( n1930 ) ? ( n45654 ) : ( n45658 ) ;
assign n45660 =  ( n879 ) ? ( n45649 ) : ( n45659 ) ;
assign n45661 =  ( n172 ) ? ( n17879 ) : ( VREG_29_15 ) ;
assign n45662 =  ( n170 ) ? ( n17878 ) : ( n45661 ) ;
assign n45663 =  ( n168 ) ? ( n17877 ) : ( n45662 ) ;
assign n45664 =  ( n166 ) ? ( n17876 ) : ( n45663 ) ;
assign n45665 =  ( n162 ) ? ( n17875 ) : ( n45664 ) ;
assign n45666 =  ( n172 ) ? ( n17889 ) : ( VREG_29_15 ) ;
assign n45667 =  ( n170 ) ? ( n17888 ) : ( n45666 ) ;
assign n45668 =  ( n168 ) ? ( n17887 ) : ( n45667 ) ;
assign n45669 =  ( n166 ) ? ( n17886 ) : ( n45668 ) ;
assign n45670 =  ( n162 ) ? ( n17885 ) : ( n45669 ) ;
assign n45671 =  ( n17868 ) ? ( VREG_29_15 ) : ( n45670 ) ;
assign n45672 =  ( n3051 ) ? ( n45671 ) : ( VREG_29_15 ) ;
assign n45673 =  ( n3040 ) ? ( n45665 ) : ( n45672 ) ;
assign n45674 =  ( n192 ) ? ( VREG_29_15 ) : ( VREG_29_15 ) ;
assign n45675 =  ( n157 ) ? ( n45673 ) : ( n45674 ) ;
assign n45676 =  ( n6 ) ? ( n45660 ) : ( n45675 ) ;
assign n45677 =  ( n659 ) ? ( n45676 ) : ( VREG_29_15 ) ;
assign n45678 =  ( n148 ) ? ( n18946 ) : ( VREG_29_2 ) ;
assign n45679 =  ( n146 ) ? ( n18945 ) : ( n45678 ) ;
assign n45680 =  ( n144 ) ? ( n18944 ) : ( n45679 ) ;
assign n45681 =  ( n142 ) ? ( n18943 ) : ( n45680 ) ;
assign n45682 =  ( n10 ) ? ( n18942 ) : ( n45681 ) ;
assign n45683 =  ( n148 ) ? ( n19980 ) : ( VREG_29_2 ) ;
assign n45684 =  ( n146 ) ? ( n19979 ) : ( n45683 ) ;
assign n45685 =  ( n144 ) ? ( n19978 ) : ( n45684 ) ;
assign n45686 =  ( n142 ) ? ( n19977 ) : ( n45685 ) ;
assign n45687 =  ( n10 ) ? ( n19976 ) : ( n45686 ) ;
assign n45688 =  ( n19987 ) ? ( VREG_29_2 ) : ( n45682 ) ;
assign n45689 =  ( n19987 ) ? ( VREG_29_2 ) : ( n45687 ) ;
assign n45690 =  ( n3034 ) ? ( n45689 ) : ( VREG_29_2 ) ;
assign n45691 =  ( n2965 ) ? ( n45688 ) : ( n45690 ) ;
assign n45692 =  ( n1930 ) ? ( n45687 ) : ( n45691 ) ;
assign n45693 =  ( n879 ) ? ( n45682 ) : ( n45692 ) ;
assign n45694 =  ( n172 ) ? ( n19998 ) : ( VREG_29_2 ) ;
assign n45695 =  ( n170 ) ? ( n19997 ) : ( n45694 ) ;
assign n45696 =  ( n168 ) ? ( n19996 ) : ( n45695 ) ;
assign n45697 =  ( n166 ) ? ( n19995 ) : ( n45696 ) ;
assign n45698 =  ( n162 ) ? ( n19994 ) : ( n45697 ) ;
assign n45699 =  ( n172 ) ? ( n20008 ) : ( VREG_29_2 ) ;
assign n45700 =  ( n170 ) ? ( n20007 ) : ( n45699 ) ;
assign n45701 =  ( n168 ) ? ( n20006 ) : ( n45700 ) ;
assign n45702 =  ( n166 ) ? ( n20005 ) : ( n45701 ) ;
assign n45703 =  ( n162 ) ? ( n20004 ) : ( n45702 ) ;
assign n45704 =  ( n19987 ) ? ( VREG_29_2 ) : ( n45703 ) ;
assign n45705 =  ( n3051 ) ? ( n45704 ) : ( VREG_29_2 ) ;
assign n45706 =  ( n3040 ) ? ( n45698 ) : ( n45705 ) ;
assign n45707 =  ( n192 ) ? ( VREG_29_2 ) : ( VREG_29_2 ) ;
assign n45708 =  ( n157 ) ? ( n45706 ) : ( n45707 ) ;
assign n45709 =  ( n6 ) ? ( n45693 ) : ( n45708 ) ;
assign n45710 =  ( n659 ) ? ( n45709 ) : ( VREG_29_2 ) ;
assign n45711 =  ( n148 ) ? ( n21065 ) : ( VREG_29_3 ) ;
assign n45712 =  ( n146 ) ? ( n21064 ) : ( n45711 ) ;
assign n45713 =  ( n144 ) ? ( n21063 ) : ( n45712 ) ;
assign n45714 =  ( n142 ) ? ( n21062 ) : ( n45713 ) ;
assign n45715 =  ( n10 ) ? ( n21061 ) : ( n45714 ) ;
assign n45716 =  ( n148 ) ? ( n22099 ) : ( VREG_29_3 ) ;
assign n45717 =  ( n146 ) ? ( n22098 ) : ( n45716 ) ;
assign n45718 =  ( n144 ) ? ( n22097 ) : ( n45717 ) ;
assign n45719 =  ( n142 ) ? ( n22096 ) : ( n45718 ) ;
assign n45720 =  ( n10 ) ? ( n22095 ) : ( n45719 ) ;
assign n45721 =  ( n22106 ) ? ( VREG_29_3 ) : ( n45715 ) ;
assign n45722 =  ( n22106 ) ? ( VREG_29_3 ) : ( n45720 ) ;
assign n45723 =  ( n3034 ) ? ( n45722 ) : ( VREG_29_3 ) ;
assign n45724 =  ( n2965 ) ? ( n45721 ) : ( n45723 ) ;
assign n45725 =  ( n1930 ) ? ( n45720 ) : ( n45724 ) ;
assign n45726 =  ( n879 ) ? ( n45715 ) : ( n45725 ) ;
assign n45727 =  ( n172 ) ? ( n22117 ) : ( VREG_29_3 ) ;
assign n45728 =  ( n170 ) ? ( n22116 ) : ( n45727 ) ;
assign n45729 =  ( n168 ) ? ( n22115 ) : ( n45728 ) ;
assign n45730 =  ( n166 ) ? ( n22114 ) : ( n45729 ) ;
assign n45731 =  ( n162 ) ? ( n22113 ) : ( n45730 ) ;
assign n45732 =  ( n172 ) ? ( n22127 ) : ( VREG_29_3 ) ;
assign n45733 =  ( n170 ) ? ( n22126 ) : ( n45732 ) ;
assign n45734 =  ( n168 ) ? ( n22125 ) : ( n45733 ) ;
assign n45735 =  ( n166 ) ? ( n22124 ) : ( n45734 ) ;
assign n45736 =  ( n162 ) ? ( n22123 ) : ( n45735 ) ;
assign n45737 =  ( n22106 ) ? ( VREG_29_3 ) : ( n45736 ) ;
assign n45738 =  ( n3051 ) ? ( n45737 ) : ( VREG_29_3 ) ;
assign n45739 =  ( n3040 ) ? ( n45731 ) : ( n45738 ) ;
assign n45740 =  ( n192 ) ? ( VREG_29_3 ) : ( VREG_29_3 ) ;
assign n45741 =  ( n157 ) ? ( n45739 ) : ( n45740 ) ;
assign n45742 =  ( n6 ) ? ( n45726 ) : ( n45741 ) ;
assign n45743 =  ( n659 ) ? ( n45742 ) : ( VREG_29_3 ) ;
assign n45744 =  ( n148 ) ? ( n23184 ) : ( VREG_29_4 ) ;
assign n45745 =  ( n146 ) ? ( n23183 ) : ( n45744 ) ;
assign n45746 =  ( n144 ) ? ( n23182 ) : ( n45745 ) ;
assign n45747 =  ( n142 ) ? ( n23181 ) : ( n45746 ) ;
assign n45748 =  ( n10 ) ? ( n23180 ) : ( n45747 ) ;
assign n45749 =  ( n148 ) ? ( n24218 ) : ( VREG_29_4 ) ;
assign n45750 =  ( n146 ) ? ( n24217 ) : ( n45749 ) ;
assign n45751 =  ( n144 ) ? ( n24216 ) : ( n45750 ) ;
assign n45752 =  ( n142 ) ? ( n24215 ) : ( n45751 ) ;
assign n45753 =  ( n10 ) ? ( n24214 ) : ( n45752 ) ;
assign n45754 =  ( n24225 ) ? ( VREG_29_4 ) : ( n45748 ) ;
assign n45755 =  ( n24225 ) ? ( VREG_29_4 ) : ( n45753 ) ;
assign n45756 =  ( n3034 ) ? ( n45755 ) : ( VREG_29_4 ) ;
assign n45757 =  ( n2965 ) ? ( n45754 ) : ( n45756 ) ;
assign n45758 =  ( n1930 ) ? ( n45753 ) : ( n45757 ) ;
assign n45759 =  ( n879 ) ? ( n45748 ) : ( n45758 ) ;
assign n45760 =  ( n172 ) ? ( n24236 ) : ( VREG_29_4 ) ;
assign n45761 =  ( n170 ) ? ( n24235 ) : ( n45760 ) ;
assign n45762 =  ( n168 ) ? ( n24234 ) : ( n45761 ) ;
assign n45763 =  ( n166 ) ? ( n24233 ) : ( n45762 ) ;
assign n45764 =  ( n162 ) ? ( n24232 ) : ( n45763 ) ;
assign n45765 =  ( n172 ) ? ( n24246 ) : ( VREG_29_4 ) ;
assign n45766 =  ( n170 ) ? ( n24245 ) : ( n45765 ) ;
assign n45767 =  ( n168 ) ? ( n24244 ) : ( n45766 ) ;
assign n45768 =  ( n166 ) ? ( n24243 ) : ( n45767 ) ;
assign n45769 =  ( n162 ) ? ( n24242 ) : ( n45768 ) ;
assign n45770 =  ( n24225 ) ? ( VREG_29_4 ) : ( n45769 ) ;
assign n45771 =  ( n3051 ) ? ( n45770 ) : ( VREG_29_4 ) ;
assign n45772 =  ( n3040 ) ? ( n45764 ) : ( n45771 ) ;
assign n45773 =  ( n192 ) ? ( VREG_29_4 ) : ( VREG_29_4 ) ;
assign n45774 =  ( n157 ) ? ( n45772 ) : ( n45773 ) ;
assign n45775 =  ( n6 ) ? ( n45759 ) : ( n45774 ) ;
assign n45776 =  ( n659 ) ? ( n45775 ) : ( VREG_29_4 ) ;
assign n45777 =  ( n148 ) ? ( n25303 ) : ( VREG_29_5 ) ;
assign n45778 =  ( n146 ) ? ( n25302 ) : ( n45777 ) ;
assign n45779 =  ( n144 ) ? ( n25301 ) : ( n45778 ) ;
assign n45780 =  ( n142 ) ? ( n25300 ) : ( n45779 ) ;
assign n45781 =  ( n10 ) ? ( n25299 ) : ( n45780 ) ;
assign n45782 =  ( n148 ) ? ( n26337 ) : ( VREG_29_5 ) ;
assign n45783 =  ( n146 ) ? ( n26336 ) : ( n45782 ) ;
assign n45784 =  ( n144 ) ? ( n26335 ) : ( n45783 ) ;
assign n45785 =  ( n142 ) ? ( n26334 ) : ( n45784 ) ;
assign n45786 =  ( n10 ) ? ( n26333 ) : ( n45785 ) ;
assign n45787 =  ( n26344 ) ? ( VREG_29_5 ) : ( n45781 ) ;
assign n45788 =  ( n26344 ) ? ( VREG_29_5 ) : ( n45786 ) ;
assign n45789 =  ( n3034 ) ? ( n45788 ) : ( VREG_29_5 ) ;
assign n45790 =  ( n2965 ) ? ( n45787 ) : ( n45789 ) ;
assign n45791 =  ( n1930 ) ? ( n45786 ) : ( n45790 ) ;
assign n45792 =  ( n879 ) ? ( n45781 ) : ( n45791 ) ;
assign n45793 =  ( n172 ) ? ( n26355 ) : ( VREG_29_5 ) ;
assign n45794 =  ( n170 ) ? ( n26354 ) : ( n45793 ) ;
assign n45795 =  ( n168 ) ? ( n26353 ) : ( n45794 ) ;
assign n45796 =  ( n166 ) ? ( n26352 ) : ( n45795 ) ;
assign n45797 =  ( n162 ) ? ( n26351 ) : ( n45796 ) ;
assign n45798 =  ( n172 ) ? ( n26365 ) : ( VREG_29_5 ) ;
assign n45799 =  ( n170 ) ? ( n26364 ) : ( n45798 ) ;
assign n45800 =  ( n168 ) ? ( n26363 ) : ( n45799 ) ;
assign n45801 =  ( n166 ) ? ( n26362 ) : ( n45800 ) ;
assign n45802 =  ( n162 ) ? ( n26361 ) : ( n45801 ) ;
assign n45803 =  ( n26344 ) ? ( VREG_29_5 ) : ( n45802 ) ;
assign n45804 =  ( n3051 ) ? ( n45803 ) : ( VREG_29_5 ) ;
assign n45805 =  ( n3040 ) ? ( n45797 ) : ( n45804 ) ;
assign n45806 =  ( n192 ) ? ( VREG_29_5 ) : ( VREG_29_5 ) ;
assign n45807 =  ( n157 ) ? ( n45805 ) : ( n45806 ) ;
assign n45808 =  ( n6 ) ? ( n45792 ) : ( n45807 ) ;
assign n45809 =  ( n659 ) ? ( n45808 ) : ( VREG_29_5 ) ;
assign n45810 =  ( n148 ) ? ( n27422 ) : ( VREG_29_6 ) ;
assign n45811 =  ( n146 ) ? ( n27421 ) : ( n45810 ) ;
assign n45812 =  ( n144 ) ? ( n27420 ) : ( n45811 ) ;
assign n45813 =  ( n142 ) ? ( n27419 ) : ( n45812 ) ;
assign n45814 =  ( n10 ) ? ( n27418 ) : ( n45813 ) ;
assign n45815 =  ( n148 ) ? ( n28456 ) : ( VREG_29_6 ) ;
assign n45816 =  ( n146 ) ? ( n28455 ) : ( n45815 ) ;
assign n45817 =  ( n144 ) ? ( n28454 ) : ( n45816 ) ;
assign n45818 =  ( n142 ) ? ( n28453 ) : ( n45817 ) ;
assign n45819 =  ( n10 ) ? ( n28452 ) : ( n45818 ) ;
assign n45820 =  ( n28463 ) ? ( VREG_29_6 ) : ( n45814 ) ;
assign n45821 =  ( n28463 ) ? ( VREG_29_6 ) : ( n45819 ) ;
assign n45822 =  ( n3034 ) ? ( n45821 ) : ( VREG_29_6 ) ;
assign n45823 =  ( n2965 ) ? ( n45820 ) : ( n45822 ) ;
assign n45824 =  ( n1930 ) ? ( n45819 ) : ( n45823 ) ;
assign n45825 =  ( n879 ) ? ( n45814 ) : ( n45824 ) ;
assign n45826 =  ( n172 ) ? ( n28474 ) : ( VREG_29_6 ) ;
assign n45827 =  ( n170 ) ? ( n28473 ) : ( n45826 ) ;
assign n45828 =  ( n168 ) ? ( n28472 ) : ( n45827 ) ;
assign n45829 =  ( n166 ) ? ( n28471 ) : ( n45828 ) ;
assign n45830 =  ( n162 ) ? ( n28470 ) : ( n45829 ) ;
assign n45831 =  ( n172 ) ? ( n28484 ) : ( VREG_29_6 ) ;
assign n45832 =  ( n170 ) ? ( n28483 ) : ( n45831 ) ;
assign n45833 =  ( n168 ) ? ( n28482 ) : ( n45832 ) ;
assign n45834 =  ( n166 ) ? ( n28481 ) : ( n45833 ) ;
assign n45835 =  ( n162 ) ? ( n28480 ) : ( n45834 ) ;
assign n45836 =  ( n28463 ) ? ( VREG_29_6 ) : ( n45835 ) ;
assign n45837 =  ( n3051 ) ? ( n45836 ) : ( VREG_29_6 ) ;
assign n45838 =  ( n3040 ) ? ( n45830 ) : ( n45837 ) ;
assign n45839 =  ( n192 ) ? ( VREG_29_6 ) : ( VREG_29_6 ) ;
assign n45840 =  ( n157 ) ? ( n45838 ) : ( n45839 ) ;
assign n45841 =  ( n6 ) ? ( n45825 ) : ( n45840 ) ;
assign n45842 =  ( n659 ) ? ( n45841 ) : ( VREG_29_6 ) ;
assign n45843 =  ( n148 ) ? ( n29541 ) : ( VREG_29_7 ) ;
assign n45844 =  ( n146 ) ? ( n29540 ) : ( n45843 ) ;
assign n45845 =  ( n144 ) ? ( n29539 ) : ( n45844 ) ;
assign n45846 =  ( n142 ) ? ( n29538 ) : ( n45845 ) ;
assign n45847 =  ( n10 ) ? ( n29537 ) : ( n45846 ) ;
assign n45848 =  ( n148 ) ? ( n30575 ) : ( VREG_29_7 ) ;
assign n45849 =  ( n146 ) ? ( n30574 ) : ( n45848 ) ;
assign n45850 =  ( n144 ) ? ( n30573 ) : ( n45849 ) ;
assign n45851 =  ( n142 ) ? ( n30572 ) : ( n45850 ) ;
assign n45852 =  ( n10 ) ? ( n30571 ) : ( n45851 ) ;
assign n45853 =  ( n30582 ) ? ( VREG_29_7 ) : ( n45847 ) ;
assign n45854 =  ( n30582 ) ? ( VREG_29_7 ) : ( n45852 ) ;
assign n45855 =  ( n3034 ) ? ( n45854 ) : ( VREG_29_7 ) ;
assign n45856 =  ( n2965 ) ? ( n45853 ) : ( n45855 ) ;
assign n45857 =  ( n1930 ) ? ( n45852 ) : ( n45856 ) ;
assign n45858 =  ( n879 ) ? ( n45847 ) : ( n45857 ) ;
assign n45859 =  ( n172 ) ? ( n30593 ) : ( VREG_29_7 ) ;
assign n45860 =  ( n170 ) ? ( n30592 ) : ( n45859 ) ;
assign n45861 =  ( n168 ) ? ( n30591 ) : ( n45860 ) ;
assign n45862 =  ( n166 ) ? ( n30590 ) : ( n45861 ) ;
assign n45863 =  ( n162 ) ? ( n30589 ) : ( n45862 ) ;
assign n45864 =  ( n172 ) ? ( n30603 ) : ( VREG_29_7 ) ;
assign n45865 =  ( n170 ) ? ( n30602 ) : ( n45864 ) ;
assign n45866 =  ( n168 ) ? ( n30601 ) : ( n45865 ) ;
assign n45867 =  ( n166 ) ? ( n30600 ) : ( n45866 ) ;
assign n45868 =  ( n162 ) ? ( n30599 ) : ( n45867 ) ;
assign n45869 =  ( n30582 ) ? ( VREG_29_7 ) : ( n45868 ) ;
assign n45870 =  ( n3051 ) ? ( n45869 ) : ( VREG_29_7 ) ;
assign n45871 =  ( n3040 ) ? ( n45863 ) : ( n45870 ) ;
assign n45872 =  ( n192 ) ? ( VREG_29_7 ) : ( VREG_29_7 ) ;
assign n45873 =  ( n157 ) ? ( n45871 ) : ( n45872 ) ;
assign n45874 =  ( n6 ) ? ( n45858 ) : ( n45873 ) ;
assign n45875 =  ( n659 ) ? ( n45874 ) : ( VREG_29_7 ) ;
assign n45876 =  ( n148 ) ? ( n31660 ) : ( VREG_29_8 ) ;
assign n45877 =  ( n146 ) ? ( n31659 ) : ( n45876 ) ;
assign n45878 =  ( n144 ) ? ( n31658 ) : ( n45877 ) ;
assign n45879 =  ( n142 ) ? ( n31657 ) : ( n45878 ) ;
assign n45880 =  ( n10 ) ? ( n31656 ) : ( n45879 ) ;
assign n45881 =  ( n148 ) ? ( n32694 ) : ( VREG_29_8 ) ;
assign n45882 =  ( n146 ) ? ( n32693 ) : ( n45881 ) ;
assign n45883 =  ( n144 ) ? ( n32692 ) : ( n45882 ) ;
assign n45884 =  ( n142 ) ? ( n32691 ) : ( n45883 ) ;
assign n45885 =  ( n10 ) ? ( n32690 ) : ( n45884 ) ;
assign n45886 =  ( n32701 ) ? ( VREG_29_8 ) : ( n45880 ) ;
assign n45887 =  ( n32701 ) ? ( VREG_29_8 ) : ( n45885 ) ;
assign n45888 =  ( n3034 ) ? ( n45887 ) : ( VREG_29_8 ) ;
assign n45889 =  ( n2965 ) ? ( n45886 ) : ( n45888 ) ;
assign n45890 =  ( n1930 ) ? ( n45885 ) : ( n45889 ) ;
assign n45891 =  ( n879 ) ? ( n45880 ) : ( n45890 ) ;
assign n45892 =  ( n172 ) ? ( n32712 ) : ( VREG_29_8 ) ;
assign n45893 =  ( n170 ) ? ( n32711 ) : ( n45892 ) ;
assign n45894 =  ( n168 ) ? ( n32710 ) : ( n45893 ) ;
assign n45895 =  ( n166 ) ? ( n32709 ) : ( n45894 ) ;
assign n45896 =  ( n162 ) ? ( n32708 ) : ( n45895 ) ;
assign n45897 =  ( n172 ) ? ( n32722 ) : ( VREG_29_8 ) ;
assign n45898 =  ( n170 ) ? ( n32721 ) : ( n45897 ) ;
assign n45899 =  ( n168 ) ? ( n32720 ) : ( n45898 ) ;
assign n45900 =  ( n166 ) ? ( n32719 ) : ( n45899 ) ;
assign n45901 =  ( n162 ) ? ( n32718 ) : ( n45900 ) ;
assign n45902 =  ( n32701 ) ? ( VREG_29_8 ) : ( n45901 ) ;
assign n45903 =  ( n3051 ) ? ( n45902 ) : ( VREG_29_8 ) ;
assign n45904 =  ( n3040 ) ? ( n45896 ) : ( n45903 ) ;
assign n45905 =  ( n192 ) ? ( VREG_29_8 ) : ( VREG_29_8 ) ;
assign n45906 =  ( n157 ) ? ( n45904 ) : ( n45905 ) ;
assign n45907 =  ( n6 ) ? ( n45891 ) : ( n45906 ) ;
assign n45908 =  ( n659 ) ? ( n45907 ) : ( VREG_29_8 ) ;
assign n45909 =  ( n148 ) ? ( n33779 ) : ( VREG_29_9 ) ;
assign n45910 =  ( n146 ) ? ( n33778 ) : ( n45909 ) ;
assign n45911 =  ( n144 ) ? ( n33777 ) : ( n45910 ) ;
assign n45912 =  ( n142 ) ? ( n33776 ) : ( n45911 ) ;
assign n45913 =  ( n10 ) ? ( n33775 ) : ( n45912 ) ;
assign n45914 =  ( n148 ) ? ( n34813 ) : ( VREG_29_9 ) ;
assign n45915 =  ( n146 ) ? ( n34812 ) : ( n45914 ) ;
assign n45916 =  ( n144 ) ? ( n34811 ) : ( n45915 ) ;
assign n45917 =  ( n142 ) ? ( n34810 ) : ( n45916 ) ;
assign n45918 =  ( n10 ) ? ( n34809 ) : ( n45917 ) ;
assign n45919 =  ( n34820 ) ? ( VREG_29_9 ) : ( n45913 ) ;
assign n45920 =  ( n34820 ) ? ( VREG_29_9 ) : ( n45918 ) ;
assign n45921 =  ( n3034 ) ? ( n45920 ) : ( VREG_29_9 ) ;
assign n45922 =  ( n2965 ) ? ( n45919 ) : ( n45921 ) ;
assign n45923 =  ( n1930 ) ? ( n45918 ) : ( n45922 ) ;
assign n45924 =  ( n879 ) ? ( n45913 ) : ( n45923 ) ;
assign n45925 =  ( n172 ) ? ( n34831 ) : ( VREG_29_9 ) ;
assign n45926 =  ( n170 ) ? ( n34830 ) : ( n45925 ) ;
assign n45927 =  ( n168 ) ? ( n34829 ) : ( n45926 ) ;
assign n45928 =  ( n166 ) ? ( n34828 ) : ( n45927 ) ;
assign n45929 =  ( n162 ) ? ( n34827 ) : ( n45928 ) ;
assign n45930 =  ( n172 ) ? ( n34841 ) : ( VREG_29_9 ) ;
assign n45931 =  ( n170 ) ? ( n34840 ) : ( n45930 ) ;
assign n45932 =  ( n168 ) ? ( n34839 ) : ( n45931 ) ;
assign n45933 =  ( n166 ) ? ( n34838 ) : ( n45932 ) ;
assign n45934 =  ( n162 ) ? ( n34837 ) : ( n45933 ) ;
assign n45935 =  ( n34820 ) ? ( VREG_29_9 ) : ( n45934 ) ;
assign n45936 =  ( n3051 ) ? ( n45935 ) : ( VREG_29_9 ) ;
assign n45937 =  ( n3040 ) ? ( n45929 ) : ( n45936 ) ;
assign n45938 =  ( n192 ) ? ( VREG_29_9 ) : ( VREG_29_9 ) ;
assign n45939 =  ( n157 ) ? ( n45937 ) : ( n45938 ) ;
assign n45940 =  ( n6 ) ? ( n45924 ) : ( n45939 ) ;
assign n45941 =  ( n659 ) ? ( n45940 ) : ( VREG_29_9 ) ;
assign n45942 =  ( n148 ) ? ( n1924 ) : ( VREG_2_0 ) ;
assign n45943 =  ( n146 ) ? ( n1923 ) : ( n45942 ) ;
assign n45944 =  ( n144 ) ? ( n1922 ) : ( n45943 ) ;
assign n45945 =  ( n142 ) ? ( n1921 ) : ( n45944 ) ;
assign n45946 =  ( n10 ) ? ( n1920 ) : ( n45945 ) ;
assign n45947 =  ( n148 ) ? ( n2959 ) : ( VREG_2_0 ) ;
assign n45948 =  ( n146 ) ? ( n2958 ) : ( n45947 ) ;
assign n45949 =  ( n144 ) ? ( n2957 ) : ( n45948 ) ;
assign n45950 =  ( n142 ) ? ( n2956 ) : ( n45949 ) ;
assign n45951 =  ( n10 ) ? ( n2955 ) : ( n45950 ) ;
assign n45952 =  ( n3032 ) ? ( VREG_2_0 ) : ( n45946 ) ;
assign n45953 =  ( n3032 ) ? ( VREG_2_0 ) : ( n45951 ) ;
assign n45954 =  ( n3034 ) ? ( n45953 ) : ( VREG_2_0 ) ;
assign n45955 =  ( n2965 ) ? ( n45952 ) : ( n45954 ) ;
assign n45956 =  ( n1930 ) ? ( n45951 ) : ( n45955 ) ;
assign n45957 =  ( n879 ) ? ( n45946 ) : ( n45956 ) ;
assign n45958 =  ( n172 ) ? ( n3045 ) : ( VREG_2_0 ) ;
assign n45959 =  ( n170 ) ? ( n3044 ) : ( n45958 ) ;
assign n45960 =  ( n168 ) ? ( n3043 ) : ( n45959 ) ;
assign n45961 =  ( n166 ) ? ( n3042 ) : ( n45960 ) ;
assign n45962 =  ( n162 ) ? ( n3041 ) : ( n45961 ) ;
assign n45963 =  ( n172 ) ? ( n3056 ) : ( VREG_2_0 ) ;
assign n45964 =  ( n170 ) ? ( n3055 ) : ( n45963 ) ;
assign n45965 =  ( n168 ) ? ( n3054 ) : ( n45964 ) ;
assign n45966 =  ( n166 ) ? ( n3053 ) : ( n45965 ) ;
assign n45967 =  ( n162 ) ? ( n3052 ) : ( n45966 ) ;
assign n45968 =  ( n3032 ) ? ( VREG_2_0 ) : ( n45967 ) ;
assign n45969 =  ( n3051 ) ? ( n45968 ) : ( VREG_2_0 ) ;
assign n45970 =  ( n3040 ) ? ( n45962 ) : ( n45969 ) ;
assign n45971 =  ( n192 ) ? ( VREG_2_0 ) : ( VREG_2_0 ) ;
assign n45972 =  ( n157 ) ? ( n45970 ) : ( n45971 ) ;
assign n45973 =  ( n6 ) ? ( n45957 ) : ( n45972 ) ;
assign n45974 =  ( n439 ) ? ( n45973 ) : ( VREG_2_0 ) ;
assign n45975 =  ( n148 ) ? ( n4113 ) : ( VREG_2_1 ) ;
assign n45976 =  ( n146 ) ? ( n4112 ) : ( n45975 ) ;
assign n45977 =  ( n144 ) ? ( n4111 ) : ( n45976 ) ;
assign n45978 =  ( n142 ) ? ( n4110 ) : ( n45977 ) ;
assign n45979 =  ( n10 ) ? ( n4109 ) : ( n45978 ) ;
assign n45980 =  ( n148 ) ? ( n5147 ) : ( VREG_2_1 ) ;
assign n45981 =  ( n146 ) ? ( n5146 ) : ( n45980 ) ;
assign n45982 =  ( n144 ) ? ( n5145 ) : ( n45981 ) ;
assign n45983 =  ( n142 ) ? ( n5144 ) : ( n45982 ) ;
assign n45984 =  ( n10 ) ? ( n5143 ) : ( n45983 ) ;
assign n45985 =  ( n5154 ) ? ( VREG_2_1 ) : ( n45979 ) ;
assign n45986 =  ( n5154 ) ? ( VREG_2_1 ) : ( n45984 ) ;
assign n45987 =  ( n3034 ) ? ( n45986 ) : ( VREG_2_1 ) ;
assign n45988 =  ( n2965 ) ? ( n45985 ) : ( n45987 ) ;
assign n45989 =  ( n1930 ) ? ( n45984 ) : ( n45988 ) ;
assign n45990 =  ( n879 ) ? ( n45979 ) : ( n45989 ) ;
assign n45991 =  ( n172 ) ? ( n5165 ) : ( VREG_2_1 ) ;
assign n45992 =  ( n170 ) ? ( n5164 ) : ( n45991 ) ;
assign n45993 =  ( n168 ) ? ( n5163 ) : ( n45992 ) ;
assign n45994 =  ( n166 ) ? ( n5162 ) : ( n45993 ) ;
assign n45995 =  ( n162 ) ? ( n5161 ) : ( n45994 ) ;
assign n45996 =  ( n172 ) ? ( n5175 ) : ( VREG_2_1 ) ;
assign n45997 =  ( n170 ) ? ( n5174 ) : ( n45996 ) ;
assign n45998 =  ( n168 ) ? ( n5173 ) : ( n45997 ) ;
assign n45999 =  ( n166 ) ? ( n5172 ) : ( n45998 ) ;
assign n46000 =  ( n162 ) ? ( n5171 ) : ( n45999 ) ;
assign n46001 =  ( n5154 ) ? ( VREG_2_1 ) : ( n46000 ) ;
assign n46002 =  ( n3051 ) ? ( n46001 ) : ( VREG_2_1 ) ;
assign n46003 =  ( n3040 ) ? ( n45995 ) : ( n46002 ) ;
assign n46004 =  ( n192 ) ? ( VREG_2_1 ) : ( VREG_2_1 ) ;
assign n46005 =  ( n157 ) ? ( n46003 ) : ( n46004 ) ;
assign n46006 =  ( n6 ) ? ( n45990 ) : ( n46005 ) ;
assign n46007 =  ( n439 ) ? ( n46006 ) : ( VREG_2_1 ) ;
assign n46008 =  ( n148 ) ? ( n6232 ) : ( VREG_2_10 ) ;
assign n46009 =  ( n146 ) ? ( n6231 ) : ( n46008 ) ;
assign n46010 =  ( n144 ) ? ( n6230 ) : ( n46009 ) ;
assign n46011 =  ( n142 ) ? ( n6229 ) : ( n46010 ) ;
assign n46012 =  ( n10 ) ? ( n6228 ) : ( n46011 ) ;
assign n46013 =  ( n148 ) ? ( n7266 ) : ( VREG_2_10 ) ;
assign n46014 =  ( n146 ) ? ( n7265 ) : ( n46013 ) ;
assign n46015 =  ( n144 ) ? ( n7264 ) : ( n46014 ) ;
assign n46016 =  ( n142 ) ? ( n7263 ) : ( n46015 ) ;
assign n46017 =  ( n10 ) ? ( n7262 ) : ( n46016 ) ;
assign n46018 =  ( n7273 ) ? ( VREG_2_10 ) : ( n46012 ) ;
assign n46019 =  ( n7273 ) ? ( VREG_2_10 ) : ( n46017 ) ;
assign n46020 =  ( n3034 ) ? ( n46019 ) : ( VREG_2_10 ) ;
assign n46021 =  ( n2965 ) ? ( n46018 ) : ( n46020 ) ;
assign n46022 =  ( n1930 ) ? ( n46017 ) : ( n46021 ) ;
assign n46023 =  ( n879 ) ? ( n46012 ) : ( n46022 ) ;
assign n46024 =  ( n172 ) ? ( n7284 ) : ( VREG_2_10 ) ;
assign n46025 =  ( n170 ) ? ( n7283 ) : ( n46024 ) ;
assign n46026 =  ( n168 ) ? ( n7282 ) : ( n46025 ) ;
assign n46027 =  ( n166 ) ? ( n7281 ) : ( n46026 ) ;
assign n46028 =  ( n162 ) ? ( n7280 ) : ( n46027 ) ;
assign n46029 =  ( n172 ) ? ( n7294 ) : ( VREG_2_10 ) ;
assign n46030 =  ( n170 ) ? ( n7293 ) : ( n46029 ) ;
assign n46031 =  ( n168 ) ? ( n7292 ) : ( n46030 ) ;
assign n46032 =  ( n166 ) ? ( n7291 ) : ( n46031 ) ;
assign n46033 =  ( n162 ) ? ( n7290 ) : ( n46032 ) ;
assign n46034 =  ( n7273 ) ? ( VREG_2_10 ) : ( n46033 ) ;
assign n46035 =  ( n3051 ) ? ( n46034 ) : ( VREG_2_10 ) ;
assign n46036 =  ( n3040 ) ? ( n46028 ) : ( n46035 ) ;
assign n46037 =  ( n192 ) ? ( VREG_2_10 ) : ( VREG_2_10 ) ;
assign n46038 =  ( n157 ) ? ( n46036 ) : ( n46037 ) ;
assign n46039 =  ( n6 ) ? ( n46023 ) : ( n46038 ) ;
assign n46040 =  ( n439 ) ? ( n46039 ) : ( VREG_2_10 ) ;
assign n46041 =  ( n148 ) ? ( n8351 ) : ( VREG_2_11 ) ;
assign n46042 =  ( n146 ) ? ( n8350 ) : ( n46041 ) ;
assign n46043 =  ( n144 ) ? ( n8349 ) : ( n46042 ) ;
assign n46044 =  ( n142 ) ? ( n8348 ) : ( n46043 ) ;
assign n46045 =  ( n10 ) ? ( n8347 ) : ( n46044 ) ;
assign n46046 =  ( n148 ) ? ( n9385 ) : ( VREG_2_11 ) ;
assign n46047 =  ( n146 ) ? ( n9384 ) : ( n46046 ) ;
assign n46048 =  ( n144 ) ? ( n9383 ) : ( n46047 ) ;
assign n46049 =  ( n142 ) ? ( n9382 ) : ( n46048 ) ;
assign n46050 =  ( n10 ) ? ( n9381 ) : ( n46049 ) ;
assign n46051 =  ( n9392 ) ? ( VREG_2_11 ) : ( n46045 ) ;
assign n46052 =  ( n9392 ) ? ( VREG_2_11 ) : ( n46050 ) ;
assign n46053 =  ( n3034 ) ? ( n46052 ) : ( VREG_2_11 ) ;
assign n46054 =  ( n2965 ) ? ( n46051 ) : ( n46053 ) ;
assign n46055 =  ( n1930 ) ? ( n46050 ) : ( n46054 ) ;
assign n46056 =  ( n879 ) ? ( n46045 ) : ( n46055 ) ;
assign n46057 =  ( n172 ) ? ( n9403 ) : ( VREG_2_11 ) ;
assign n46058 =  ( n170 ) ? ( n9402 ) : ( n46057 ) ;
assign n46059 =  ( n168 ) ? ( n9401 ) : ( n46058 ) ;
assign n46060 =  ( n166 ) ? ( n9400 ) : ( n46059 ) ;
assign n46061 =  ( n162 ) ? ( n9399 ) : ( n46060 ) ;
assign n46062 =  ( n172 ) ? ( n9413 ) : ( VREG_2_11 ) ;
assign n46063 =  ( n170 ) ? ( n9412 ) : ( n46062 ) ;
assign n46064 =  ( n168 ) ? ( n9411 ) : ( n46063 ) ;
assign n46065 =  ( n166 ) ? ( n9410 ) : ( n46064 ) ;
assign n46066 =  ( n162 ) ? ( n9409 ) : ( n46065 ) ;
assign n46067 =  ( n9392 ) ? ( VREG_2_11 ) : ( n46066 ) ;
assign n46068 =  ( n3051 ) ? ( n46067 ) : ( VREG_2_11 ) ;
assign n46069 =  ( n3040 ) ? ( n46061 ) : ( n46068 ) ;
assign n46070 =  ( n192 ) ? ( VREG_2_11 ) : ( VREG_2_11 ) ;
assign n46071 =  ( n157 ) ? ( n46069 ) : ( n46070 ) ;
assign n46072 =  ( n6 ) ? ( n46056 ) : ( n46071 ) ;
assign n46073 =  ( n439 ) ? ( n46072 ) : ( VREG_2_11 ) ;
assign n46074 =  ( n148 ) ? ( n10470 ) : ( VREG_2_12 ) ;
assign n46075 =  ( n146 ) ? ( n10469 ) : ( n46074 ) ;
assign n46076 =  ( n144 ) ? ( n10468 ) : ( n46075 ) ;
assign n46077 =  ( n142 ) ? ( n10467 ) : ( n46076 ) ;
assign n46078 =  ( n10 ) ? ( n10466 ) : ( n46077 ) ;
assign n46079 =  ( n148 ) ? ( n11504 ) : ( VREG_2_12 ) ;
assign n46080 =  ( n146 ) ? ( n11503 ) : ( n46079 ) ;
assign n46081 =  ( n144 ) ? ( n11502 ) : ( n46080 ) ;
assign n46082 =  ( n142 ) ? ( n11501 ) : ( n46081 ) ;
assign n46083 =  ( n10 ) ? ( n11500 ) : ( n46082 ) ;
assign n46084 =  ( n11511 ) ? ( VREG_2_12 ) : ( n46078 ) ;
assign n46085 =  ( n11511 ) ? ( VREG_2_12 ) : ( n46083 ) ;
assign n46086 =  ( n3034 ) ? ( n46085 ) : ( VREG_2_12 ) ;
assign n46087 =  ( n2965 ) ? ( n46084 ) : ( n46086 ) ;
assign n46088 =  ( n1930 ) ? ( n46083 ) : ( n46087 ) ;
assign n46089 =  ( n879 ) ? ( n46078 ) : ( n46088 ) ;
assign n46090 =  ( n172 ) ? ( n11522 ) : ( VREG_2_12 ) ;
assign n46091 =  ( n170 ) ? ( n11521 ) : ( n46090 ) ;
assign n46092 =  ( n168 ) ? ( n11520 ) : ( n46091 ) ;
assign n46093 =  ( n166 ) ? ( n11519 ) : ( n46092 ) ;
assign n46094 =  ( n162 ) ? ( n11518 ) : ( n46093 ) ;
assign n46095 =  ( n172 ) ? ( n11532 ) : ( VREG_2_12 ) ;
assign n46096 =  ( n170 ) ? ( n11531 ) : ( n46095 ) ;
assign n46097 =  ( n168 ) ? ( n11530 ) : ( n46096 ) ;
assign n46098 =  ( n166 ) ? ( n11529 ) : ( n46097 ) ;
assign n46099 =  ( n162 ) ? ( n11528 ) : ( n46098 ) ;
assign n46100 =  ( n11511 ) ? ( VREG_2_12 ) : ( n46099 ) ;
assign n46101 =  ( n3051 ) ? ( n46100 ) : ( VREG_2_12 ) ;
assign n46102 =  ( n3040 ) ? ( n46094 ) : ( n46101 ) ;
assign n46103 =  ( n192 ) ? ( VREG_2_12 ) : ( VREG_2_12 ) ;
assign n46104 =  ( n157 ) ? ( n46102 ) : ( n46103 ) ;
assign n46105 =  ( n6 ) ? ( n46089 ) : ( n46104 ) ;
assign n46106 =  ( n439 ) ? ( n46105 ) : ( VREG_2_12 ) ;
assign n46107 =  ( n148 ) ? ( n12589 ) : ( VREG_2_13 ) ;
assign n46108 =  ( n146 ) ? ( n12588 ) : ( n46107 ) ;
assign n46109 =  ( n144 ) ? ( n12587 ) : ( n46108 ) ;
assign n46110 =  ( n142 ) ? ( n12586 ) : ( n46109 ) ;
assign n46111 =  ( n10 ) ? ( n12585 ) : ( n46110 ) ;
assign n46112 =  ( n148 ) ? ( n13623 ) : ( VREG_2_13 ) ;
assign n46113 =  ( n146 ) ? ( n13622 ) : ( n46112 ) ;
assign n46114 =  ( n144 ) ? ( n13621 ) : ( n46113 ) ;
assign n46115 =  ( n142 ) ? ( n13620 ) : ( n46114 ) ;
assign n46116 =  ( n10 ) ? ( n13619 ) : ( n46115 ) ;
assign n46117 =  ( n13630 ) ? ( VREG_2_13 ) : ( n46111 ) ;
assign n46118 =  ( n13630 ) ? ( VREG_2_13 ) : ( n46116 ) ;
assign n46119 =  ( n3034 ) ? ( n46118 ) : ( VREG_2_13 ) ;
assign n46120 =  ( n2965 ) ? ( n46117 ) : ( n46119 ) ;
assign n46121 =  ( n1930 ) ? ( n46116 ) : ( n46120 ) ;
assign n46122 =  ( n879 ) ? ( n46111 ) : ( n46121 ) ;
assign n46123 =  ( n172 ) ? ( n13641 ) : ( VREG_2_13 ) ;
assign n46124 =  ( n170 ) ? ( n13640 ) : ( n46123 ) ;
assign n46125 =  ( n168 ) ? ( n13639 ) : ( n46124 ) ;
assign n46126 =  ( n166 ) ? ( n13638 ) : ( n46125 ) ;
assign n46127 =  ( n162 ) ? ( n13637 ) : ( n46126 ) ;
assign n46128 =  ( n172 ) ? ( n13651 ) : ( VREG_2_13 ) ;
assign n46129 =  ( n170 ) ? ( n13650 ) : ( n46128 ) ;
assign n46130 =  ( n168 ) ? ( n13649 ) : ( n46129 ) ;
assign n46131 =  ( n166 ) ? ( n13648 ) : ( n46130 ) ;
assign n46132 =  ( n162 ) ? ( n13647 ) : ( n46131 ) ;
assign n46133 =  ( n13630 ) ? ( VREG_2_13 ) : ( n46132 ) ;
assign n46134 =  ( n3051 ) ? ( n46133 ) : ( VREG_2_13 ) ;
assign n46135 =  ( n3040 ) ? ( n46127 ) : ( n46134 ) ;
assign n46136 =  ( n192 ) ? ( VREG_2_13 ) : ( VREG_2_13 ) ;
assign n46137 =  ( n157 ) ? ( n46135 ) : ( n46136 ) ;
assign n46138 =  ( n6 ) ? ( n46122 ) : ( n46137 ) ;
assign n46139 =  ( n439 ) ? ( n46138 ) : ( VREG_2_13 ) ;
assign n46140 =  ( n148 ) ? ( n14708 ) : ( VREG_2_14 ) ;
assign n46141 =  ( n146 ) ? ( n14707 ) : ( n46140 ) ;
assign n46142 =  ( n144 ) ? ( n14706 ) : ( n46141 ) ;
assign n46143 =  ( n142 ) ? ( n14705 ) : ( n46142 ) ;
assign n46144 =  ( n10 ) ? ( n14704 ) : ( n46143 ) ;
assign n46145 =  ( n148 ) ? ( n15742 ) : ( VREG_2_14 ) ;
assign n46146 =  ( n146 ) ? ( n15741 ) : ( n46145 ) ;
assign n46147 =  ( n144 ) ? ( n15740 ) : ( n46146 ) ;
assign n46148 =  ( n142 ) ? ( n15739 ) : ( n46147 ) ;
assign n46149 =  ( n10 ) ? ( n15738 ) : ( n46148 ) ;
assign n46150 =  ( n15749 ) ? ( VREG_2_14 ) : ( n46144 ) ;
assign n46151 =  ( n15749 ) ? ( VREG_2_14 ) : ( n46149 ) ;
assign n46152 =  ( n3034 ) ? ( n46151 ) : ( VREG_2_14 ) ;
assign n46153 =  ( n2965 ) ? ( n46150 ) : ( n46152 ) ;
assign n46154 =  ( n1930 ) ? ( n46149 ) : ( n46153 ) ;
assign n46155 =  ( n879 ) ? ( n46144 ) : ( n46154 ) ;
assign n46156 =  ( n172 ) ? ( n15760 ) : ( VREG_2_14 ) ;
assign n46157 =  ( n170 ) ? ( n15759 ) : ( n46156 ) ;
assign n46158 =  ( n168 ) ? ( n15758 ) : ( n46157 ) ;
assign n46159 =  ( n166 ) ? ( n15757 ) : ( n46158 ) ;
assign n46160 =  ( n162 ) ? ( n15756 ) : ( n46159 ) ;
assign n46161 =  ( n172 ) ? ( n15770 ) : ( VREG_2_14 ) ;
assign n46162 =  ( n170 ) ? ( n15769 ) : ( n46161 ) ;
assign n46163 =  ( n168 ) ? ( n15768 ) : ( n46162 ) ;
assign n46164 =  ( n166 ) ? ( n15767 ) : ( n46163 ) ;
assign n46165 =  ( n162 ) ? ( n15766 ) : ( n46164 ) ;
assign n46166 =  ( n15749 ) ? ( VREG_2_14 ) : ( n46165 ) ;
assign n46167 =  ( n3051 ) ? ( n46166 ) : ( VREG_2_14 ) ;
assign n46168 =  ( n3040 ) ? ( n46160 ) : ( n46167 ) ;
assign n46169 =  ( n192 ) ? ( VREG_2_14 ) : ( VREG_2_14 ) ;
assign n46170 =  ( n157 ) ? ( n46168 ) : ( n46169 ) ;
assign n46171 =  ( n6 ) ? ( n46155 ) : ( n46170 ) ;
assign n46172 =  ( n439 ) ? ( n46171 ) : ( VREG_2_14 ) ;
assign n46173 =  ( n148 ) ? ( n16827 ) : ( VREG_2_15 ) ;
assign n46174 =  ( n146 ) ? ( n16826 ) : ( n46173 ) ;
assign n46175 =  ( n144 ) ? ( n16825 ) : ( n46174 ) ;
assign n46176 =  ( n142 ) ? ( n16824 ) : ( n46175 ) ;
assign n46177 =  ( n10 ) ? ( n16823 ) : ( n46176 ) ;
assign n46178 =  ( n148 ) ? ( n17861 ) : ( VREG_2_15 ) ;
assign n46179 =  ( n146 ) ? ( n17860 ) : ( n46178 ) ;
assign n46180 =  ( n144 ) ? ( n17859 ) : ( n46179 ) ;
assign n46181 =  ( n142 ) ? ( n17858 ) : ( n46180 ) ;
assign n46182 =  ( n10 ) ? ( n17857 ) : ( n46181 ) ;
assign n46183 =  ( n17868 ) ? ( VREG_2_15 ) : ( n46177 ) ;
assign n46184 =  ( n17868 ) ? ( VREG_2_15 ) : ( n46182 ) ;
assign n46185 =  ( n3034 ) ? ( n46184 ) : ( VREG_2_15 ) ;
assign n46186 =  ( n2965 ) ? ( n46183 ) : ( n46185 ) ;
assign n46187 =  ( n1930 ) ? ( n46182 ) : ( n46186 ) ;
assign n46188 =  ( n879 ) ? ( n46177 ) : ( n46187 ) ;
assign n46189 =  ( n172 ) ? ( n17879 ) : ( VREG_2_15 ) ;
assign n46190 =  ( n170 ) ? ( n17878 ) : ( n46189 ) ;
assign n46191 =  ( n168 ) ? ( n17877 ) : ( n46190 ) ;
assign n46192 =  ( n166 ) ? ( n17876 ) : ( n46191 ) ;
assign n46193 =  ( n162 ) ? ( n17875 ) : ( n46192 ) ;
assign n46194 =  ( n172 ) ? ( n17889 ) : ( VREG_2_15 ) ;
assign n46195 =  ( n170 ) ? ( n17888 ) : ( n46194 ) ;
assign n46196 =  ( n168 ) ? ( n17887 ) : ( n46195 ) ;
assign n46197 =  ( n166 ) ? ( n17886 ) : ( n46196 ) ;
assign n46198 =  ( n162 ) ? ( n17885 ) : ( n46197 ) ;
assign n46199 =  ( n17868 ) ? ( VREG_2_15 ) : ( n46198 ) ;
assign n46200 =  ( n3051 ) ? ( n46199 ) : ( VREG_2_15 ) ;
assign n46201 =  ( n3040 ) ? ( n46193 ) : ( n46200 ) ;
assign n46202 =  ( n192 ) ? ( VREG_2_15 ) : ( VREG_2_15 ) ;
assign n46203 =  ( n157 ) ? ( n46201 ) : ( n46202 ) ;
assign n46204 =  ( n6 ) ? ( n46188 ) : ( n46203 ) ;
assign n46205 =  ( n439 ) ? ( n46204 ) : ( VREG_2_15 ) ;
assign n46206 =  ( n148 ) ? ( n18946 ) : ( VREG_2_2 ) ;
assign n46207 =  ( n146 ) ? ( n18945 ) : ( n46206 ) ;
assign n46208 =  ( n144 ) ? ( n18944 ) : ( n46207 ) ;
assign n46209 =  ( n142 ) ? ( n18943 ) : ( n46208 ) ;
assign n46210 =  ( n10 ) ? ( n18942 ) : ( n46209 ) ;
assign n46211 =  ( n148 ) ? ( n19980 ) : ( VREG_2_2 ) ;
assign n46212 =  ( n146 ) ? ( n19979 ) : ( n46211 ) ;
assign n46213 =  ( n144 ) ? ( n19978 ) : ( n46212 ) ;
assign n46214 =  ( n142 ) ? ( n19977 ) : ( n46213 ) ;
assign n46215 =  ( n10 ) ? ( n19976 ) : ( n46214 ) ;
assign n46216 =  ( n19987 ) ? ( VREG_2_2 ) : ( n46210 ) ;
assign n46217 =  ( n19987 ) ? ( VREG_2_2 ) : ( n46215 ) ;
assign n46218 =  ( n3034 ) ? ( n46217 ) : ( VREG_2_2 ) ;
assign n46219 =  ( n2965 ) ? ( n46216 ) : ( n46218 ) ;
assign n46220 =  ( n1930 ) ? ( n46215 ) : ( n46219 ) ;
assign n46221 =  ( n879 ) ? ( n46210 ) : ( n46220 ) ;
assign n46222 =  ( n172 ) ? ( n19998 ) : ( VREG_2_2 ) ;
assign n46223 =  ( n170 ) ? ( n19997 ) : ( n46222 ) ;
assign n46224 =  ( n168 ) ? ( n19996 ) : ( n46223 ) ;
assign n46225 =  ( n166 ) ? ( n19995 ) : ( n46224 ) ;
assign n46226 =  ( n162 ) ? ( n19994 ) : ( n46225 ) ;
assign n46227 =  ( n172 ) ? ( n20008 ) : ( VREG_2_2 ) ;
assign n46228 =  ( n170 ) ? ( n20007 ) : ( n46227 ) ;
assign n46229 =  ( n168 ) ? ( n20006 ) : ( n46228 ) ;
assign n46230 =  ( n166 ) ? ( n20005 ) : ( n46229 ) ;
assign n46231 =  ( n162 ) ? ( n20004 ) : ( n46230 ) ;
assign n46232 =  ( n19987 ) ? ( VREG_2_2 ) : ( n46231 ) ;
assign n46233 =  ( n3051 ) ? ( n46232 ) : ( VREG_2_2 ) ;
assign n46234 =  ( n3040 ) ? ( n46226 ) : ( n46233 ) ;
assign n46235 =  ( n192 ) ? ( VREG_2_2 ) : ( VREG_2_2 ) ;
assign n46236 =  ( n157 ) ? ( n46234 ) : ( n46235 ) ;
assign n46237 =  ( n6 ) ? ( n46221 ) : ( n46236 ) ;
assign n46238 =  ( n439 ) ? ( n46237 ) : ( VREG_2_2 ) ;
assign n46239 =  ( n148 ) ? ( n21065 ) : ( VREG_2_3 ) ;
assign n46240 =  ( n146 ) ? ( n21064 ) : ( n46239 ) ;
assign n46241 =  ( n144 ) ? ( n21063 ) : ( n46240 ) ;
assign n46242 =  ( n142 ) ? ( n21062 ) : ( n46241 ) ;
assign n46243 =  ( n10 ) ? ( n21061 ) : ( n46242 ) ;
assign n46244 =  ( n148 ) ? ( n22099 ) : ( VREG_2_3 ) ;
assign n46245 =  ( n146 ) ? ( n22098 ) : ( n46244 ) ;
assign n46246 =  ( n144 ) ? ( n22097 ) : ( n46245 ) ;
assign n46247 =  ( n142 ) ? ( n22096 ) : ( n46246 ) ;
assign n46248 =  ( n10 ) ? ( n22095 ) : ( n46247 ) ;
assign n46249 =  ( n22106 ) ? ( VREG_2_3 ) : ( n46243 ) ;
assign n46250 =  ( n22106 ) ? ( VREG_2_3 ) : ( n46248 ) ;
assign n46251 =  ( n3034 ) ? ( n46250 ) : ( VREG_2_3 ) ;
assign n46252 =  ( n2965 ) ? ( n46249 ) : ( n46251 ) ;
assign n46253 =  ( n1930 ) ? ( n46248 ) : ( n46252 ) ;
assign n46254 =  ( n879 ) ? ( n46243 ) : ( n46253 ) ;
assign n46255 =  ( n172 ) ? ( n22117 ) : ( VREG_2_3 ) ;
assign n46256 =  ( n170 ) ? ( n22116 ) : ( n46255 ) ;
assign n46257 =  ( n168 ) ? ( n22115 ) : ( n46256 ) ;
assign n46258 =  ( n166 ) ? ( n22114 ) : ( n46257 ) ;
assign n46259 =  ( n162 ) ? ( n22113 ) : ( n46258 ) ;
assign n46260 =  ( n172 ) ? ( n22127 ) : ( VREG_2_3 ) ;
assign n46261 =  ( n170 ) ? ( n22126 ) : ( n46260 ) ;
assign n46262 =  ( n168 ) ? ( n22125 ) : ( n46261 ) ;
assign n46263 =  ( n166 ) ? ( n22124 ) : ( n46262 ) ;
assign n46264 =  ( n162 ) ? ( n22123 ) : ( n46263 ) ;
assign n46265 =  ( n22106 ) ? ( VREG_2_3 ) : ( n46264 ) ;
assign n46266 =  ( n3051 ) ? ( n46265 ) : ( VREG_2_3 ) ;
assign n46267 =  ( n3040 ) ? ( n46259 ) : ( n46266 ) ;
assign n46268 =  ( n192 ) ? ( VREG_2_3 ) : ( VREG_2_3 ) ;
assign n46269 =  ( n157 ) ? ( n46267 ) : ( n46268 ) ;
assign n46270 =  ( n6 ) ? ( n46254 ) : ( n46269 ) ;
assign n46271 =  ( n439 ) ? ( n46270 ) : ( VREG_2_3 ) ;
assign n46272 =  ( n148 ) ? ( n23184 ) : ( VREG_2_4 ) ;
assign n46273 =  ( n146 ) ? ( n23183 ) : ( n46272 ) ;
assign n46274 =  ( n144 ) ? ( n23182 ) : ( n46273 ) ;
assign n46275 =  ( n142 ) ? ( n23181 ) : ( n46274 ) ;
assign n46276 =  ( n10 ) ? ( n23180 ) : ( n46275 ) ;
assign n46277 =  ( n148 ) ? ( n24218 ) : ( VREG_2_4 ) ;
assign n46278 =  ( n146 ) ? ( n24217 ) : ( n46277 ) ;
assign n46279 =  ( n144 ) ? ( n24216 ) : ( n46278 ) ;
assign n46280 =  ( n142 ) ? ( n24215 ) : ( n46279 ) ;
assign n46281 =  ( n10 ) ? ( n24214 ) : ( n46280 ) ;
assign n46282 =  ( n24225 ) ? ( VREG_2_4 ) : ( n46276 ) ;
assign n46283 =  ( n24225 ) ? ( VREG_2_4 ) : ( n46281 ) ;
assign n46284 =  ( n3034 ) ? ( n46283 ) : ( VREG_2_4 ) ;
assign n46285 =  ( n2965 ) ? ( n46282 ) : ( n46284 ) ;
assign n46286 =  ( n1930 ) ? ( n46281 ) : ( n46285 ) ;
assign n46287 =  ( n879 ) ? ( n46276 ) : ( n46286 ) ;
assign n46288 =  ( n172 ) ? ( n24236 ) : ( VREG_2_4 ) ;
assign n46289 =  ( n170 ) ? ( n24235 ) : ( n46288 ) ;
assign n46290 =  ( n168 ) ? ( n24234 ) : ( n46289 ) ;
assign n46291 =  ( n166 ) ? ( n24233 ) : ( n46290 ) ;
assign n46292 =  ( n162 ) ? ( n24232 ) : ( n46291 ) ;
assign n46293 =  ( n172 ) ? ( n24246 ) : ( VREG_2_4 ) ;
assign n46294 =  ( n170 ) ? ( n24245 ) : ( n46293 ) ;
assign n46295 =  ( n168 ) ? ( n24244 ) : ( n46294 ) ;
assign n46296 =  ( n166 ) ? ( n24243 ) : ( n46295 ) ;
assign n46297 =  ( n162 ) ? ( n24242 ) : ( n46296 ) ;
assign n46298 =  ( n24225 ) ? ( VREG_2_4 ) : ( n46297 ) ;
assign n46299 =  ( n3051 ) ? ( n46298 ) : ( VREG_2_4 ) ;
assign n46300 =  ( n3040 ) ? ( n46292 ) : ( n46299 ) ;
assign n46301 =  ( n192 ) ? ( VREG_2_4 ) : ( VREG_2_4 ) ;
assign n46302 =  ( n157 ) ? ( n46300 ) : ( n46301 ) ;
assign n46303 =  ( n6 ) ? ( n46287 ) : ( n46302 ) ;
assign n46304 =  ( n439 ) ? ( n46303 ) : ( VREG_2_4 ) ;
assign n46305 =  ( n148 ) ? ( n25303 ) : ( VREG_2_5 ) ;
assign n46306 =  ( n146 ) ? ( n25302 ) : ( n46305 ) ;
assign n46307 =  ( n144 ) ? ( n25301 ) : ( n46306 ) ;
assign n46308 =  ( n142 ) ? ( n25300 ) : ( n46307 ) ;
assign n46309 =  ( n10 ) ? ( n25299 ) : ( n46308 ) ;
assign n46310 =  ( n148 ) ? ( n26337 ) : ( VREG_2_5 ) ;
assign n46311 =  ( n146 ) ? ( n26336 ) : ( n46310 ) ;
assign n46312 =  ( n144 ) ? ( n26335 ) : ( n46311 ) ;
assign n46313 =  ( n142 ) ? ( n26334 ) : ( n46312 ) ;
assign n46314 =  ( n10 ) ? ( n26333 ) : ( n46313 ) ;
assign n46315 =  ( n26344 ) ? ( VREG_2_5 ) : ( n46309 ) ;
assign n46316 =  ( n26344 ) ? ( VREG_2_5 ) : ( n46314 ) ;
assign n46317 =  ( n3034 ) ? ( n46316 ) : ( VREG_2_5 ) ;
assign n46318 =  ( n2965 ) ? ( n46315 ) : ( n46317 ) ;
assign n46319 =  ( n1930 ) ? ( n46314 ) : ( n46318 ) ;
assign n46320 =  ( n879 ) ? ( n46309 ) : ( n46319 ) ;
assign n46321 =  ( n172 ) ? ( n26355 ) : ( VREG_2_5 ) ;
assign n46322 =  ( n170 ) ? ( n26354 ) : ( n46321 ) ;
assign n46323 =  ( n168 ) ? ( n26353 ) : ( n46322 ) ;
assign n46324 =  ( n166 ) ? ( n26352 ) : ( n46323 ) ;
assign n46325 =  ( n162 ) ? ( n26351 ) : ( n46324 ) ;
assign n46326 =  ( n172 ) ? ( n26365 ) : ( VREG_2_5 ) ;
assign n46327 =  ( n170 ) ? ( n26364 ) : ( n46326 ) ;
assign n46328 =  ( n168 ) ? ( n26363 ) : ( n46327 ) ;
assign n46329 =  ( n166 ) ? ( n26362 ) : ( n46328 ) ;
assign n46330 =  ( n162 ) ? ( n26361 ) : ( n46329 ) ;
assign n46331 =  ( n26344 ) ? ( VREG_2_5 ) : ( n46330 ) ;
assign n46332 =  ( n3051 ) ? ( n46331 ) : ( VREG_2_5 ) ;
assign n46333 =  ( n3040 ) ? ( n46325 ) : ( n46332 ) ;
assign n46334 =  ( n192 ) ? ( VREG_2_5 ) : ( VREG_2_5 ) ;
assign n46335 =  ( n157 ) ? ( n46333 ) : ( n46334 ) ;
assign n46336 =  ( n6 ) ? ( n46320 ) : ( n46335 ) ;
assign n46337 =  ( n439 ) ? ( n46336 ) : ( VREG_2_5 ) ;
assign n46338 =  ( n148 ) ? ( n27422 ) : ( VREG_2_6 ) ;
assign n46339 =  ( n146 ) ? ( n27421 ) : ( n46338 ) ;
assign n46340 =  ( n144 ) ? ( n27420 ) : ( n46339 ) ;
assign n46341 =  ( n142 ) ? ( n27419 ) : ( n46340 ) ;
assign n46342 =  ( n10 ) ? ( n27418 ) : ( n46341 ) ;
assign n46343 =  ( n148 ) ? ( n28456 ) : ( VREG_2_6 ) ;
assign n46344 =  ( n146 ) ? ( n28455 ) : ( n46343 ) ;
assign n46345 =  ( n144 ) ? ( n28454 ) : ( n46344 ) ;
assign n46346 =  ( n142 ) ? ( n28453 ) : ( n46345 ) ;
assign n46347 =  ( n10 ) ? ( n28452 ) : ( n46346 ) ;
assign n46348 =  ( n28463 ) ? ( VREG_2_6 ) : ( n46342 ) ;
assign n46349 =  ( n28463 ) ? ( VREG_2_6 ) : ( n46347 ) ;
assign n46350 =  ( n3034 ) ? ( n46349 ) : ( VREG_2_6 ) ;
assign n46351 =  ( n2965 ) ? ( n46348 ) : ( n46350 ) ;
assign n46352 =  ( n1930 ) ? ( n46347 ) : ( n46351 ) ;
assign n46353 =  ( n879 ) ? ( n46342 ) : ( n46352 ) ;
assign n46354 =  ( n172 ) ? ( n28474 ) : ( VREG_2_6 ) ;
assign n46355 =  ( n170 ) ? ( n28473 ) : ( n46354 ) ;
assign n46356 =  ( n168 ) ? ( n28472 ) : ( n46355 ) ;
assign n46357 =  ( n166 ) ? ( n28471 ) : ( n46356 ) ;
assign n46358 =  ( n162 ) ? ( n28470 ) : ( n46357 ) ;
assign n46359 =  ( n172 ) ? ( n28484 ) : ( VREG_2_6 ) ;
assign n46360 =  ( n170 ) ? ( n28483 ) : ( n46359 ) ;
assign n46361 =  ( n168 ) ? ( n28482 ) : ( n46360 ) ;
assign n46362 =  ( n166 ) ? ( n28481 ) : ( n46361 ) ;
assign n46363 =  ( n162 ) ? ( n28480 ) : ( n46362 ) ;
assign n46364 =  ( n28463 ) ? ( VREG_2_6 ) : ( n46363 ) ;
assign n46365 =  ( n3051 ) ? ( n46364 ) : ( VREG_2_6 ) ;
assign n46366 =  ( n3040 ) ? ( n46358 ) : ( n46365 ) ;
assign n46367 =  ( n192 ) ? ( VREG_2_6 ) : ( VREG_2_6 ) ;
assign n46368 =  ( n157 ) ? ( n46366 ) : ( n46367 ) ;
assign n46369 =  ( n6 ) ? ( n46353 ) : ( n46368 ) ;
assign n46370 =  ( n439 ) ? ( n46369 ) : ( VREG_2_6 ) ;
assign n46371 =  ( n148 ) ? ( n29541 ) : ( VREG_2_7 ) ;
assign n46372 =  ( n146 ) ? ( n29540 ) : ( n46371 ) ;
assign n46373 =  ( n144 ) ? ( n29539 ) : ( n46372 ) ;
assign n46374 =  ( n142 ) ? ( n29538 ) : ( n46373 ) ;
assign n46375 =  ( n10 ) ? ( n29537 ) : ( n46374 ) ;
assign n46376 =  ( n148 ) ? ( n30575 ) : ( VREG_2_7 ) ;
assign n46377 =  ( n146 ) ? ( n30574 ) : ( n46376 ) ;
assign n46378 =  ( n144 ) ? ( n30573 ) : ( n46377 ) ;
assign n46379 =  ( n142 ) ? ( n30572 ) : ( n46378 ) ;
assign n46380 =  ( n10 ) ? ( n30571 ) : ( n46379 ) ;
assign n46381 =  ( n30582 ) ? ( VREG_2_7 ) : ( n46375 ) ;
assign n46382 =  ( n30582 ) ? ( VREG_2_7 ) : ( n46380 ) ;
assign n46383 =  ( n3034 ) ? ( n46382 ) : ( VREG_2_7 ) ;
assign n46384 =  ( n2965 ) ? ( n46381 ) : ( n46383 ) ;
assign n46385 =  ( n1930 ) ? ( n46380 ) : ( n46384 ) ;
assign n46386 =  ( n879 ) ? ( n46375 ) : ( n46385 ) ;
assign n46387 =  ( n172 ) ? ( n30593 ) : ( VREG_2_7 ) ;
assign n46388 =  ( n170 ) ? ( n30592 ) : ( n46387 ) ;
assign n46389 =  ( n168 ) ? ( n30591 ) : ( n46388 ) ;
assign n46390 =  ( n166 ) ? ( n30590 ) : ( n46389 ) ;
assign n46391 =  ( n162 ) ? ( n30589 ) : ( n46390 ) ;
assign n46392 =  ( n172 ) ? ( n30603 ) : ( VREG_2_7 ) ;
assign n46393 =  ( n170 ) ? ( n30602 ) : ( n46392 ) ;
assign n46394 =  ( n168 ) ? ( n30601 ) : ( n46393 ) ;
assign n46395 =  ( n166 ) ? ( n30600 ) : ( n46394 ) ;
assign n46396 =  ( n162 ) ? ( n30599 ) : ( n46395 ) ;
assign n46397 =  ( n30582 ) ? ( VREG_2_7 ) : ( n46396 ) ;
assign n46398 =  ( n3051 ) ? ( n46397 ) : ( VREG_2_7 ) ;
assign n46399 =  ( n3040 ) ? ( n46391 ) : ( n46398 ) ;
assign n46400 =  ( n192 ) ? ( VREG_2_7 ) : ( VREG_2_7 ) ;
assign n46401 =  ( n157 ) ? ( n46399 ) : ( n46400 ) ;
assign n46402 =  ( n6 ) ? ( n46386 ) : ( n46401 ) ;
assign n46403 =  ( n439 ) ? ( n46402 ) : ( VREG_2_7 ) ;
assign n46404 =  ( n148 ) ? ( n31660 ) : ( VREG_2_8 ) ;
assign n46405 =  ( n146 ) ? ( n31659 ) : ( n46404 ) ;
assign n46406 =  ( n144 ) ? ( n31658 ) : ( n46405 ) ;
assign n46407 =  ( n142 ) ? ( n31657 ) : ( n46406 ) ;
assign n46408 =  ( n10 ) ? ( n31656 ) : ( n46407 ) ;
assign n46409 =  ( n148 ) ? ( n32694 ) : ( VREG_2_8 ) ;
assign n46410 =  ( n146 ) ? ( n32693 ) : ( n46409 ) ;
assign n46411 =  ( n144 ) ? ( n32692 ) : ( n46410 ) ;
assign n46412 =  ( n142 ) ? ( n32691 ) : ( n46411 ) ;
assign n46413 =  ( n10 ) ? ( n32690 ) : ( n46412 ) ;
assign n46414 =  ( n32701 ) ? ( VREG_2_8 ) : ( n46408 ) ;
assign n46415 =  ( n32701 ) ? ( VREG_2_8 ) : ( n46413 ) ;
assign n46416 =  ( n3034 ) ? ( n46415 ) : ( VREG_2_8 ) ;
assign n46417 =  ( n2965 ) ? ( n46414 ) : ( n46416 ) ;
assign n46418 =  ( n1930 ) ? ( n46413 ) : ( n46417 ) ;
assign n46419 =  ( n879 ) ? ( n46408 ) : ( n46418 ) ;
assign n46420 =  ( n172 ) ? ( n32712 ) : ( VREG_2_8 ) ;
assign n46421 =  ( n170 ) ? ( n32711 ) : ( n46420 ) ;
assign n46422 =  ( n168 ) ? ( n32710 ) : ( n46421 ) ;
assign n46423 =  ( n166 ) ? ( n32709 ) : ( n46422 ) ;
assign n46424 =  ( n162 ) ? ( n32708 ) : ( n46423 ) ;
assign n46425 =  ( n172 ) ? ( n32722 ) : ( VREG_2_8 ) ;
assign n46426 =  ( n170 ) ? ( n32721 ) : ( n46425 ) ;
assign n46427 =  ( n168 ) ? ( n32720 ) : ( n46426 ) ;
assign n46428 =  ( n166 ) ? ( n32719 ) : ( n46427 ) ;
assign n46429 =  ( n162 ) ? ( n32718 ) : ( n46428 ) ;
assign n46430 =  ( n32701 ) ? ( VREG_2_8 ) : ( n46429 ) ;
assign n46431 =  ( n3051 ) ? ( n46430 ) : ( VREG_2_8 ) ;
assign n46432 =  ( n3040 ) ? ( n46424 ) : ( n46431 ) ;
assign n46433 =  ( n192 ) ? ( VREG_2_8 ) : ( VREG_2_8 ) ;
assign n46434 =  ( n157 ) ? ( n46432 ) : ( n46433 ) ;
assign n46435 =  ( n6 ) ? ( n46419 ) : ( n46434 ) ;
assign n46436 =  ( n439 ) ? ( n46435 ) : ( VREG_2_8 ) ;
assign n46437 =  ( n148 ) ? ( n33779 ) : ( VREG_2_9 ) ;
assign n46438 =  ( n146 ) ? ( n33778 ) : ( n46437 ) ;
assign n46439 =  ( n144 ) ? ( n33777 ) : ( n46438 ) ;
assign n46440 =  ( n142 ) ? ( n33776 ) : ( n46439 ) ;
assign n46441 =  ( n10 ) ? ( n33775 ) : ( n46440 ) ;
assign n46442 =  ( n148 ) ? ( n34813 ) : ( VREG_2_9 ) ;
assign n46443 =  ( n146 ) ? ( n34812 ) : ( n46442 ) ;
assign n46444 =  ( n144 ) ? ( n34811 ) : ( n46443 ) ;
assign n46445 =  ( n142 ) ? ( n34810 ) : ( n46444 ) ;
assign n46446 =  ( n10 ) ? ( n34809 ) : ( n46445 ) ;
assign n46447 =  ( n34820 ) ? ( VREG_2_9 ) : ( n46441 ) ;
assign n46448 =  ( n34820 ) ? ( VREG_2_9 ) : ( n46446 ) ;
assign n46449 =  ( n3034 ) ? ( n46448 ) : ( VREG_2_9 ) ;
assign n46450 =  ( n2965 ) ? ( n46447 ) : ( n46449 ) ;
assign n46451 =  ( n1930 ) ? ( n46446 ) : ( n46450 ) ;
assign n46452 =  ( n879 ) ? ( n46441 ) : ( n46451 ) ;
assign n46453 =  ( n172 ) ? ( n34831 ) : ( VREG_2_9 ) ;
assign n46454 =  ( n170 ) ? ( n34830 ) : ( n46453 ) ;
assign n46455 =  ( n168 ) ? ( n34829 ) : ( n46454 ) ;
assign n46456 =  ( n166 ) ? ( n34828 ) : ( n46455 ) ;
assign n46457 =  ( n162 ) ? ( n34827 ) : ( n46456 ) ;
assign n46458 =  ( n172 ) ? ( n34841 ) : ( VREG_2_9 ) ;
assign n46459 =  ( n170 ) ? ( n34840 ) : ( n46458 ) ;
assign n46460 =  ( n168 ) ? ( n34839 ) : ( n46459 ) ;
assign n46461 =  ( n166 ) ? ( n34838 ) : ( n46460 ) ;
assign n46462 =  ( n162 ) ? ( n34837 ) : ( n46461 ) ;
assign n46463 =  ( n34820 ) ? ( VREG_2_9 ) : ( n46462 ) ;
assign n46464 =  ( n3051 ) ? ( n46463 ) : ( VREG_2_9 ) ;
assign n46465 =  ( n3040 ) ? ( n46457 ) : ( n46464 ) ;
assign n46466 =  ( n192 ) ? ( VREG_2_9 ) : ( VREG_2_9 ) ;
assign n46467 =  ( n157 ) ? ( n46465 ) : ( n46466 ) ;
assign n46468 =  ( n6 ) ? ( n46452 ) : ( n46467 ) ;
assign n46469 =  ( n439 ) ? ( n46468 ) : ( VREG_2_9 ) ;
assign n46470 =  ( n148 ) ? ( n1924 ) : ( VREG_30_0 ) ;
assign n46471 =  ( n146 ) ? ( n1923 ) : ( n46470 ) ;
assign n46472 =  ( n144 ) ? ( n1922 ) : ( n46471 ) ;
assign n46473 =  ( n142 ) ? ( n1921 ) : ( n46472 ) ;
assign n46474 =  ( n10 ) ? ( n1920 ) : ( n46473 ) ;
assign n46475 =  ( n148 ) ? ( n2959 ) : ( VREG_30_0 ) ;
assign n46476 =  ( n146 ) ? ( n2958 ) : ( n46475 ) ;
assign n46477 =  ( n144 ) ? ( n2957 ) : ( n46476 ) ;
assign n46478 =  ( n142 ) ? ( n2956 ) : ( n46477 ) ;
assign n46479 =  ( n10 ) ? ( n2955 ) : ( n46478 ) ;
assign n46480 =  ( n3032 ) ? ( VREG_30_0 ) : ( n46474 ) ;
assign n46481 =  ( n3032 ) ? ( VREG_30_0 ) : ( n46479 ) ;
assign n46482 =  ( n3034 ) ? ( n46481 ) : ( VREG_30_0 ) ;
assign n46483 =  ( n2965 ) ? ( n46480 ) : ( n46482 ) ;
assign n46484 =  ( n1930 ) ? ( n46479 ) : ( n46483 ) ;
assign n46485 =  ( n879 ) ? ( n46474 ) : ( n46484 ) ;
assign n46486 =  ( n172 ) ? ( n3045 ) : ( VREG_30_0 ) ;
assign n46487 =  ( n170 ) ? ( n3044 ) : ( n46486 ) ;
assign n46488 =  ( n168 ) ? ( n3043 ) : ( n46487 ) ;
assign n46489 =  ( n166 ) ? ( n3042 ) : ( n46488 ) ;
assign n46490 =  ( n162 ) ? ( n3041 ) : ( n46489 ) ;
assign n46491 =  ( n172 ) ? ( n3056 ) : ( VREG_30_0 ) ;
assign n46492 =  ( n170 ) ? ( n3055 ) : ( n46491 ) ;
assign n46493 =  ( n168 ) ? ( n3054 ) : ( n46492 ) ;
assign n46494 =  ( n166 ) ? ( n3053 ) : ( n46493 ) ;
assign n46495 =  ( n162 ) ? ( n3052 ) : ( n46494 ) ;
assign n46496 =  ( n3032 ) ? ( VREG_30_0 ) : ( n46495 ) ;
assign n46497 =  ( n3051 ) ? ( n46496 ) : ( VREG_30_0 ) ;
assign n46498 =  ( n3040 ) ? ( n46490 ) : ( n46497 ) ;
assign n46499 =  ( n192 ) ? ( VREG_30_0 ) : ( VREG_30_0 ) ;
assign n46500 =  ( n157 ) ? ( n46498 ) : ( n46499 ) ;
assign n46501 =  ( n6 ) ? ( n46485 ) : ( n46500 ) ;
assign n46502 =  ( n703 ) ? ( n46501 ) : ( VREG_30_0 ) ;
assign n46503 =  ( n148 ) ? ( n4113 ) : ( VREG_30_1 ) ;
assign n46504 =  ( n146 ) ? ( n4112 ) : ( n46503 ) ;
assign n46505 =  ( n144 ) ? ( n4111 ) : ( n46504 ) ;
assign n46506 =  ( n142 ) ? ( n4110 ) : ( n46505 ) ;
assign n46507 =  ( n10 ) ? ( n4109 ) : ( n46506 ) ;
assign n46508 =  ( n148 ) ? ( n5147 ) : ( VREG_30_1 ) ;
assign n46509 =  ( n146 ) ? ( n5146 ) : ( n46508 ) ;
assign n46510 =  ( n144 ) ? ( n5145 ) : ( n46509 ) ;
assign n46511 =  ( n142 ) ? ( n5144 ) : ( n46510 ) ;
assign n46512 =  ( n10 ) ? ( n5143 ) : ( n46511 ) ;
assign n46513 =  ( n5154 ) ? ( VREG_30_1 ) : ( n46507 ) ;
assign n46514 =  ( n5154 ) ? ( VREG_30_1 ) : ( n46512 ) ;
assign n46515 =  ( n3034 ) ? ( n46514 ) : ( VREG_30_1 ) ;
assign n46516 =  ( n2965 ) ? ( n46513 ) : ( n46515 ) ;
assign n46517 =  ( n1930 ) ? ( n46512 ) : ( n46516 ) ;
assign n46518 =  ( n879 ) ? ( n46507 ) : ( n46517 ) ;
assign n46519 =  ( n172 ) ? ( n5165 ) : ( VREG_30_1 ) ;
assign n46520 =  ( n170 ) ? ( n5164 ) : ( n46519 ) ;
assign n46521 =  ( n168 ) ? ( n5163 ) : ( n46520 ) ;
assign n46522 =  ( n166 ) ? ( n5162 ) : ( n46521 ) ;
assign n46523 =  ( n162 ) ? ( n5161 ) : ( n46522 ) ;
assign n46524 =  ( n172 ) ? ( n5175 ) : ( VREG_30_1 ) ;
assign n46525 =  ( n170 ) ? ( n5174 ) : ( n46524 ) ;
assign n46526 =  ( n168 ) ? ( n5173 ) : ( n46525 ) ;
assign n46527 =  ( n166 ) ? ( n5172 ) : ( n46526 ) ;
assign n46528 =  ( n162 ) ? ( n5171 ) : ( n46527 ) ;
assign n46529 =  ( n5154 ) ? ( VREG_30_1 ) : ( n46528 ) ;
assign n46530 =  ( n3051 ) ? ( n46529 ) : ( VREG_30_1 ) ;
assign n46531 =  ( n3040 ) ? ( n46523 ) : ( n46530 ) ;
assign n46532 =  ( n192 ) ? ( VREG_30_1 ) : ( VREG_30_1 ) ;
assign n46533 =  ( n157 ) ? ( n46531 ) : ( n46532 ) ;
assign n46534 =  ( n6 ) ? ( n46518 ) : ( n46533 ) ;
assign n46535 =  ( n703 ) ? ( n46534 ) : ( VREG_30_1 ) ;
assign n46536 =  ( n148 ) ? ( n6232 ) : ( VREG_30_10 ) ;
assign n46537 =  ( n146 ) ? ( n6231 ) : ( n46536 ) ;
assign n46538 =  ( n144 ) ? ( n6230 ) : ( n46537 ) ;
assign n46539 =  ( n142 ) ? ( n6229 ) : ( n46538 ) ;
assign n46540 =  ( n10 ) ? ( n6228 ) : ( n46539 ) ;
assign n46541 =  ( n148 ) ? ( n7266 ) : ( VREG_30_10 ) ;
assign n46542 =  ( n146 ) ? ( n7265 ) : ( n46541 ) ;
assign n46543 =  ( n144 ) ? ( n7264 ) : ( n46542 ) ;
assign n46544 =  ( n142 ) ? ( n7263 ) : ( n46543 ) ;
assign n46545 =  ( n10 ) ? ( n7262 ) : ( n46544 ) ;
assign n46546 =  ( n7273 ) ? ( VREG_30_10 ) : ( n46540 ) ;
assign n46547 =  ( n7273 ) ? ( VREG_30_10 ) : ( n46545 ) ;
assign n46548 =  ( n3034 ) ? ( n46547 ) : ( VREG_30_10 ) ;
assign n46549 =  ( n2965 ) ? ( n46546 ) : ( n46548 ) ;
assign n46550 =  ( n1930 ) ? ( n46545 ) : ( n46549 ) ;
assign n46551 =  ( n879 ) ? ( n46540 ) : ( n46550 ) ;
assign n46552 =  ( n172 ) ? ( n7284 ) : ( VREG_30_10 ) ;
assign n46553 =  ( n170 ) ? ( n7283 ) : ( n46552 ) ;
assign n46554 =  ( n168 ) ? ( n7282 ) : ( n46553 ) ;
assign n46555 =  ( n166 ) ? ( n7281 ) : ( n46554 ) ;
assign n46556 =  ( n162 ) ? ( n7280 ) : ( n46555 ) ;
assign n46557 =  ( n172 ) ? ( n7294 ) : ( VREG_30_10 ) ;
assign n46558 =  ( n170 ) ? ( n7293 ) : ( n46557 ) ;
assign n46559 =  ( n168 ) ? ( n7292 ) : ( n46558 ) ;
assign n46560 =  ( n166 ) ? ( n7291 ) : ( n46559 ) ;
assign n46561 =  ( n162 ) ? ( n7290 ) : ( n46560 ) ;
assign n46562 =  ( n7273 ) ? ( VREG_30_10 ) : ( n46561 ) ;
assign n46563 =  ( n3051 ) ? ( n46562 ) : ( VREG_30_10 ) ;
assign n46564 =  ( n3040 ) ? ( n46556 ) : ( n46563 ) ;
assign n46565 =  ( n192 ) ? ( VREG_30_10 ) : ( VREG_30_10 ) ;
assign n46566 =  ( n157 ) ? ( n46564 ) : ( n46565 ) ;
assign n46567 =  ( n6 ) ? ( n46551 ) : ( n46566 ) ;
assign n46568 =  ( n703 ) ? ( n46567 ) : ( VREG_30_10 ) ;
assign n46569 =  ( n148 ) ? ( n8351 ) : ( VREG_30_11 ) ;
assign n46570 =  ( n146 ) ? ( n8350 ) : ( n46569 ) ;
assign n46571 =  ( n144 ) ? ( n8349 ) : ( n46570 ) ;
assign n46572 =  ( n142 ) ? ( n8348 ) : ( n46571 ) ;
assign n46573 =  ( n10 ) ? ( n8347 ) : ( n46572 ) ;
assign n46574 =  ( n148 ) ? ( n9385 ) : ( VREG_30_11 ) ;
assign n46575 =  ( n146 ) ? ( n9384 ) : ( n46574 ) ;
assign n46576 =  ( n144 ) ? ( n9383 ) : ( n46575 ) ;
assign n46577 =  ( n142 ) ? ( n9382 ) : ( n46576 ) ;
assign n46578 =  ( n10 ) ? ( n9381 ) : ( n46577 ) ;
assign n46579 =  ( n9392 ) ? ( VREG_30_11 ) : ( n46573 ) ;
assign n46580 =  ( n9392 ) ? ( VREG_30_11 ) : ( n46578 ) ;
assign n46581 =  ( n3034 ) ? ( n46580 ) : ( VREG_30_11 ) ;
assign n46582 =  ( n2965 ) ? ( n46579 ) : ( n46581 ) ;
assign n46583 =  ( n1930 ) ? ( n46578 ) : ( n46582 ) ;
assign n46584 =  ( n879 ) ? ( n46573 ) : ( n46583 ) ;
assign n46585 =  ( n172 ) ? ( n9403 ) : ( VREG_30_11 ) ;
assign n46586 =  ( n170 ) ? ( n9402 ) : ( n46585 ) ;
assign n46587 =  ( n168 ) ? ( n9401 ) : ( n46586 ) ;
assign n46588 =  ( n166 ) ? ( n9400 ) : ( n46587 ) ;
assign n46589 =  ( n162 ) ? ( n9399 ) : ( n46588 ) ;
assign n46590 =  ( n172 ) ? ( n9413 ) : ( VREG_30_11 ) ;
assign n46591 =  ( n170 ) ? ( n9412 ) : ( n46590 ) ;
assign n46592 =  ( n168 ) ? ( n9411 ) : ( n46591 ) ;
assign n46593 =  ( n166 ) ? ( n9410 ) : ( n46592 ) ;
assign n46594 =  ( n162 ) ? ( n9409 ) : ( n46593 ) ;
assign n46595 =  ( n9392 ) ? ( VREG_30_11 ) : ( n46594 ) ;
assign n46596 =  ( n3051 ) ? ( n46595 ) : ( VREG_30_11 ) ;
assign n46597 =  ( n3040 ) ? ( n46589 ) : ( n46596 ) ;
assign n46598 =  ( n192 ) ? ( VREG_30_11 ) : ( VREG_30_11 ) ;
assign n46599 =  ( n157 ) ? ( n46597 ) : ( n46598 ) ;
assign n46600 =  ( n6 ) ? ( n46584 ) : ( n46599 ) ;
assign n46601 =  ( n703 ) ? ( n46600 ) : ( VREG_30_11 ) ;
assign n46602 =  ( n148 ) ? ( n10470 ) : ( VREG_30_12 ) ;
assign n46603 =  ( n146 ) ? ( n10469 ) : ( n46602 ) ;
assign n46604 =  ( n144 ) ? ( n10468 ) : ( n46603 ) ;
assign n46605 =  ( n142 ) ? ( n10467 ) : ( n46604 ) ;
assign n46606 =  ( n10 ) ? ( n10466 ) : ( n46605 ) ;
assign n46607 =  ( n148 ) ? ( n11504 ) : ( VREG_30_12 ) ;
assign n46608 =  ( n146 ) ? ( n11503 ) : ( n46607 ) ;
assign n46609 =  ( n144 ) ? ( n11502 ) : ( n46608 ) ;
assign n46610 =  ( n142 ) ? ( n11501 ) : ( n46609 ) ;
assign n46611 =  ( n10 ) ? ( n11500 ) : ( n46610 ) ;
assign n46612 =  ( n11511 ) ? ( VREG_30_12 ) : ( n46606 ) ;
assign n46613 =  ( n11511 ) ? ( VREG_30_12 ) : ( n46611 ) ;
assign n46614 =  ( n3034 ) ? ( n46613 ) : ( VREG_30_12 ) ;
assign n46615 =  ( n2965 ) ? ( n46612 ) : ( n46614 ) ;
assign n46616 =  ( n1930 ) ? ( n46611 ) : ( n46615 ) ;
assign n46617 =  ( n879 ) ? ( n46606 ) : ( n46616 ) ;
assign n46618 =  ( n172 ) ? ( n11522 ) : ( VREG_30_12 ) ;
assign n46619 =  ( n170 ) ? ( n11521 ) : ( n46618 ) ;
assign n46620 =  ( n168 ) ? ( n11520 ) : ( n46619 ) ;
assign n46621 =  ( n166 ) ? ( n11519 ) : ( n46620 ) ;
assign n46622 =  ( n162 ) ? ( n11518 ) : ( n46621 ) ;
assign n46623 =  ( n172 ) ? ( n11532 ) : ( VREG_30_12 ) ;
assign n46624 =  ( n170 ) ? ( n11531 ) : ( n46623 ) ;
assign n46625 =  ( n168 ) ? ( n11530 ) : ( n46624 ) ;
assign n46626 =  ( n166 ) ? ( n11529 ) : ( n46625 ) ;
assign n46627 =  ( n162 ) ? ( n11528 ) : ( n46626 ) ;
assign n46628 =  ( n11511 ) ? ( VREG_30_12 ) : ( n46627 ) ;
assign n46629 =  ( n3051 ) ? ( n46628 ) : ( VREG_30_12 ) ;
assign n46630 =  ( n3040 ) ? ( n46622 ) : ( n46629 ) ;
assign n46631 =  ( n192 ) ? ( VREG_30_12 ) : ( VREG_30_12 ) ;
assign n46632 =  ( n157 ) ? ( n46630 ) : ( n46631 ) ;
assign n46633 =  ( n6 ) ? ( n46617 ) : ( n46632 ) ;
assign n46634 =  ( n703 ) ? ( n46633 ) : ( VREG_30_12 ) ;
assign n46635 =  ( n148 ) ? ( n12589 ) : ( VREG_30_13 ) ;
assign n46636 =  ( n146 ) ? ( n12588 ) : ( n46635 ) ;
assign n46637 =  ( n144 ) ? ( n12587 ) : ( n46636 ) ;
assign n46638 =  ( n142 ) ? ( n12586 ) : ( n46637 ) ;
assign n46639 =  ( n10 ) ? ( n12585 ) : ( n46638 ) ;
assign n46640 =  ( n148 ) ? ( n13623 ) : ( VREG_30_13 ) ;
assign n46641 =  ( n146 ) ? ( n13622 ) : ( n46640 ) ;
assign n46642 =  ( n144 ) ? ( n13621 ) : ( n46641 ) ;
assign n46643 =  ( n142 ) ? ( n13620 ) : ( n46642 ) ;
assign n46644 =  ( n10 ) ? ( n13619 ) : ( n46643 ) ;
assign n46645 =  ( n13630 ) ? ( VREG_30_13 ) : ( n46639 ) ;
assign n46646 =  ( n13630 ) ? ( VREG_30_13 ) : ( n46644 ) ;
assign n46647 =  ( n3034 ) ? ( n46646 ) : ( VREG_30_13 ) ;
assign n46648 =  ( n2965 ) ? ( n46645 ) : ( n46647 ) ;
assign n46649 =  ( n1930 ) ? ( n46644 ) : ( n46648 ) ;
assign n46650 =  ( n879 ) ? ( n46639 ) : ( n46649 ) ;
assign n46651 =  ( n172 ) ? ( n13641 ) : ( VREG_30_13 ) ;
assign n46652 =  ( n170 ) ? ( n13640 ) : ( n46651 ) ;
assign n46653 =  ( n168 ) ? ( n13639 ) : ( n46652 ) ;
assign n46654 =  ( n166 ) ? ( n13638 ) : ( n46653 ) ;
assign n46655 =  ( n162 ) ? ( n13637 ) : ( n46654 ) ;
assign n46656 =  ( n172 ) ? ( n13651 ) : ( VREG_30_13 ) ;
assign n46657 =  ( n170 ) ? ( n13650 ) : ( n46656 ) ;
assign n46658 =  ( n168 ) ? ( n13649 ) : ( n46657 ) ;
assign n46659 =  ( n166 ) ? ( n13648 ) : ( n46658 ) ;
assign n46660 =  ( n162 ) ? ( n13647 ) : ( n46659 ) ;
assign n46661 =  ( n13630 ) ? ( VREG_30_13 ) : ( n46660 ) ;
assign n46662 =  ( n3051 ) ? ( n46661 ) : ( VREG_30_13 ) ;
assign n46663 =  ( n3040 ) ? ( n46655 ) : ( n46662 ) ;
assign n46664 =  ( n192 ) ? ( VREG_30_13 ) : ( VREG_30_13 ) ;
assign n46665 =  ( n157 ) ? ( n46663 ) : ( n46664 ) ;
assign n46666 =  ( n6 ) ? ( n46650 ) : ( n46665 ) ;
assign n46667 =  ( n703 ) ? ( n46666 ) : ( VREG_30_13 ) ;
assign n46668 =  ( n148 ) ? ( n14708 ) : ( VREG_30_14 ) ;
assign n46669 =  ( n146 ) ? ( n14707 ) : ( n46668 ) ;
assign n46670 =  ( n144 ) ? ( n14706 ) : ( n46669 ) ;
assign n46671 =  ( n142 ) ? ( n14705 ) : ( n46670 ) ;
assign n46672 =  ( n10 ) ? ( n14704 ) : ( n46671 ) ;
assign n46673 =  ( n148 ) ? ( n15742 ) : ( VREG_30_14 ) ;
assign n46674 =  ( n146 ) ? ( n15741 ) : ( n46673 ) ;
assign n46675 =  ( n144 ) ? ( n15740 ) : ( n46674 ) ;
assign n46676 =  ( n142 ) ? ( n15739 ) : ( n46675 ) ;
assign n46677 =  ( n10 ) ? ( n15738 ) : ( n46676 ) ;
assign n46678 =  ( n15749 ) ? ( VREG_30_14 ) : ( n46672 ) ;
assign n46679 =  ( n15749 ) ? ( VREG_30_14 ) : ( n46677 ) ;
assign n46680 =  ( n3034 ) ? ( n46679 ) : ( VREG_30_14 ) ;
assign n46681 =  ( n2965 ) ? ( n46678 ) : ( n46680 ) ;
assign n46682 =  ( n1930 ) ? ( n46677 ) : ( n46681 ) ;
assign n46683 =  ( n879 ) ? ( n46672 ) : ( n46682 ) ;
assign n46684 =  ( n172 ) ? ( n15760 ) : ( VREG_30_14 ) ;
assign n46685 =  ( n170 ) ? ( n15759 ) : ( n46684 ) ;
assign n46686 =  ( n168 ) ? ( n15758 ) : ( n46685 ) ;
assign n46687 =  ( n166 ) ? ( n15757 ) : ( n46686 ) ;
assign n46688 =  ( n162 ) ? ( n15756 ) : ( n46687 ) ;
assign n46689 =  ( n172 ) ? ( n15770 ) : ( VREG_30_14 ) ;
assign n46690 =  ( n170 ) ? ( n15769 ) : ( n46689 ) ;
assign n46691 =  ( n168 ) ? ( n15768 ) : ( n46690 ) ;
assign n46692 =  ( n166 ) ? ( n15767 ) : ( n46691 ) ;
assign n46693 =  ( n162 ) ? ( n15766 ) : ( n46692 ) ;
assign n46694 =  ( n15749 ) ? ( VREG_30_14 ) : ( n46693 ) ;
assign n46695 =  ( n3051 ) ? ( n46694 ) : ( VREG_30_14 ) ;
assign n46696 =  ( n3040 ) ? ( n46688 ) : ( n46695 ) ;
assign n46697 =  ( n192 ) ? ( VREG_30_14 ) : ( VREG_30_14 ) ;
assign n46698 =  ( n157 ) ? ( n46696 ) : ( n46697 ) ;
assign n46699 =  ( n6 ) ? ( n46683 ) : ( n46698 ) ;
assign n46700 =  ( n703 ) ? ( n46699 ) : ( VREG_30_14 ) ;
assign n46701 =  ( n148 ) ? ( n16827 ) : ( VREG_30_15 ) ;
assign n46702 =  ( n146 ) ? ( n16826 ) : ( n46701 ) ;
assign n46703 =  ( n144 ) ? ( n16825 ) : ( n46702 ) ;
assign n46704 =  ( n142 ) ? ( n16824 ) : ( n46703 ) ;
assign n46705 =  ( n10 ) ? ( n16823 ) : ( n46704 ) ;
assign n46706 =  ( n148 ) ? ( n17861 ) : ( VREG_30_15 ) ;
assign n46707 =  ( n146 ) ? ( n17860 ) : ( n46706 ) ;
assign n46708 =  ( n144 ) ? ( n17859 ) : ( n46707 ) ;
assign n46709 =  ( n142 ) ? ( n17858 ) : ( n46708 ) ;
assign n46710 =  ( n10 ) ? ( n17857 ) : ( n46709 ) ;
assign n46711 =  ( n17868 ) ? ( VREG_30_15 ) : ( n46705 ) ;
assign n46712 =  ( n17868 ) ? ( VREG_30_15 ) : ( n46710 ) ;
assign n46713 =  ( n3034 ) ? ( n46712 ) : ( VREG_30_15 ) ;
assign n46714 =  ( n2965 ) ? ( n46711 ) : ( n46713 ) ;
assign n46715 =  ( n1930 ) ? ( n46710 ) : ( n46714 ) ;
assign n46716 =  ( n879 ) ? ( n46705 ) : ( n46715 ) ;
assign n46717 =  ( n172 ) ? ( n17879 ) : ( VREG_30_15 ) ;
assign n46718 =  ( n170 ) ? ( n17878 ) : ( n46717 ) ;
assign n46719 =  ( n168 ) ? ( n17877 ) : ( n46718 ) ;
assign n46720 =  ( n166 ) ? ( n17876 ) : ( n46719 ) ;
assign n46721 =  ( n162 ) ? ( n17875 ) : ( n46720 ) ;
assign n46722 =  ( n172 ) ? ( n17889 ) : ( VREG_30_15 ) ;
assign n46723 =  ( n170 ) ? ( n17888 ) : ( n46722 ) ;
assign n46724 =  ( n168 ) ? ( n17887 ) : ( n46723 ) ;
assign n46725 =  ( n166 ) ? ( n17886 ) : ( n46724 ) ;
assign n46726 =  ( n162 ) ? ( n17885 ) : ( n46725 ) ;
assign n46727 =  ( n17868 ) ? ( VREG_30_15 ) : ( n46726 ) ;
assign n46728 =  ( n3051 ) ? ( n46727 ) : ( VREG_30_15 ) ;
assign n46729 =  ( n3040 ) ? ( n46721 ) : ( n46728 ) ;
assign n46730 =  ( n192 ) ? ( VREG_30_15 ) : ( VREG_30_15 ) ;
assign n46731 =  ( n157 ) ? ( n46729 ) : ( n46730 ) ;
assign n46732 =  ( n6 ) ? ( n46716 ) : ( n46731 ) ;
assign n46733 =  ( n703 ) ? ( n46732 ) : ( VREG_30_15 ) ;
assign n46734 =  ( n148 ) ? ( n18946 ) : ( VREG_30_2 ) ;
assign n46735 =  ( n146 ) ? ( n18945 ) : ( n46734 ) ;
assign n46736 =  ( n144 ) ? ( n18944 ) : ( n46735 ) ;
assign n46737 =  ( n142 ) ? ( n18943 ) : ( n46736 ) ;
assign n46738 =  ( n10 ) ? ( n18942 ) : ( n46737 ) ;
assign n46739 =  ( n148 ) ? ( n19980 ) : ( VREG_30_2 ) ;
assign n46740 =  ( n146 ) ? ( n19979 ) : ( n46739 ) ;
assign n46741 =  ( n144 ) ? ( n19978 ) : ( n46740 ) ;
assign n46742 =  ( n142 ) ? ( n19977 ) : ( n46741 ) ;
assign n46743 =  ( n10 ) ? ( n19976 ) : ( n46742 ) ;
assign n46744 =  ( n19987 ) ? ( VREG_30_2 ) : ( n46738 ) ;
assign n46745 =  ( n19987 ) ? ( VREG_30_2 ) : ( n46743 ) ;
assign n46746 =  ( n3034 ) ? ( n46745 ) : ( VREG_30_2 ) ;
assign n46747 =  ( n2965 ) ? ( n46744 ) : ( n46746 ) ;
assign n46748 =  ( n1930 ) ? ( n46743 ) : ( n46747 ) ;
assign n46749 =  ( n879 ) ? ( n46738 ) : ( n46748 ) ;
assign n46750 =  ( n172 ) ? ( n19998 ) : ( VREG_30_2 ) ;
assign n46751 =  ( n170 ) ? ( n19997 ) : ( n46750 ) ;
assign n46752 =  ( n168 ) ? ( n19996 ) : ( n46751 ) ;
assign n46753 =  ( n166 ) ? ( n19995 ) : ( n46752 ) ;
assign n46754 =  ( n162 ) ? ( n19994 ) : ( n46753 ) ;
assign n46755 =  ( n172 ) ? ( n20008 ) : ( VREG_30_2 ) ;
assign n46756 =  ( n170 ) ? ( n20007 ) : ( n46755 ) ;
assign n46757 =  ( n168 ) ? ( n20006 ) : ( n46756 ) ;
assign n46758 =  ( n166 ) ? ( n20005 ) : ( n46757 ) ;
assign n46759 =  ( n162 ) ? ( n20004 ) : ( n46758 ) ;
assign n46760 =  ( n19987 ) ? ( VREG_30_2 ) : ( n46759 ) ;
assign n46761 =  ( n3051 ) ? ( n46760 ) : ( VREG_30_2 ) ;
assign n46762 =  ( n3040 ) ? ( n46754 ) : ( n46761 ) ;
assign n46763 =  ( n192 ) ? ( VREG_30_2 ) : ( VREG_30_2 ) ;
assign n46764 =  ( n157 ) ? ( n46762 ) : ( n46763 ) ;
assign n46765 =  ( n6 ) ? ( n46749 ) : ( n46764 ) ;
assign n46766 =  ( n703 ) ? ( n46765 ) : ( VREG_30_2 ) ;
assign n46767 =  ( n148 ) ? ( n21065 ) : ( VREG_30_3 ) ;
assign n46768 =  ( n146 ) ? ( n21064 ) : ( n46767 ) ;
assign n46769 =  ( n144 ) ? ( n21063 ) : ( n46768 ) ;
assign n46770 =  ( n142 ) ? ( n21062 ) : ( n46769 ) ;
assign n46771 =  ( n10 ) ? ( n21061 ) : ( n46770 ) ;
assign n46772 =  ( n148 ) ? ( n22099 ) : ( VREG_30_3 ) ;
assign n46773 =  ( n146 ) ? ( n22098 ) : ( n46772 ) ;
assign n46774 =  ( n144 ) ? ( n22097 ) : ( n46773 ) ;
assign n46775 =  ( n142 ) ? ( n22096 ) : ( n46774 ) ;
assign n46776 =  ( n10 ) ? ( n22095 ) : ( n46775 ) ;
assign n46777 =  ( n22106 ) ? ( VREG_30_3 ) : ( n46771 ) ;
assign n46778 =  ( n22106 ) ? ( VREG_30_3 ) : ( n46776 ) ;
assign n46779 =  ( n3034 ) ? ( n46778 ) : ( VREG_30_3 ) ;
assign n46780 =  ( n2965 ) ? ( n46777 ) : ( n46779 ) ;
assign n46781 =  ( n1930 ) ? ( n46776 ) : ( n46780 ) ;
assign n46782 =  ( n879 ) ? ( n46771 ) : ( n46781 ) ;
assign n46783 =  ( n172 ) ? ( n22117 ) : ( VREG_30_3 ) ;
assign n46784 =  ( n170 ) ? ( n22116 ) : ( n46783 ) ;
assign n46785 =  ( n168 ) ? ( n22115 ) : ( n46784 ) ;
assign n46786 =  ( n166 ) ? ( n22114 ) : ( n46785 ) ;
assign n46787 =  ( n162 ) ? ( n22113 ) : ( n46786 ) ;
assign n46788 =  ( n172 ) ? ( n22127 ) : ( VREG_30_3 ) ;
assign n46789 =  ( n170 ) ? ( n22126 ) : ( n46788 ) ;
assign n46790 =  ( n168 ) ? ( n22125 ) : ( n46789 ) ;
assign n46791 =  ( n166 ) ? ( n22124 ) : ( n46790 ) ;
assign n46792 =  ( n162 ) ? ( n22123 ) : ( n46791 ) ;
assign n46793 =  ( n22106 ) ? ( VREG_30_3 ) : ( n46792 ) ;
assign n46794 =  ( n3051 ) ? ( n46793 ) : ( VREG_30_3 ) ;
assign n46795 =  ( n3040 ) ? ( n46787 ) : ( n46794 ) ;
assign n46796 =  ( n192 ) ? ( VREG_30_3 ) : ( VREG_30_3 ) ;
assign n46797 =  ( n157 ) ? ( n46795 ) : ( n46796 ) ;
assign n46798 =  ( n6 ) ? ( n46782 ) : ( n46797 ) ;
assign n46799 =  ( n703 ) ? ( n46798 ) : ( VREG_30_3 ) ;
assign n46800 =  ( n148 ) ? ( n23184 ) : ( VREG_30_4 ) ;
assign n46801 =  ( n146 ) ? ( n23183 ) : ( n46800 ) ;
assign n46802 =  ( n144 ) ? ( n23182 ) : ( n46801 ) ;
assign n46803 =  ( n142 ) ? ( n23181 ) : ( n46802 ) ;
assign n46804 =  ( n10 ) ? ( n23180 ) : ( n46803 ) ;
assign n46805 =  ( n148 ) ? ( n24218 ) : ( VREG_30_4 ) ;
assign n46806 =  ( n146 ) ? ( n24217 ) : ( n46805 ) ;
assign n46807 =  ( n144 ) ? ( n24216 ) : ( n46806 ) ;
assign n46808 =  ( n142 ) ? ( n24215 ) : ( n46807 ) ;
assign n46809 =  ( n10 ) ? ( n24214 ) : ( n46808 ) ;
assign n46810 =  ( n24225 ) ? ( VREG_30_4 ) : ( n46804 ) ;
assign n46811 =  ( n24225 ) ? ( VREG_30_4 ) : ( n46809 ) ;
assign n46812 =  ( n3034 ) ? ( n46811 ) : ( VREG_30_4 ) ;
assign n46813 =  ( n2965 ) ? ( n46810 ) : ( n46812 ) ;
assign n46814 =  ( n1930 ) ? ( n46809 ) : ( n46813 ) ;
assign n46815 =  ( n879 ) ? ( n46804 ) : ( n46814 ) ;
assign n46816 =  ( n172 ) ? ( n24236 ) : ( VREG_30_4 ) ;
assign n46817 =  ( n170 ) ? ( n24235 ) : ( n46816 ) ;
assign n46818 =  ( n168 ) ? ( n24234 ) : ( n46817 ) ;
assign n46819 =  ( n166 ) ? ( n24233 ) : ( n46818 ) ;
assign n46820 =  ( n162 ) ? ( n24232 ) : ( n46819 ) ;
assign n46821 =  ( n172 ) ? ( n24246 ) : ( VREG_30_4 ) ;
assign n46822 =  ( n170 ) ? ( n24245 ) : ( n46821 ) ;
assign n46823 =  ( n168 ) ? ( n24244 ) : ( n46822 ) ;
assign n46824 =  ( n166 ) ? ( n24243 ) : ( n46823 ) ;
assign n46825 =  ( n162 ) ? ( n24242 ) : ( n46824 ) ;
assign n46826 =  ( n24225 ) ? ( VREG_30_4 ) : ( n46825 ) ;
assign n46827 =  ( n3051 ) ? ( n46826 ) : ( VREG_30_4 ) ;
assign n46828 =  ( n3040 ) ? ( n46820 ) : ( n46827 ) ;
assign n46829 =  ( n192 ) ? ( VREG_30_4 ) : ( VREG_30_4 ) ;
assign n46830 =  ( n157 ) ? ( n46828 ) : ( n46829 ) ;
assign n46831 =  ( n6 ) ? ( n46815 ) : ( n46830 ) ;
assign n46832 =  ( n703 ) ? ( n46831 ) : ( VREG_30_4 ) ;
assign n46833 =  ( n148 ) ? ( n25303 ) : ( VREG_30_5 ) ;
assign n46834 =  ( n146 ) ? ( n25302 ) : ( n46833 ) ;
assign n46835 =  ( n144 ) ? ( n25301 ) : ( n46834 ) ;
assign n46836 =  ( n142 ) ? ( n25300 ) : ( n46835 ) ;
assign n46837 =  ( n10 ) ? ( n25299 ) : ( n46836 ) ;
assign n46838 =  ( n148 ) ? ( n26337 ) : ( VREG_30_5 ) ;
assign n46839 =  ( n146 ) ? ( n26336 ) : ( n46838 ) ;
assign n46840 =  ( n144 ) ? ( n26335 ) : ( n46839 ) ;
assign n46841 =  ( n142 ) ? ( n26334 ) : ( n46840 ) ;
assign n46842 =  ( n10 ) ? ( n26333 ) : ( n46841 ) ;
assign n46843 =  ( n26344 ) ? ( VREG_30_5 ) : ( n46837 ) ;
assign n46844 =  ( n26344 ) ? ( VREG_30_5 ) : ( n46842 ) ;
assign n46845 =  ( n3034 ) ? ( n46844 ) : ( VREG_30_5 ) ;
assign n46846 =  ( n2965 ) ? ( n46843 ) : ( n46845 ) ;
assign n46847 =  ( n1930 ) ? ( n46842 ) : ( n46846 ) ;
assign n46848 =  ( n879 ) ? ( n46837 ) : ( n46847 ) ;
assign n46849 =  ( n172 ) ? ( n26355 ) : ( VREG_30_5 ) ;
assign n46850 =  ( n170 ) ? ( n26354 ) : ( n46849 ) ;
assign n46851 =  ( n168 ) ? ( n26353 ) : ( n46850 ) ;
assign n46852 =  ( n166 ) ? ( n26352 ) : ( n46851 ) ;
assign n46853 =  ( n162 ) ? ( n26351 ) : ( n46852 ) ;
assign n46854 =  ( n172 ) ? ( n26365 ) : ( VREG_30_5 ) ;
assign n46855 =  ( n170 ) ? ( n26364 ) : ( n46854 ) ;
assign n46856 =  ( n168 ) ? ( n26363 ) : ( n46855 ) ;
assign n46857 =  ( n166 ) ? ( n26362 ) : ( n46856 ) ;
assign n46858 =  ( n162 ) ? ( n26361 ) : ( n46857 ) ;
assign n46859 =  ( n26344 ) ? ( VREG_30_5 ) : ( n46858 ) ;
assign n46860 =  ( n3051 ) ? ( n46859 ) : ( VREG_30_5 ) ;
assign n46861 =  ( n3040 ) ? ( n46853 ) : ( n46860 ) ;
assign n46862 =  ( n192 ) ? ( VREG_30_5 ) : ( VREG_30_5 ) ;
assign n46863 =  ( n157 ) ? ( n46861 ) : ( n46862 ) ;
assign n46864 =  ( n6 ) ? ( n46848 ) : ( n46863 ) ;
assign n46865 =  ( n703 ) ? ( n46864 ) : ( VREG_30_5 ) ;
assign n46866 =  ( n148 ) ? ( n27422 ) : ( VREG_30_6 ) ;
assign n46867 =  ( n146 ) ? ( n27421 ) : ( n46866 ) ;
assign n46868 =  ( n144 ) ? ( n27420 ) : ( n46867 ) ;
assign n46869 =  ( n142 ) ? ( n27419 ) : ( n46868 ) ;
assign n46870 =  ( n10 ) ? ( n27418 ) : ( n46869 ) ;
assign n46871 =  ( n148 ) ? ( n28456 ) : ( VREG_30_6 ) ;
assign n46872 =  ( n146 ) ? ( n28455 ) : ( n46871 ) ;
assign n46873 =  ( n144 ) ? ( n28454 ) : ( n46872 ) ;
assign n46874 =  ( n142 ) ? ( n28453 ) : ( n46873 ) ;
assign n46875 =  ( n10 ) ? ( n28452 ) : ( n46874 ) ;
assign n46876 =  ( n28463 ) ? ( VREG_30_6 ) : ( n46870 ) ;
assign n46877 =  ( n28463 ) ? ( VREG_30_6 ) : ( n46875 ) ;
assign n46878 =  ( n3034 ) ? ( n46877 ) : ( VREG_30_6 ) ;
assign n46879 =  ( n2965 ) ? ( n46876 ) : ( n46878 ) ;
assign n46880 =  ( n1930 ) ? ( n46875 ) : ( n46879 ) ;
assign n46881 =  ( n879 ) ? ( n46870 ) : ( n46880 ) ;
assign n46882 =  ( n172 ) ? ( n28474 ) : ( VREG_30_6 ) ;
assign n46883 =  ( n170 ) ? ( n28473 ) : ( n46882 ) ;
assign n46884 =  ( n168 ) ? ( n28472 ) : ( n46883 ) ;
assign n46885 =  ( n166 ) ? ( n28471 ) : ( n46884 ) ;
assign n46886 =  ( n162 ) ? ( n28470 ) : ( n46885 ) ;
assign n46887 =  ( n172 ) ? ( n28484 ) : ( VREG_30_6 ) ;
assign n46888 =  ( n170 ) ? ( n28483 ) : ( n46887 ) ;
assign n46889 =  ( n168 ) ? ( n28482 ) : ( n46888 ) ;
assign n46890 =  ( n166 ) ? ( n28481 ) : ( n46889 ) ;
assign n46891 =  ( n162 ) ? ( n28480 ) : ( n46890 ) ;
assign n46892 =  ( n28463 ) ? ( VREG_30_6 ) : ( n46891 ) ;
assign n46893 =  ( n3051 ) ? ( n46892 ) : ( VREG_30_6 ) ;
assign n46894 =  ( n3040 ) ? ( n46886 ) : ( n46893 ) ;
assign n46895 =  ( n192 ) ? ( VREG_30_6 ) : ( VREG_30_6 ) ;
assign n46896 =  ( n157 ) ? ( n46894 ) : ( n46895 ) ;
assign n46897 =  ( n6 ) ? ( n46881 ) : ( n46896 ) ;
assign n46898 =  ( n703 ) ? ( n46897 ) : ( VREG_30_6 ) ;
assign n46899 =  ( n148 ) ? ( n29541 ) : ( VREG_30_7 ) ;
assign n46900 =  ( n146 ) ? ( n29540 ) : ( n46899 ) ;
assign n46901 =  ( n144 ) ? ( n29539 ) : ( n46900 ) ;
assign n46902 =  ( n142 ) ? ( n29538 ) : ( n46901 ) ;
assign n46903 =  ( n10 ) ? ( n29537 ) : ( n46902 ) ;
assign n46904 =  ( n148 ) ? ( n30575 ) : ( VREG_30_7 ) ;
assign n46905 =  ( n146 ) ? ( n30574 ) : ( n46904 ) ;
assign n46906 =  ( n144 ) ? ( n30573 ) : ( n46905 ) ;
assign n46907 =  ( n142 ) ? ( n30572 ) : ( n46906 ) ;
assign n46908 =  ( n10 ) ? ( n30571 ) : ( n46907 ) ;
assign n46909 =  ( n30582 ) ? ( VREG_30_7 ) : ( n46903 ) ;
assign n46910 =  ( n30582 ) ? ( VREG_30_7 ) : ( n46908 ) ;
assign n46911 =  ( n3034 ) ? ( n46910 ) : ( VREG_30_7 ) ;
assign n46912 =  ( n2965 ) ? ( n46909 ) : ( n46911 ) ;
assign n46913 =  ( n1930 ) ? ( n46908 ) : ( n46912 ) ;
assign n46914 =  ( n879 ) ? ( n46903 ) : ( n46913 ) ;
assign n46915 =  ( n172 ) ? ( n30593 ) : ( VREG_30_7 ) ;
assign n46916 =  ( n170 ) ? ( n30592 ) : ( n46915 ) ;
assign n46917 =  ( n168 ) ? ( n30591 ) : ( n46916 ) ;
assign n46918 =  ( n166 ) ? ( n30590 ) : ( n46917 ) ;
assign n46919 =  ( n162 ) ? ( n30589 ) : ( n46918 ) ;
assign n46920 =  ( n172 ) ? ( n30603 ) : ( VREG_30_7 ) ;
assign n46921 =  ( n170 ) ? ( n30602 ) : ( n46920 ) ;
assign n46922 =  ( n168 ) ? ( n30601 ) : ( n46921 ) ;
assign n46923 =  ( n166 ) ? ( n30600 ) : ( n46922 ) ;
assign n46924 =  ( n162 ) ? ( n30599 ) : ( n46923 ) ;
assign n46925 =  ( n30582 ) ? ( VREG_30_7 ) : ( n46924 ) ;
assign n46926 =  ( n3051 ) ? ( n46925 ) : ( VREG_30_7 ) ;
assign n46927 =  ( n3040 ) ? ( n46919 ) : ( n46926 ) ;
assign n46928 =  ( n192 ) ? ( VREG_30_7 ) : ( VREG_30_7 ) ;
assign n46929 =  ( n157 ) ? ( n46927 ) : ( n46928 ) ;
assign n46930 =  ( n6 ) ? ( n46914 ) : ( n46929 ) ;
assign n46931 =  ( n703 ) ? ( n46930 ) : ( VREG_30_7 ) ;
assign n46932 =  ( n148 ) ? ( n31660 ) : ( VREG_30_8 ) ;
assign n46933 =  ( n146 ) ? ( n31659 ) : ( n46932 ) ;
assign n46934 =  ( n144 ) ? ( n31658 ) : ( n46933 ) ;
assign n46935 =  ( n142 ) ? ( n31657 ) : ( n46934 ) ;
assign n46936 =  ( n10 ) ? ( n31656 ) : ( n46935 ) ;
assign n46937 =  ( n148 ) ? ( n32694 ) : ( VREG_30_8 ) ;
assign n46938 =  ( n146 ) ? ( n32693 ) : ( n46937 ) ;
assign n46939 =  ( n144 ) ? ( n32692 ) : ( n46938 ) ;
assign n46940 =  ( n142 ) ? ( n32691 ) : ( n46939 ) ;
assign n46941 =  ( n10 ) ? ( n32690 ) : ( n46940 ) ;
assign n46942 =  ( n32701 ) ? ( VREG_30_8 ) : ( n46936 ) ;
assign n46943 =  ( n32701 ) ? ( VREG_30_8 ) : ( n46941 ) ;
assign n46944 =  ( n3034 ) ? ( n46943 ) : ( VREG_30_8 ) ;
assign n46945 =  ( n2965 ) ? ( n46942 ) : ( n46944 ) ;
assign n46946 =  ( n1930 ) ? ( n46941 ) : ( n46945 ) ;
assign n46947 =  ( n879 ) ? ( n46936 ) : ( n46946 ) ;
assign n46948 =  ( n172 ) ? ( n32712 ) : ( VREG_30_8 ) ;
assign n46949 =  ( n170 ) ? ( n32711 ) : ( n46948 ) ;
assign n46950 =  ( n168 ) ? ( n32710 ) : ( n46949 ) ;
assign n46951 =  ( n166 ) ? ( n32709 ) : ( n46950 ) ;
assign n46952 =  ( n162 ) ? ( n32708 ) : ( n46951 ) ;
assign n46953 =  ( n172 ) ? ( n32722 ) : ( VREG_30_8 ) ;
assign n46954 =  ( n170 ) ? ( n32721 ) : ( n46953 ) ;
assign n46955 =  ( n168 ) ? ( n32720 ) : ( n46954 ) ;
assign n46956 =  ( n166 ) ? ( n32719 ) : ( n46955 ) ;
assign n46957 =  ( n162 ) ? ( n32718 ) : ( n46956 ) ;
assign n46958 =  ( n32701 ) ? ( VREG_30_8 ) : ( n46957 ) ;
assign n46959 =  ( n3051 ) ? ( n46958 ) : ( VREG_30_8 ) ;
assign n46960 =  ( n3040 ) ? ( n46952 ) : ( n46959 ) ;
assign n46961 =  ( n192 ) ? ( VREG_30_8 ) : ( VREG_30_8 ) ;
assign n46962 =  ( n157 ) ? ( n46960 ) : ( n46961 ) ;
assign n46963 =  ( n6 ) ? ( n46947 ) : ( n46962 ) ;
assign n46964 =  ( n703 ) ? ( n46963 ) : ( VREG_30_8 ) ;
assign n46965 =  ( n148 ) ? ( n33779 ) : ( VREG_30_9 ) ;
assign n46966 =  ( n146 ) ? ( n33778 ) : ( n46965 ) ;
assign n46967 =  ( n144 ) ? ( n33777 ) : ( n46966 ) ;
assign n46968 =  ( n142 ) ? ( n33776 ) : ( n46967 ) ;
assign n46969 =  ( n10 ) ? ( n33775 ) : ( n46968 ) ;
assign n46970 =  ( n148 ) ? ( n34813 ) : ( VREG_30_9 ) ;
assign n46971 =  ( n146 ) ? ( n34812 ) : ( n46970 ) ;
assign n46972 =  ( n144 ) ? ( n34811 ) : ( n46971 ) ;
assign n46973 =  ( n142 ) ? ( n34810 ) : ( n46972 ) ;
assign n46974 =  ( n10 ) ? ( n34809 ) : ( n46973 ) ;
assign n46975 =  ( n34820 ) ? ( VREG_30_9 ) : ( n46969 ) ;
assign n46976 =  ( n34820 ) ? ( VREG_30_9 ) : ( n46974 ) ;
assign n46977 =  ( n3034 ) ? ( n46976 ) : ( VREG_30_9 ) ;
assign n46978 =  ( n2965 ) ? ( n46975 ) : ( n46977 ) ;
assign n46979 =  ( n1930 ) ? ( n46974 ) : ( n46978 ) ;
assign n46980 =  ( n879 ) ? ( n46969 ) : ( n46979 ) ;
assign n46981 =  ( n172 ) ? ( n34831 ) : ( VREG_30_9 ) ;
assign n46982 =  ( n170 ) ? ( n34830 ) : ( n46981 ) ;
assign n46983 =  ( n168 ) ? ( n34829 ) : ( n46982 ) ;
assign n46984 =  ( n166 ) ? ( n34828 ) : ( n46983 ) ;
assign n46985 =  ( n162 ) ? ( n34827 ) : ( n46984 ) ;
assign n46986 =  ( n172 ) ? ( n34841 ) : ( VREG_30_9 ) ;
assign n46987 =  ( n170 ) ? ( n34840 ) : ( n46986 ) ;
assign n46988 =  ( n168 ) ? ( n34839 ) : ( n46987 ) ;
assign n46989 =  ( n166 ) ? ( n34838 ) : ( n46988 ) ;
assign n46990 =  ( n162 ) ? ( n34837 ) : ( n46989 ) ;
assign n46991 =  ( n34820 ) ? ( VREG_30_9 ) : ( n46990 ) ;
assign n46992 =  ( n3051 ) ? ( n46991 ) : ( VREG_30_9 ) ;
assign n46993 =  ( n3040 ) ? ( n46985 ) : ( n46992 ) ;
assign n46994 =  ( n192 ) ? ( VREG_30_9 ) : ( VREG_30_9 ) ;
assign n46995 =  ( n157 ) ? ( n46993 ) : ( n46994 ) ;
assign n46996 =  ( n6 ) ? ( n46980 ) : ( n46995 ) ;
assign n46997 =  ( n703 ) ? ( n46996 ) : ( VREG_30_9 ) ;
assign n46998 =  ( n148 ) ? ( n1924 ) : ( VREG_31_0 ) ;
assign n46999 =  ( n146 ) ? ( n1923 ) : ( n46998 ) ;
assign n47000 =  ( n144 ) ? ( n1922 ) : ( n46999 ) ;
assign n47001 =  ( n142 ) ? ( n1921 ) : ( n47000 ) ;
assign n47002 =  ( n10 ) ? ( n1920 ) : ( n47001 ) ;
assign n47003 =  ( n148 ) ? ( n2959 ) : ( VREG_31_0 ) ;
assign n47004 =  ( n146 ) ? ( n2958 ) : ( n47003 ) ;
assign n47005 =  ( n144 ) ? ( n2957 ) : ( n47004 ) ;
assign n47006 =  ( n142 ) ? ( n2956 ) : ( n47005 ) ;
assign n47007 =  ( n10 ) ? ( n2955 ) : ( n47006 ) ;
assign n47008 =  ( n3032 ) ? ( VREG_31_0 ) : ( n47002 ) ;
assign n47009 =  ( n3032 ) ? ( VREG_31_0 ) : ( n47007 ) ;
assign n47010 =  ( n3034 ) ? ( n47009 ) : ( VREG_31_0 ) ;
assign n47011 =  ( n2965 ) ? ( n47008 ) : ( n47010 ) ;
assign n47012 =  ( n1930 ) ? ( n47007 ) : ( n47011 ) ;
assign n47013 =  ( n879 ) ? ( n47002 ) : ( n47012 ) ;
assign n47014 =  ( n172 ) ? ( n3045 ) : ( VREG_31_0 ) ;
assign n47015 =  ( n170 ) ? ( n3044 ) : ( n47014 ) ;
assign n47016 =  ( n168 ) ? ( n3043 ) : ( n47015 ) ;
assign n47017 =  ( n166 ) ? ( n3042 ) : ( n47016 ) ;
assign n47018 =  ( n162 ) ? ( n3041 ) : ( n47017 ) ;
assign n47019 =  ( n172 ) ? ( n3056 ) : ( VREG_31_0 ) ;
assign n47020 =  ( n170 ) ? ( n3055 ) : ( n47019 ) ;
assign n47021 =  ( n168 ) ? ( n3054 ) : ( n47020 ) ;
assign n47022 =  ( n166 ) ? ( n3053 ) : ( n47021 ) ;
assign n47023 =  ( n162 ) ? ( n3052 ) : ( n47022 ) ;
assign n47024 =  ( n3032 ) ? ( VREG_31_0 ) : ( n47023 ) ;
assign n47025 =  ( n3051 ) ? ( n47024 ) : ( VREG_31_0 ) ;
assign n47026 =  ( n3040 ) ? ( n47018 ) : ( n47025 ) ;
assign n47027 =  ( n192 ) ? ( VREG_31_0 ) : ( VREG_31_0 ) ;
assign n47028 =  ( n157 ) ? ( n47026 ) : ( n47027 ) ;
assign n47029 =  ( n6 ) ? ( n47013 ) : ( n47028 ) ;
assign n47030 =  ( n725 ) ? ( n47029 ) : ( VREG_31_0 ) ;
assign n47031 =  ( n148 ) ? ( n4113 ) : ( VREG_31_1 ) ;
assign n47032 =  ( n146 ) ? ( n4112 ) : ( n47031 ) ;
assign n47033 =  ( n144 ) ? ( n4111 ) : ( n47032 ) ;
assign n47034 =  ( n142 ) ? ( n4110 ) : ( n47033 ) ;
assign n47035 =  ( n10 ) ? ( n4109 ) : ( n47034 ) ;
assign n47036 =  ( n148 ) ? ( n5147 ) : ( VREG_31_1 ) ;
assign n47037 =  ( n146 ) ? ( n5146 ) : ( n47036 ) ;
assign n47038 =  ( n144 ) ? ( n5145 ) : ( n47037 ) ;
assign n47039 =  ( n142 ) ? ( n5144 ) : ( n47038 ) ;
assign n47040 =  ( n10 ) ? ( n5143 ) : ( n47039 ) ;
assign n47041 =  ( n5154 ) ? ( VREG_31_1 ) : ( n47035 ) ;
assign n47042 =  ( n5154 ) ? ( VREG_31_1 ) : ( n47040 ) ;
assign n47043 =  ( n3034 ) ? ( n47042 ) : ( VREG_31_1 ) ;
assign n47044 =  ( n2965 ) ? ( n47041 ) : ( n47043 ) ;
assign n47045 =  ( n1930 ) ? ( n47040 ) : ( n47044 ) ;
assign n47046 =  ( n879 ) ? ( n47035 ) : ( n47045 ) ;
assign n47047 =  ( n172 ) ? ( n5165 ) : ( VREG_31_1 ) ;
assign n47048 =  ( n170 ) ? ( n5164 ) : ( n47047 ) ;
assign n47049 =  ( n168 ) ? ( n5163 ) : ( n47048 ) ;
assign n47050 =  ( n166 ) ? ( n5162 ) : ( n47049 ) ;
assign n47051 =  ( n162 ) ? ( n5161 ) : ( n47050 ) ;
assign n47052 =  ( n172 ) ? ( n5175 ) : ( VREG_31_1 ) ;
assign n47053 =  ( n170 ) ? ( n5174 ) : ( n47052 ) ;
assign n47054 =  ( n168 ) ? ( n5173 ) : ( n47053 ) ;
assign n47055 =  ( n166 ) ? ( n5172 ) : ( n47054 ) ;
assign n47056 =  ( n162 ) ? ( n5171 ) : ( n47055 ) ;
assign n47057 =  ( n5154 ) ? ( VREG_31_1 ) : ( n47056 ) ;
assign n47058 =  ( n3051 ) ? ( n47057 ) : ( VREG_31_1 ) ;
assign n47059 =  ( n3040 ) ? ( n47051 ) : ( n47058 ) ;
assign n47060 =  ( n192 ) ? ( VREG_31_1 ) : ( VREG_31_1 ) ;
assign n47061 =  ( n157 ) ? ( n47059 ) : ( n47060 ) ;
assign n47062 =  ( n6 ) ? ( n47046 ) : ( n47061 ) ;
assign n47063 =  ( n725 ) ? ( n47062 ) : ( VREG_31_1 ) ;
assign n47064 =  ( n148 ) ? ( n6232 ) : ( VREG_31_10 ) ;
assign n47065 =  ( n146 ) ? ( n6231 ) : ( n47064 ) ;
assign n47066 =  ( n144 ) ? ( n6230 ) : ( n47065 ) ;
assign n47067 =  ( n142 ) ? ( n6229 ) : ( n47066 ) ;
assign n47068 =  ( n10 ) ? ( n6228 ) : ( n47067 ) ;
assign n47069 =  ( n148 ) ? ( n7266 ) : ( VREG_31_10 ) ;
assign n47070 =  ( n146 ) ? ( n7265 ) : ( n47069 ) ;
assign n47071 =  ( n144 ) ? ( n7264 ) : ( n47070 ) ;
assign n47072 =  ( n142 ) ? ( n7263 ) : ( n47071 ) ;
assign n47073 =  ( n10 ) ? ( n7262 ) : ( n47072 ) ;
assign n47074 =  ( n7273 ) ? ( VREG_31_10 ) : ( n47068 ) ;
assign n47075 =  ( n7273 ) ? ( VREG_31_10 ) : ( n47073 ) ;
assign n47076 =  ( n3034 ) ? ( n47075 ) : ( VREG_31_10 ) ;
assign n47077 =  ( n2965 ) ? ( n47074 ) : ( n47076 ) ;
assign n47078 =  ( n1930 ) ? ( n47073 ) : ( n47077 ) ;
assign n47079 =  ( n879 ) ? ( n47068 ) : ( n47078 ) ;
assign n47080 =  ( n172 ) ? ( n7284 ) : ( VREG_31_10 ) ;
assign n47081 =  ( n170 ) ? ( n7283 ) : ( n47080 ) ;
assign n47082 =  ( n168 ) ? ( n7282 ) : ( n47081 ) ;
assign n47083 =  ( n166 ) ? ( n7281 ) : ( n47082 ) ;
assign n47084 =  ( n162 ) ? ( n7280 ) : ( n47083 ) ;
assign n47085 =  ( n172 ) ? ( n7294 ) : ( VREG_31_10 ) ;
assign n47086 =  ( n170 ) ? ( n7293 ) : ( n47085 ) ;
assign n47087 =  ( n168 ) ? ( n7292 ) : ( n47086 ) ;
assign n47088 =  ( n166 ) ? ( n7291 ) : ( n47087 ) ;
assign n47089 =  ( n162 ) ? ( n7290 ) : ( n47088 ) ;
assign n47090 =  ( n7273 ) ? ( VREG_31_10 ) : ( n47089 ) ;
assign n47091 =  ( n3051 ) ? ( n47090 ) : ( VREG_31_10 ) ;
assign n47092 =  ( n3040 ) ? ( n47084 ) : ( n47091 ) ;
assign n47093 =  ( n192 ) ? ( VREG_31_10 ) : ( VREG_31_10 ) ;
assign n47094 =  ( n157 ) ? ( n47092 ) : ( n47093 ) ;
assign n47095 =  ( n6 ) ? ( n47079 ) : ( n47094 ) ;
assign n47096 =  ( n725 ) ? ( n47095 ) : ( VREG_31_10 ) ;
assign n47097 =  ( n148 ) ? ( n8351 ) : ( VREG_31_11 ) ;
assign n47098 =  ( n146 ) ? ( n8350 ) : ( n47097 ) ;
assign n47099 =  ( n144 ) ? ( n8349 ) : ( n47098 ) ;
assign n47100 =  ( n142 ) ? ( n8348 ) : ( n47099 ) ;
assign n47101 =  ( n10 ) ? ( n8347 ) : ( n47100 ) ;
assign n47102 =  ( n148 ) ? ( n9385 ) : ( VREG_31_11 ) ;
assign n47103 =  ( n146 ) ? ( n9384 ) : ( n47102 ) ;
assign n47104 =  ( n144 ) ? ( n9383 ) : ( n47103 ) ;
assign n47105 =  ( n142 ) ? ( n9382 ) : ( n47104 ) ;
assign n47106 =  ( n10 ) ? ( n9381 ) : ( n47105 ) ;
assign n47107 =  ( n9392 ) ? ( VREG_31_11 ) : ( n47101 ) ;
assign n47108 =  ( n9392 ) ? ( VREG_31_11 ) : ( n47106 ) ;
assign n47109 =  ( n3034 ) ? ( n47108 ) : ( VREG_31_11 ) ;
assign n47110 =  ( n2965 ) ? ( n47107 ) : ( n47109 ) ;
assign n47111 =  ( n1930 ) ? ( n47106 ) : ( n47110 ) ;
assign n47112 =  ( n879 ) ? ( n47101 ) : ( n47111 ) ;
assign n47113 =  ( n172 ) ? ( n9403 ) : ( VREG_31_11 ) ;
assign n47114 =  ( n170 ) ? ( n9402 ) : ( n47113 ) ;
assign n47115 =  ( n168 ) ? ( n9401 ) : ( n47114 ) ;
assign n47116 =  ( n166 ) ? ( n9400 ) : ( n47115 ) ;
assign n47117 =  ( n162 ) ? ( n9399 ) : ( n47116 ) ;
assign n47118 =  ( n172 ) ? ( n9413 ) : ( VREG_31_11 ) ;
assign n47119 =  ( n170 ) ? ( n9412 ) : ( n47118 ) ;
assign n47120 =  ( n168 ) ? ( n9411 ) : ( n47119 ) ;
assign n47121 =  ( n166 ) ? ( n9410 ) : ( n47120 ) ;
assign n47122 =  ( n162 ) ? ( n9409 ) : ( n47121 ) ;
assign n47123 =  ( n9392 ) ? ( VREG_31_11 ) : ( n47122 ) ;
assign n47124 =  ( n3051 ) ? ( n47123 ) : ( VREG_31_11 ) ;
assign n47125 =  ( n3040 ) ? ( n47117 ) : ( n47124 ) ;
assign n47126 =  ( n192 ) ? ( VREG_31_11 ) : ( VREG_31_11 ) ;
assign n47127 =  ( n157 ) ? ( n47125 ) : ( n47126 ) ;
assign n47128 =  ( n6 ) ? ( n47112 ) : ( n47127 ) ;
assign n47129 =  ( n725 ) ? ( n47128 ) : ( VREG_31_11 ) ;
assign n47130 =  ( n148 ) ? ( n10470 ) : ( VREG_31_12 ) ;
assign n47131 =  ( n146 ) ? ( n10469 ) : ( n47130 ) ;
assign n47132 =  ( n144 ) ? ( n10468 ) : ( n47131 ) ;
assign n47133 =  ( n142 ) ? ( n10467 ) : ( n47132 ) ;
assign n47134 =  ( n10 ) ? ( n10466 ) : ( n47133 ) ;
assign n47135 =  ( n148 ) ? ( n11504 ) : ( VREG_31_12 ) ;
assign n47136 =  ( n146 ) ? ( n11503 ) : ( n47135 ) ;
assign n47137 =  ( n144 ) ? ( n11502 ) : ( n47136 ) ;
assign n47138 =  ( n142 ) ? ( n11501 ) : ( n47137 ) ;
assign n47139 =  ( n10 ) ? ( n11500 ) : ( n47138 ) ;
assign n47140 =  ( n11511 ) ? ( VREG_31_12 ) : ( n47134 ) ;
assign n47141 =  ( n11511 ) ? ( VREG_31_12 ) : ( n47139 ) ;
assign n47142 =  ( n3034 ) ? ( n47141 ) : ( VREG_31_12 ) ;
assign n47143 =  ( n2965 ) ? ( n47140 ) : ( n47142 ) ;
assign n47144 =  ( n1930 ) ? ( n47139 ) : ( n47143 ) ;
assign n47145 =  ( n879 ) ? ( n47134 ) : ( n47144 ) ;
assign n47146 =  ( n172 ) ? ( n11522 ) : ( VREG_31_12 ) ;
assign n47147 =  ( n170 ) ? ( n11521 ) : ( n47146 ) ;
assign n47148 =  ( n168 ) ? ( n11520 ) : ( n47147 ) ;
assign n47149 =  ( n166 ) ? ( n11519 ) : ( n47148 ) ;
assign n47150 =  ( n162 ) ? ( n11518 ) : ( n47149 ) ;
assign n47151 =  ( n172 ) ? ( n11532 ) : ( VREG_31_12 ) ;
assign n47152 =  ( n170 ) ? ( n11531 ) : ( n47151 ) ;
assign n47153 =  ( n168 ) ? ( n11530 ) : ( n47152 ) ;
assign n47154 =  ( n166 ) ? ( n11529 ) : ( n47153 ) ;
assign n47155 =  ( n162 ) ? ( n11528 ) : ( n47154 ) ;
assign n47156 =  ( n11511 ) ? ( VREG_31_12 ) : ( n47155 ) ;
assign n47157 =  ( n3051 ) ? ( n47156 ) : ( VREG_31_12 ) ;
assign n47158 =  ( n3040 ) ? ( n47150 ) : ( n47157 ) ;
assign n47159 =  ( n192 ) ? ( VREG_31_12 ) : ( VREG_31_12 ) ;
assign n47160 =  ( n157 ) ? ( n47158 ) : ( n47159 ) ;
assign n47161 =  ( n6 ) ? ( n47145 ) : ( n47160 ) ;
assign n47162 =  ( n725 ) ? ( n47161 ) : ( VREG_31_12 ) ;
assign n47163 =  ( n148 ) ? ( n12589 ) : ( VREG_31_13 ) ;
assign n47164 =  ( n146 ) ? ( n12588 ) : ( n47163 ) ;
assign n47165 =  ( n144 ) ? ( n12587 ) : ( n47164 ) ;
assign n47166 =  ( n142 ) ? ( n12586 ) : ( n47165 ) ;
assign n47167 =  ( n10 ) ? ( n12585 ) : ( n47166 ) ;
assign n47168 =  ( n148 ) ? ( n13623 ) : ( VREG_31_13 ) ;
assign n47169 =  ( n146 ) ? ( n13622 ) : ( n47168 ) ;
assign n47170 =  ( n144 ) ? ( n13621 ) : ( n47169 ) ;
assign n47171 =  ( n142 ) ? ( n13620 ) : ( n47170 ) ;
assign n47172 =  ( n10 ) ? ( n13619 ) : ( n47171 ) ;
assign n47173 =  ( n13630 ) ? ( VREG_31_13 ) : ( n47167 ) ;
assign n47174 =  ( n13630 ) ? ( VREG_31_13 ) : ( n47172 ) ;
assign n47175 =  ( n3034 ) ? ( n47174 ) : ( VREG_31_13 ) ;
assign n47176 =  ( n2965 ) ? ( n47173 ) : ( n47175 ) ;
assign n47177 =  ( n1930 ) ? ( n47172 ) : ( n47176 ) ;
assign n47178 =  ( n879 ) ? ( n47167 ) : ( n47177 ) ;
assign n47179 =  ( n172 ) ? ( n13641 ) : ( VREG_31_13 ) ;
assign n47180 =  ( n170 ) ? ( n13640 ) : ( n47179 ) ;
assign n47181 =  ( n168 ) ? ( n13639 ) : ( n47180 ) ;
assign n47182 =  ( n166 ) ? ( n13638 ) : ( n47181 ) ;
assign n47183 =  ( n162 ) ? ( n13637 ) : ( n47182 ) ;
assign n47184 =  ( n172 ) ? ( n13651 ) : ( VREG_31_13 ) ;
assign n47185 =  ( n170 ) ? ( n13650 ) : ( n47184 ) ;
assign n47186 =  ( n168 ) ? ( n13649 ) : ( n47185 ) ;
assign n47187 =  ( n166 ) ? ( n13648 ) : ( n47186 ) ;
assign n47188 =  ( n162 ) ? ( n13647 ) : ( n47187 ) ;
assign n47189 =  ( n13630 ) ? ( VREG_31_13 ) : ( n47188 ) ;
assign n47190 =  ( n3051 ) ? ( n47189 ) : ( VREG_31_13 ) ;
assign n47191 =  ( n3040 ) ? ( n47183 ) : ( n47190 ) ;
assign n47192 =  ( n192 ) ? ( VREG_31_13 ) : ( VREG_31_13 ) ;
assign n47193 =  ( n157 ) ? ( n47191 ) : ( n47192 ) ;
assign n47194 =  ( n6 ) ? ( n47178 ) : ( n47193 ) ;
assign n47195 =  ( n725 ) ? ( n47194 ) : ( VREG_31_13 ) ;
assign n47196 =  ( n148 ) ? ( n14708 ) : ( VREG_31_14 ) ;
assign n47197 =  ( n146 ) ? ( n14707 ) : ( n47196 ) ;
assign n47198 =  ( n144 ) ? ( n14706 ) : ( n47197 ) ;
assign n47199 =  ( n142 ) ? ( n14705 ) : ( n47198 ) ;
assign n47200 =  ( n10 ) ? ( n14704 ) : ( n47199 ) ;
assign n47201 =  ( n148 ) ? ( n15742 ) : ( VREG_31_14 ) ;
assign n47202 =  ( n146 ) ? ( n15741 ) : ( n47201 ) ;
assign n47203 =  ( n144 ) ? ( n15740 ) : ( n47202 ) ;
assign n47204 =  ( n142 ) ? ( n15739 ) : ( n47203 ) ;
assign n47205 =  ( n10 ) ? ( n15738 ) : ( n47204 ) ;
assign n47206 =  ( n15749 ) ? ( VREG_31_14 ) : ( n47200 ) ;
assign n47207 =  ( n15749 ) ? ( VREG_31_14 ) : ( n47205 ) ;
assign n47208 =  ( n3034 ) ? ( n47207 ) : ( VREG_31_14 ) ;
assign n47209 =  ( n2965 ) ? ( n47206 ) : ( n47208 ) ;
assign n47210 =  ( n1930 ) ? ( n47205 ) : ( n47209 ) ;
assign n47211 =  ( n879 ) ? ( n47200 ) : ( n47210 ) ;
assign n47212 =  ( n172 ) ? ( n15760 ) : ( VREG_31_14 ) ;
assign n47213 =  ( n170 ) ? ( n15759 ) : ( n47212 ) ;
assign n47214 =  ( n168 ) ? ( n15758 ) : ( n47213 ) ;
assign n47215 =  ( n166 ) ? ( n15757 ) : ( n47214 ) ;
assign n47216 =  ( n162 ) ? ( n15756 ) : ( n47215 ) ;
assign n47217 =  ( n172 ) ? ( n15770 ) : ( VREG_31_14 ) ;
assign n47218 =  ( n170 ) ? ( n15769 ) : ( n47217 ) ;
assign n47219 =  ( n168 ) ? ( n15768 ) : ( n47218 ) ;
assign n47220 =  ( n166 ) ? ( n15767 ) : ( n47219 ) ;
assign n47221 =  ( n162 ) ? ( n15766 ) : ( n47220 ) ;
assign n47222 =  ( n15749 ) ? ( VREG_31_14 ) : ( n47221 ) ;
assign n47223 =  ( n3051 ) ? ( n47222 ) : ( VREG_31_14 ) ;
assign n47224 =  ( n3040 ) ? ( n47216 ) : ( n47223 ) ;
assign n47225 =  ( n192 ) ? ( VREG_31_14 ) : ( VREG_31_14 ) ;
assign n47226 =  ( n157 ) ? ( n47224 ) : ( n47225 ) ;
assign n47227 =  ( n6 ) ? ( n47211 ) : ( n47226 ) ;
assign n47228 =  ( n725 ) ? ( n47227 ) : ( VREG_31_14 ) ;
assign n47229 =  ( n148 ) ? ( n16827 ) : ( VREG_31_15 ) ;
assign n47230 =  ( n146 ) ? ( n16826 ) : ( n47229 ) ;
assign n47231 =  ( n144 ) ? ( n16825 ) : ( n47230 ) ;
assign n47232 =  ( n142 ) ? ( n16824 ) : ( n47231 ) ;
assign n47233 =  ( n10 ) ? ( n16823 ) : ( n47232 ) ;
assign n47234 =  ( n148 ) ? ( n17861 ) : ( VREG_31_15 ) ;
assign n47235 =  ( n146 ) ? ( n17860 ) : ( n47234 ) ;
assign n47236 =  ( n144 ) ? ( n17859 ) : ( n47235 ) ;
assign n47237 =  ( n142 ) ? ( n17858 ) : ( n47236 ) ;
assign n47238 =  ( n10 ) ? ( n17857 ) : ( n47237 ) ;
assign n47239 =  ( n17868 ) ? ( VREG_31_15 ) : ( n47233 ) ;
assign n47240 =  ( n17868 ) ? ( VREG_31_15 ) : ( n47238 ) ;
assign n47241 =  ( n3034 ) ? ( n47240 ) : ( VREG_31_15 ) ;
assign n47242 =  ( n2965 ) ? ( n47239 ) : ( n47241 ) ;
assign n47243 =  ( n1930 ) ? ( n47238 ) : ( n47242 ) ;
assign n47244 =  ( n879 ) ? ( n47233 ) : ( n47243 ) ;
assign n47245 =  ( n172 ) ? ( n17879 ) : ( VREG_31_15 ) ;
assign n47246 =  ( n170 ) ? ( n17878 ) : ( n47245 ) ;
assign n47247 =  ( n168 ) ? ( n17877 ) : ( n47246 ) ;
assign n47248 =  ( n166 ) ? ( n17876 ) : ( n47247 ) ;
assign n47249 =  ( n162 ) ? ( n17875 ) : ( n47248 ) ;
assign n47250 =  ( n172 ) ? ( n17889 ) : ( VREG_31_15 ) ;
assign n47251 =  ( n170 ) ? ( n17888 ) : ( n47250 ) ;
assign n47252 =  ( n168 ) ? ( n17887 ) : ( n47251 ) ;
assign n47253 =  ( n166 ) ? ( n17886 ) : ( n47252 ) ;
assign n47254 =  ( n162 ) ? ( n17885 ) : ( n47253 ) ;
assign n47255 =  ( n17868 ) ? ( VREG_31_15 ) : ( n47254 ) ;
assign n47256 =  ( n3051 ) ? ( n47255 ) : ( VREG_31_15 ) ;
assign n47257 =  ( n3040 ) ? ( n47249 ) : ( n47256 ) ;
assign n47258 =  ( n192 ) ? ( VREG_31_15 ) : ( VREG_31_15 ) ;
assign n47259 =  ( n157 ) ? ( n47257 ) : ( n47258 ) ;
assign n47260 =  ( n6 ) ? ( n47244 ) : ( n47259 ) ;
assign n47261 =  ( n725 ) ? ( n47260 ) : ( VREG_31_15 ) ;
assign n47262 =  ( n148 ) ? ( n18946 ) : ( VREG_31_2 ) ;
assign n47263 =  ( n146 ) ? ( n18945 ) : ( n47262 ) ;
assign n47264 =  ( n144 ) ? ( n18944 ) : ( n47263 ) ;
assign n47265 =  ( n142 ) ? ( n18943 ) : ( n47264 ) ;
assign n47266 =  ( n10 ) ? ( n18942 ) : ( n47265 ) ;
assign n47267 =  ( n148 ) ? ( n19980 ) : ( VREG_31_2 ) ;
assign n47268 =  ( n146 ) ? ( n19979 ) : ( n47267 ) ;
assign n47269 =  ( n144 ) ? ( n19978 ) : ( n47268 ) ;
assign n47270 =  ( n142 ) ? ( n19977 ) : ( n47269 ) ;
assign n47271 =  ( n10 ) ? ( n19976 ) : ( n47270 ) ;
assign n47272 =  ( n19987 ) ? ( VREG_31_2 ) : ( n47266 ) ;
assign n47273 =  ( n19987 ) ? ( VREG_31_2 ) : ( n47271 ) ;
assign n47274 =  ( n3034 ) ? ( n47273 ) : ( VREG_31_2 ) ;
assign n47275 =  ( n2965 ) ? ( n47272 ) : ( n47274 ) ;
assign n47276 =  ( n1930 ) ? ( n47271 ) : ( n47275 ) ;
assign n47277 =  ( n879 ) ? ( n47266 ) : ( n47276 ) ;
assign n47278 =  ( n172 ) ? ( n19998 ) : ( VREG_31_2 ) ;
assign n47279 =  ( n170 ) ? ( n19997 ) : ( n47278 ) ;
assign n47280 =  ( n168 ) ? ( n19996 ) : ( n47279 ) ;
assign n47281 =  ( n166 ) ? ( n19995 ) : ( n47280 ) ;
assign n47282 =  ( n162 ) ? ( n19994 ) : ( n47281 ) ;
assign n47283 =  ( n172 ) ? ( n20008 ) : ( VREG_31_2 ) ;
assign n47284 =  ( n170 ) ? ( n20007 ) : ( n47283 ) ;
assign n47285 =  ( n168 ) ? ( n20006 ) : ( n47284 ) ;
assign n47286 =  ( n166 ) ? ( n20005 ) : ( n47285 ) ;
assign n47287 =  ( n162 ) ? ( n20004 ) : ( n47286 ) ;
assign n47288 =  ( n19987 ) ? ( VREG_31_2 ) : ( n47287 ) ;
assign n47289 =  ( n3051 ) ? ( n47288 ) : ( VREG_31_2 ) ;
assign n47290 =  ( n3040 ) ? ( n47282 ) : ( n47289 ) ;
assign n47291 =  ( n192 ) ? ( VREG_31_2 ) : ( VREG_31_2 ) ;
assign n47292 =  ( n157 ) ? ( n47290 ) : ( n47291 ) ;
assign n47293 =  ( n6 ) ? ( n47277 ) : ( n47292 ) ;
assign n47294 =  ( n725 ) ? ( n47293 ) : ( VREG_31_2 ) ;
assign n47295 =  ( n148 ) ? ( n21065 ) : ( VREG_31_3 ) ;
assign n47296 =  ( n146 ) ? ( n21064 ) : ( n47295 ) ;
assign n47297 =  ( n144 ) ? ( n21063 ) : ( n47296 ) ;
assign n47298 =  ( n142 ) ? ( n21062 ) : ( n47297 ) ;
assign n47299 =  ( n10 ) ? ( n21061 ) : ( n47298 ) ;
assign n47300 =  ( n148 ) ? ( n22099 ) : ( VREG_31_3 ) ;
assign n47301 =  ( n146 ) ? ( n22098 ) : ( n47300 ) ;
assign n47302 =  ( n144 ) ? ( n22097 ) : ( n47301 ) ;
assign n47303 =  ( n142 ) ? ( n22096 ) : ( n47302 ) ;
assign n47304 =  ( n10 ) ? ( n22095 ) : ( n47303 ) ;
assign n47305 =  ( n22106 ) ? ( VREG_31_3 ) : ( n47299 ) ;
assign n47306 =  ( n22106 ) ? ( VREG_31_3 ) : ( n47304 ) ;
assign n47307 =  ( n3034 ) ? ( n47306 ) : ( VREG_31_3 ) ;
assign n47308 =  ( n2965 ) ? ( n47305 ) : ( n47307 ) ;
assign n47309 =  ( n1930 ) ? ( n47304 ) : ( n47308 ) ;
assign n47310 =  ( n879 ) ? ( n47299 ) : ( n47309 ) ;
assign n47311 =  ( n172 ) ? ( n22117 ) : ( VREG_31_3 ) ;
assign n47312 =  ( n170 ) ? ( n22116 ) : ( n47311 ) ;
assign n47313 =  ( n168 ) ? ( n22115 ) : ( n47312 ) ;
assign n47314 =  ( n166 ) ? ( n22114 ) : ( n47313 ) ;
assign n47315 =  ( n162 ) ? ( n22113 ) : ( n47314 ) ;
assign n47316 =  ( n172 ) ? ( n22127 ) : ( VREG_31_3 ) ;
assign n47317 =  ( n170 ) ? ( n22126 ) : ( n47316 ) ;
assign n47318 =  ( n168 ) ? ( n22125 ) : ( n47317 ) ;
assign n47319 =  ( n166 ) ? ( n22124 ) : ( n47318 ) ;
assign n47320 =  ( n162 ) ? ( n22123 ) : ( n47319 ) ;
assign n47321 =  ( n22106 ) ? ( VREG_31_3 ) : ( n47320 ) ;
assign n47322 =  ( n3051 ) ? ( n47321 ) : ( VREG_31_3 ) ;
assign n47323 =  ( n3040 ) ? ( n47315 ) : ( n47322 ) ;
assign n47324 =  ( n192 ) ? ( VREG_31_3 ) : ( VREG_31_3 ) ;
assign n47325 =  ( n157 ) ? ( n47323 ) : ( n47324 ) ;
assign n47326 =  ( n6 ) ? ( n47310 ) : ( n47325 ) ;
assign n47327 =  ( n725 ) ? ( n47326 ) : ( VREG_31_3 ) ;
assign n47328 =  ( n148 ) ? ( n23184 ) : ( VREG_31_4 ) ;
assign n47329 =  ( n146 ) ? ( n23183 ) : ( n47328 ) ;
assign n47330 =  ( n144 ) ? ( n23182 ) : ( n47329 ) ;
assign n47331 =  ( n142 ) ? ( n23181 ) : ( n47330 ) ;
assign n47332 =  ( n10 ) ? ( n23180 ) : ( n47331 ) ;
assign n47333 =  ( n148 ) ? ( n24218 ) : ( VREG_31_4 ) ;
assign n47334 =  ( n146 ) ? ( n24217 ) : ( n47333 ) ;
assign n47335 =  ( n144 ) ? ( n24216 ) : ( n47334 ) ;
assign n47336 =  ( n142 ) ? ( n24215 ) : ( n47335 ) ;
assign n47337 =  ( n10 ) ? ( n24214 ) : ( n47336 ) ;
assign n47338 =  ( n24225 ) ? ( VREG_31_4 ) : ( n47332 ) ;
assign n47339 =  ( n24225 ) ? ( VREG_31_4 ) : ( n47337 ) ;
assign n47340 =  ( n3034 ) ? ( n47339 ) : ( VREG_31_4 ) ;
assign n47341 =  ( n2965 ) ? ( n47338 ) : ( n47340 ) ;
assign n47342 =  ( n1930 ) ? ( n47337 ) : ( n47341 ) ;
assign n47343 =  ( n879 ) ? ( n47332 ) : ( n47342 ) ;
assign n47344 =  ( n172 ) ? ( n24236 ) : ( VREG_31_4 ) ;
assign n47345 =  ( n170 ) ? ( n24235 ) : ( n47344 ) ;
assign n47346 =  ( n168 ) ? ( n24234 ) : ( n47345 ) ;
assign n47347 =  ( n166 ) ? ( n24233 ) : ( n47346 ) ;
assign n47348 =  ( n162 ) ? ( n24232 ) : ( n47347 ) ;
assign n47349 =  ( n172 ) ? ( n24246 ) : ( VREG_31_4 ) ;
assign n47350 =  ( n170 ) ? ( n24245 ) : ( n47349 ) ;
assign n47351 =  ( n168 ) ? ( n24244 ) : ( n47350 ) ;
assign n47352 =  ( n166 ) ? ( n24243 ) : ( n47351 ) ;
assign n47353 =  ( n162 ) ? ( n24242 ) : ( n47352 ) ;
assign n47354 =  ( n24225 ) ? ( VREG_31_4 ) : ( n47353 ) ;
assign n47355 =  ( n3051 ) ? ( n47354 ) : ( VREG_31_4 ) ;
assign n47356 =  ( n3040 ) ? ( n47348 ) : ( n47355 ) ;
assign n47357 =  ( n192 ) ? ( VREG_31_4 ) : ( VREG_31_4 ) ;
assign n47358 =  ( n157 ) ? ( n47356 ) : ( n47357 ) ;
assign n47359 =  ( n6 ) ? ( n47343 ) : ( n47358 ) ;
assign n47360 =  ( n725 ) ? ( n47359 ) : ( VREG_31_4 ) ;
assign n47361 =  ( n148 ) ? ( n25303 ) : ( VREG_31_5 ) ;
assign n47362 =  ( n146 ) ? ( n25302 ) : ( n47361 ) ;
assign n47363 =  ( n144 ) ? ( n25301 ) : ( n47362 ) ;
assign n47364 =  ( n142 ) ? ( n25300 ) : ( n47363 ) ;
assign n47365 =  ( n10 ) ? ( n25299 ) : ( n47364 ) ;
assign n47366 =  ( n148 ) ? ( n26337 ) : ( VREG_31_5 ) ;
assign n47367 =  ( n146 ) ? ( n26336 ) : ( n47366 ) ;
assign n47368 =  ( n144 ) ? ( n26335 ) : ( n47367 ) ;
assign n47369 =  ( n142 ) ? ( n26334 ) : ( n47368 ) ;
assign n47370 =  ( n10 ) ? ( n26333 ) : ( n47369 ) ;
assign n47371 =  ( n26344 ) ? ( VREG_31_5 ) : ( n47365 ) ;
assign n47372 =  ( n26344 ) ? ( VREG_31_5 ) : ( n47370 ) ;
assign n47373 =  ( n3034 ) ? ( n47372 ) : ( VREG_31_5 ) ;
assign n47374 =  ( n2965 ) ? ( n47371 ) : ( n47373 ) ;
assign n47375 =  ( n1930 ) ? ( n47370 ) : ( n47374 ) ;
assign n47376 =  ( n879 ) ? ( n47365 ) : ( n47375 ) ;
assign n47377 =  ( n172 ) ? ( n26355 ) : ( VREG_31_5 ) ;
assign n47378 =  ( n170 ) ? ( n26354 ) : ( n47377 ) ;
assign n47379 =  ( n168 ) ? ( n26353 ) : ( n47378 ) ;
assign n47380 =  ( n166 ) ? ( n26352 ) : ( n47379 ) ;
assign n47381 =  ( n162 ) ? ( n26351 ) : ( n47380 ) ;
assign n47382 =  ( n172 ) ? ( n26365 ) : ( VREG_31_5 ) ;
assign n47383 =  ( n170 ) ? ( n26364 ) : ( n47382 ) ;
assign n47384 =  ( n168 ) ? ( n26363 ) : ( n47383 ) ;
assign n47385 =  ( n166 ) ? ( n26362 ) : ( n47384 ) ;
assign n47386 =  ( n162 ) ? ( n26361 ) : ( n47385 ) ;
assign n47387 =  ( n26344 ) ? ( VREG_31_5 ) : ( n47386 ) ;
assign n47388 =  ( n3051 ) ? ( n47387 ) : ( VREG_31_5 ) ;
assign n47389 =  ( n3040 ) ? ( n47381 ) : ( n47388 ) ;
assign n47390 =  ( n192 ) ? ( VREG_31_5 ) : ( VREG_31_5 ) ;
assign n47391 =  ( n157 ) ? ( n47389 ) : ( n47390 ) ;
assign n47392 =  ( n6 ) ? ( n47376 ) : ( n47391 ) ;
assign n47393 =  ( n725 ) ? ( n47392 ) : ( VREG_31_5 ) ;
assign n47394 =  ( n148 ) ? ( n27422 ) : ( VREG_31_6 ) ;
assign n47395 =  ( n146 ) ? ( n27421 ) : ( n47394 ) ;
assign n47396 =  ( n144 ) ? ( n27420 ) : ( n47395 ) ;
assign n47397 =  ( n142 ) ? ( n27419 ) : ( n47396 ) ;
assign n47398 =  ( n10 ) ? ( n27418 ) : ( n47397 ) ;
assign n47399 =  ( n148 ) ? ( n28456 ) : ( VREG_31_6 ) ;
assign n47400 =  ( n146 ) ? ( n28455 ) : ( n47399 ) ;
assign n47401 =  ( n144 ) ? ( n28454 ) : ( n47400 ) ;
assign n47402 =  ( n142 ) ? ( n28453 ) : ( n47401 ) ;
assign n47403 =  ( n10 ) ? ( n28452 ) : ( n47402 ) ;
assign n47404 =  ( n28463 ) ? ( VREG_31_6 ) : ( n47398 ) ;
assign n47405 =  ( n28463 ) ? ( VREG_31_6 ) : ( n47403 ) ;
assign n47406 =  ( n3034 ) ? ( n47405 ) : ( VREG_31_6 ) ;
assign n47407 =  ( n2965 ) ? ( n47404 ) : ( n47406 ) ;
assign n47408 =  ( n1930 ) ? ( n47403 ) : ( n47407 ) ;
assign n47409 =  ( n879 ) ? ( n47398 ) : ( n47408 ) ;
assign n47410 =  ( n172 ) ? ( n28474 ) : ( VREG_31_6 ) ;
assign n47411 =  ( n170 ) ? ( n28473 ) : ( n47410 ) ;
assign n47412 =  ( n168 ) ? ( n28472 ) : ( n47411 ) ;
assign n47413 =  ( n166 ) ? ( n28471 ) : ( n47412 ) ;
assign n47414 =  ( n162 ) ? ( n28470 ) : ( n47413 ) ;
assign n47415 =  ( n172 ) ? ( n28484 ) : ( VREG_31_6 ) ;
assign n47416 =  ( n170 ) ? ( n28483 ) : ( n47415 ) ;
assign n47417 =  ( n168 ) ? ( n28482 ) : ( n47416 ) ;
assign n47418 =  ( n166 ) ? ( n28481 ) : ( n47417 ) ;
assign n47419 =  ( n162 ) ? ( n28480 ) : ( n47418 ) ;
assign n47420 =  ( n28463 ) ? ( VREG_31_6 ) : ( n47419 ) ;
assign n47421 =  ( n3051 ) ? ( n47420 ) : ( VREG_31_6 ) ;
assign n47422 =  ( n3040 ) ? ( n47414 ) : ( n47421 ) ;
assign n47423 =  ( n192 ) ? ( VREG_31_6 ) : ( VREG_31_6 ) ;
assign n47424 =  ( n157 ) ? ( n47422 ) : ( n47423 ) ;
assign n47425 =  ( n6 ) ? ( n47409 ) : ( n47424 ) ;
assign n47426 =  ( n725 ) ? ( n47425 ) : ( VREG_31_6 ) ;
assign n47427 =  ( n148 ) ? ( n29541 ) : ( VREG_31_7 ) ;
assign n47428 =  ( n146 ) ? ( n29540 ) : ( n47427 ) ;
assign n47429 =  ( n144 ) ? ( n29539 ) : ( n47428 ) ;
assign n47430 =  ( n142 ) ? ( n29538 ) : ( n47429 ) ;
assign n47431 =  ( n10 ) ? ( n29537 ) : ( n47430 ) ;
assign n47432 =  ( n148 ) ? ( n30575 ) : ( VREG_31_7 ) ;
assign n47433 =  ( n146 ) ? ( n30574 ) : ( n47432 ) ;
assign n47434 =  ( n144 ) ? ( n30573 ) : ( n47433 ) ;
assign n47435 =  ( n142 ) ? ( n30572 ) : ( n47434 ) ;
assign n47436 =  ( n10 ) ? ( n30571 ) : ( n47435 ) ;
assign n47437 =  ( n30582 ) ? ( VREG_31_7 ) : ( n47431 ) ;
assign n47438 =  ( n30582 ) ? ( VREG_31_7 ) : ( n47436 ) ;
assign n47439 =  ( n3034 ) ? ( n47438 ) : ( VREG_31_7 ) ;
assign n47440 =  ( n2965 ) ? ( n47437 ) : ( n47439 ) ;
assign n47441 =  ( n1930 ) ? ( n47436 ) : ( n47440 ) ;
assign n47442 =  ( n879 ) ? ( n47431 ) : ( n47441 ) ;
assign n47443 =  ( n172 ) ? ( n30593 ) : ( VREG_31_7 ) ;
assign n47444 =  ( n170 ) ? ( n30592 ) : ( n47443 ) ;
assign n47445 =  ( n168 ) ? ( n30591 ) : ( n47444 ) ;
assign n47446 =  ( n166 ) ? ( n30590 ) : ( n47445 ) ;
assign n47447 =  ( n162 ) ? ( n30589 ) : ( n47446 ) ;
assign n47448 =  ( n172 ) ? ( n30603 ) : ( VREG_31_7 ) ;
assign n47449 =  ( n170 ) ? ( n30602 ) : ( n47448 ) ;
assign n47450 =  ( n168 ) ? ( n30601 ) : ( n47449 ) ;
assign n47451 =  ( n166 ) ? ( n30600 ) : ( n47450 ) ;
assign n47452 =  ( n162 ) ? ( n30599 ) : ( n47451 ) ;
assign n47453 =  ( n30582 ) ? ( VREG_31_7 ) : ( n47452 ) ;
assign n47454 =  ( n3051 ) ? ( n47453 ) : ( VREG_31_7 ) ;
assign n47455 =  ( n3040 ) ? ( n47447 ) : ( n47454 ) ;
assign n47456 =  ( n192 ) ? ( VREG_31_7 ) : ( VREG_31_7 ) ;
assign n47457 =  ( n157 ) ? ( n47455 ) : ( n47456 ) ;
assign n47458 =  ( n6 ) ? ( n47442 ) : ( n47457 ) ;
assign n47459 =  ( n725 ) ? ( n47458 ) : ( VREG_31_7 ) ;
assign n47460 =  ( n148 ) ? ( n31660 ) : ( VREG_31_8 ) ;
assign n47461 =  ( n146 ) ? ( n31659 ) : ( n47460 ) ;
assign n47462 =  ( n144 ) ? ( n31658 ) : ( n47461 ) ;
assign n47463 =  ( n142 ) ? ( n31657 ) : ( n47462 ) ;
assign n47464 =  ( n10 ) ? ( n31656 ) : ( n47463 ) ;
assign n47465 =  ( n148 ) ? ( n32694 ) : ( VREG_31_8 ) ;
assign n47466 =  ( n146 ) ? ( n32693 ) : ( n47465 ) ;
assign n47467 =  ( n144 ) ? ( n32692 ) : ( n47466 ) ;
assign n47468 =  ( n142 ) ? ( n32691 ) : ( n47467 ) ;
assign n47469 =  ( n10 ) ? ( n32690 ) : ( n47468 ) ;
assign n47470 =  ( n32701 ) ? ( VREG_31_8 ) : ( n47464 ) ;
assign n47471 =  ( n32701 ) ? ( VREG_31_8 ) : ( n47469 ) ;
assign n47472 =  ( n3034 ) ? ( n47471 ) : ( VREG_31_8 ) ;
assign n47473 =  ( n2965 ) ? ( n47470 ) : ( n47472 ) ;
assign n47474 =  ( n1930 ) ? ( n47469 ) : ( n47473 ) ;
assign n47475 =  ( n879 ) ? ( n47464 ) : ( n47474 ) ;
assign n47476 =  ( n172 ) ? ( n32712 ) : ( VREG_31_8 ) ;
assign n47477 =  ( n170 ) ? ( n32711 ) : ( n47476 ) ;
assign n47478 =  ( n168 ) ? ( n32710 ) : ( n47477 ) ;
assign n47479 =  ( n166 ) ? ( n32709 ) : ( n47478 ) ;
assign n47480 =  ( n162 ) ? ( n32708 ) : ( n47479 ) ;
assign n47481 =  ( n172 ) ? ( n32722 ) : ( VREG_31_8 ) ;
assign n47482 =  ( n170 ) ? ( n32721 ) : ( n47481 ) ;
assign n47483 =  ( n168 ) ? ( n32720 ) : ( n47482 ) ;
assign n47484 =  ( n166 ) ? ( n32719 ) : ( n47483 ) ;
assign n47485 =  ( n162 ) ? ( n32718 ) : ( n47484 ) ;
assign n47486 =  ( n32701 ) ? ( VREG_31_8 ) : ( n47485 ) ;
assign n47487 =  ( n3051 ) ? ( n47486 ) : ( VREG_31_8 ) ;
assign n47488 =  ( n3040 ) ? ( n47480 ) : ( n47487 ) ;
assign n47489 =  ( n192 ) ? ( VREG_31_8 ) : ( VREG_31_8 ) ;
assign n47490 =  ( n157 ) ? ( n47488 ) : ( n47489 ) ;
assign n47491 =  ( n6 ) ? ( n47475 ) : ( n47490 ) ;
assign n47492 =  ( n725 ) ? ( n47491 ) : ( VREG_31_8 ) ;
assign n47493 =  ( n148 ) ? ( n33779 ) : ( VREG_31_9 ) ;
assign n47494 =  ( n146 ) ? ( n33778 ) : ( n47493 ) ;
assign n47495 =  ( n144 ) ? ( n33777 ) : ( n47494 ) ;
assign n47496 =  ( n142 ) ? ( n33776 ) : ( n47495 ) ;
assign n47497 =  ( n10 ) ? ( n33775 ) : ( n47496 ) ;
assign n47498 =  ( n148 ) ? ( n34813 ) : ( VREG_31_9 ) ;
assign n47499 =  ( n146 ) ? ( n34812 ) : ( n47498 ) ;
assign n47500 =  ( n144 ) ? ( n34811 ) : ( n47499 ) ;
assign n47501 =  ( n142 ) ? ( n34810 ) : ( n47500 ) ;
assign n47502 =  ( n10 ) ? ( n34809 ) : ( n47501 ) ;
assign n47503 =  ( n34820 ) ? ( VREG_31_9 ) : ( n47497 ) ;
assign n47504 =  ( n34820 ) ? ( VREG_31_9 ) : ( n47502 ) ;
assign n47505 =  ( n3034 ) ? ( n47504 ) : ( VREG_31_9 ) ;
assign n47506 =  ( n2965 ) ? ( n47503 ) : ( n47505 ) ;
assign n47507 =  ( n1930 ) ? ( n47502 ) : ( n47506 ) ;
assign n47508 =  ( n879 ) ? ( n47497 ) : ( n47507 ) ;
assign n47509 =  ( n172 ) ? ( n34831 ) : ( VREG_31_9 ) ;
assign n47510 =  ( n170 ) ? ( n34830 ) : ( n47509 ) ;
assign n47511 =  ( n168 ) ? ( n34829 ) : ( n47510 ) ;
assign n47512 =  ( n166 ) ? ( n34828 ) : ( n47511 ) ;
assign n47513 =  ( n162 ) ? ( n34827 ) : ( n47512 ) ;
assign n47514 =  ( n172 ) ? ( n34841 ) : ( VREG_31_9 ) ;
assign n47515 =  ( n170 ) ? ( n34840 ) : ( n47514 ) ;
assign n47516 =  ( n168 ) ? ( n34839 ) : ( n47515 ) ;
assign n47517 =  ( n166 ) ? ( n34838 ) : ( n47516 ) ;
assign n47518 =  ( n162 ) ? ( n34837 ) : ( n47517 ) ;
assign n47519 =  ( n34820 ) ? ( VREG_31_9 ) : ( n47518 ) ;
assign n47520 =  ( n3051 ) ? ( n47519 ) : ( VREG_31_9 ) ;
assign n47521 =  ( n3040 ) ? ( n47513 ) : ( n47520 ) ;
assign n47522 =  ( n192 ) ? ( VREG_31_9 ) : ( VREG_31_9 ) ;
assign n47523 =  ( n157 ) ? ( n47521 ) : ( n47522 ) ;
assign n47524 =  ( n6 ) ? ( n47508 ) : ( n47523 ) ;
assign n47525 =  ( n725 ) ? ( n47524 ) : ( VREG_31_9 ) ;
assign n47526 =  ( n148 ) ? ( n1924 ) : ( VREG_3_0 ) ;
assign n47527 =  ( n146 ) ? ( n1923 ) : ( n47526 ) ;
assign n47528 =  ( n144 ) ? ( n1922 ) : ( n47527 ) ;
assign n47529 =  ( n142 ) ? ( n1921 ) : ( n47528 ) ;
assign n47530 =  ( n10 ) ? ( n1920 ) : ( n47529 ) ;
assign n47531 =  ( n148 ) ? ( n2959 ) : ( VREG_3_0 ) ;
assign n47532 =  ( n146 ) ? ( n2958 ) : ( n47531 ) ;
assign n47533 =  ( n144 ) ? ( n2957 ) : ( n47532 ) ;
assign n47534 =  ( n142 ) ? ( n2956 ) : ( n47533 ) ;
assign n47535 =  ( n10 ) ? ( n2955 ) : ( n47534 ) ;
assign n47536 =  ( n3032 ) ? ( VREG_3_0 ) : ( n47530 ) ;
assign n47537 =  ( n3032 ) ? ( VREG_3_0 ) : ( n47535 ) ;
assign n47538 =  ( n3034 ) ? ( n47537 ) : ( VREG_3_0 ) ;
assign n47539 =  ( n2965 ) ? ( n47536 ) : ( n47538 ) ;
assign n47540 =  ( n1930 ) ? ( n47535 ) : ( n47539 ) ;
assign n47541 =  ( n879 ) ? ( n47530 ) : ( n47540 ) ;
assign n47542 =  ( n172 ) ? ( n3045 ) : ( VREG_3_0 ) ;
assign n47543 =  ( n170 ) ? ( n3044 ) : ( n47542 ) ;
assign n47544 =  ( n168 ) ? ( n3043 ) : ( n47543 ) ;
assign n47545 =  ( n166 ) ? ( n3042 ) : ( n47544 ) ;
assign n47546 =  ( n162 ) ? ( n3041 ) : ( n47545 ) ;
assign n47547 =  ( n172 ) ? ( n3056 ) : ( VREG_3_0 ) ;
assign n47548 =  ( n170 ) ? ( n3055 ) : ( n47547 ) ;
assign n47549 =  ( n168 ) ? ( n3054 ) : ( n47548 ) ;
assign n47550 =  ( n166 ) ? ( n3053 ) : ( n47549 ) ;
assign n47551 =  ( n162 ) ? ( n3052 ) : ( n47550 ) ;
assign n47552 =  ( n3032 ) ? ( VREG_3_0 ) : ( n47551 ) ;
assign n47553 =  ( n3051 ) ? ( n47552 ) : ( VREG_3_0 ) ;
assign n47554 =  ( n3040 ) ? ( n47546 ) : ( n47553 ) ;
assign n47555 =  ( n192 ) ? ( VREG_3_0 ) : ( VREG_3_0 ) ;
assign n47556 =  ( n157 ) ? ( n47554 ) : ( n47555 ) ;
assign n47557 =  ( n6 ) ? ( n47541 ) : ( n47556 ) ;
assign n47558 =  ( n681 ) ? ( n47557 ) : ( VREG_3_0 ) ;
assign n47559 =  ( n148 ) ? ( n4113 ) : ( VREG_3_1 ) ;
assign n47560 =  ( n146 ) ? ( n4112 ) : ( n47559 ) ;
assign n47561 =  ( n144 ) ? ( n4111 ) : ( n47560 ) ;
assign n47562 =  ( n142 ) ? ( n4110 ) : ( n47561 ) ;
assign n47563 =  ( n10 ) ? ( n4109 ) : ( n47562 ) ;
assign n47564 =  ( n148 ) ? ( n5147 ) : ( VREG_3_1 ) ;
assign n47565 =  ( n146 ) ? ( n5146 ) : ( n47564 ) ;
assign n47566 =  ( n144 ) ? ( n5145 ) : ( n47565 ) ;
assign n47567 =  ( n142 ) ? ( n5144 ) : ( n47566 ) ;
assign n47568 =  ( n10 ) ? ( n5143 ) : ( n47567 ) ;
assign n47569 =  ( n5154 ) ? ( VREG_3_1 ) : ( n47563 ) ;
assign n47570 =  ( n5154 ) ? ( VREG_3_1 ) : ( n47568 ) ;
assign n47571 =  ( n3034 ) ? ( n47570 ) : ( VREG_3_1 ) ;
assign n47572 =  ( n2965 ) ? ( n47569 ) : ( n47571 ) ;
assign n47573 =  ( n1930 ) ? ( n47568 ) : ( n47572 ) ;
assign n47574 =  ( n879 ) ? ( n47563 ) : ( n47573 ) ;
assign n47575 =  ( n172 ) ? ( n5165 ) : ( VREG_3_1 ) ;
assign n47576 =  ( n170 ) ? ( n5164 ) : ( n47575 ) ;
assign n47577 =  ( n168 ) ? ( n5163 ) : ( n47576 ) ;
assign n47578 =  ( n166 ) ? ( n5162 ) : ( n47577 ) ;
assign n47579 =  ( n162 ) ? ( n5161 ) : ( n47578 ) ;
assign n47580 =  ( n172 ) ? ( n5175 ) : ( VREG_3_1 ) ;
assign n47581 =  ( n170 ) ? ( n5174 ) : ( n47580 ) ;
assign n47582 =  ( n168 ) ? ( n5173 ) : ( n47581 ) ;
assign n47583 =  ( n166 ) ? ( n5172 ) : ( n47582 ) ;
assign n47584 =  ( n162 ) ? ( n5171 ) : ( n47583 ) ;
assign n47585 =  ( n5154 ) ? ( VREG_3_1 ) : ( n47584 ) ;
assign n47586 =  ( n3051 ) ? ( n47585 ) : ( VREG_3_1 ) ;
assign n47587 =  ( n3040 ) ? ( n47579 ) : ( n47586 ) ;
assign n47588 =  ( n192 ) ? ( VREG_3_1 ) : ( VREG_3_1 ) ;
assign n47589 =  ( n157 ) ? ( n47587 ) : ( n47588 ) ;
assign n47590 =  ( n6 ) ? ( n47574 ) : ( n47589 ) ;
assign n47591 =  ( n681 ) ? ( n47590 ) : ( VREG_3_1 ) ;
assign n47592 =  ( n148 ) ? ( n6232 ) : ( VREG_3_10 ) ;
assign n47593 =  ( n146 ) ? ( n6231 ) : ( n47592 ) ;
assign n47594 =  ( n144 ) ? ( n6230 ) : ( n47593 ) ;
assign n47595 =  ( n142 ) ? ( n6229 ) : ( n47594 ) ;
assign n47596 =  ( n10 ) ? ( n6228 ) : ( n47595 ) ;
assign n47597 =  ( n148 ) ? ( n7266 ) : ( VREG_3_10 ) ;
assign n47598 =  ( n146 ) ? ( n7265 ) : ( n47597 ) ;
assign n47599 =  ( n144 ) ? ( n7264 ) : ( n47598 ) ;
assign n47600 =  ( n142 ) ? ( n7263 ) : ( n47599 ) ;
assign n47601 =  ( n10 ) ? ( n7262 ) : ( n47600 ) ;
assign n47602 =  ( n7273 ) ? ( VREG_3_10 ) : ( n47596 ) ;
assign n47603 =  ( n7273 ) ? ( VREG_3_10 ) : ( n47601 ) ;
assign n47604 =  ( n3034 ) ? ( n47603 ) : ( VREG_3_10 ) ;
assign n47605 =  ( n2965 ) ? ( n47602 ) : ( n47604 ) ;
assign n47606 =  ( n1930 ) ? ( n47601 ) : ( n47605 ) ;
assign n47607 =  ( n879 ) ? ( n47596 ) : ( n47606 ) ;
assign n47608 =  ( n172 ) ? ( n7284 ) : ( VREG_3_10 ) ;
assign n47609 =  ( n170 ) ? ( n7283 ) : ( n47608 ) ;
assign n47610 =  ( n168 ) ? ( n7282 ) : ( n47609 ) ;
assign n47611 =  ( n166 ) ? ( n7281 ) : ( n47610 ) ;
assign n47612 =  ( n162 ) ? ( n7280 ) : ( n47611 ) ;
assign n47613 =  ( n172 ) ? ( n7294 ) : ( VREG_3_10 ) ;
assign n47614 =  ( n170 ) ? ( n7293 ) : ( n47613 ) ;
assign n47615 =  ( n168 ) ? ( n7292 ) : ( n47614 ) ;
assign n47616 =  ( n166 ) ? ( n7291 ) : ( n47615 ) ;
assign n47617 =  ( n162 ) ? ( n7290 ) : ( n47616 ) ;
assign n47618 =  ( n7273 ) ? ( VREG_3_10 ) : ( n47617 ) ;
assign n47619 =  ( n3051 ) ? ( n47618 ) : ( VREG_3_10 ) ;
assign n47620 =  ( n3040 ) ? ( n47612 ) : ( n47619 ) ;
assign n47621 =  ( n192 ) ? ( VREG_3_10 ) : ( VREG_3_10 ) ;
assign n47622 =  ( n157 ) ? ( n47620 ) : ( n47621 ) ;
assign n47623 =  ( n6 ) ? ( n47607 ) : ( n47622 ) ;
assign n47624 =  ( n681 ) ? ( n47623 ) : ( VREG_3_10 ) ;
assign n47625 =  ( n148 ) ? ( n8351 ) : ( VREG_3_11 ) ;
assign n47626 =  ( n146 ) ? ( n8350 ) : ( n47625 ) ;
assign n47627 =  ( n144 ) ? ( n8349 ) : ( n47626 ) ;
assign n47628 =  ( n142 ) ? ( n8348 ) : ( n47627 ) ;
assign n47629 =  ( n10 ) ? ( n8347 ) : ( n47628 ) ;
assign n47630 =  ( n148 ) ? ( n9385 ) : ( VREG_3_11 ) ;
assign n47631 =  ( n146 ) ? ( n9384 ) : ( n47630 ) ;
assign n47632 =  ( n144 ) ? ( n9383 ) : ( n47631 ) ;
assign n47633 =  ( n142 ) ? ( n9382 ) : ( n47632 ) ;
assign n47634 =  ( n10 ) ? ( n9381 ) : ( n47633 ) ;
assign n47635 =  ( n9392 ) ? ( VREG_3_11 ) : ( n47629 ) ;
assign n47636 =  ( n9392 ) ? ( VREG_3_11 ) : ( n47634 ) ;
assign n47637 =  ( n3034 ) ? ( n47636 ) : ( VREG_3_11 ) ;
assign n47638 =  ( n2965 ) ? ( n47635 ) : ( n47637 ) ;
assign n47639 =  ( n1930 ) ? ( n47634 ) : ( n47638 ) ;
assign n47640 =  ( n879 ) ? ( n47629 ) : ( n47639 ) ;
assign n47641 =  ( n172 ) ? ( n9403 ) : ( VREG_3_11 ) ;
assign n47642 =  ( n170 ) ? ( n9402 ) : ( n47641 ) ;
assign n47643 =  ( n168 ) ? ( n9401 ) : ( n47642 ) ;
assign n47644 =  ( n166 ) ? ( n9400 ) : ( n47643 ) ;
assign n47645 =  ( n162 ) ? ( n9399 ) : ( n47644 ) ;
assign n47646 =  ( n172 ) ? ( n9413 ) : ( VREG_3_11 ) ;
assign n47647 =  ( n170 ) ? ( n9412 ) : ( n47646 ) ;
assign n47648 =  ( n168 ) ? ( n9411 ) : ( n47647 ) ;
assign n47649 =  ( n166 ) ? ( n9410 ) : ( n47648 ) ;
assign n47650 =  ( n162 ) ? ( n9409 ) : ( n47649 ) ;
assign n47651 =  ( n9392 ) ? ( VREG_3_11 ) : ( n47650 ) ;
assign n47652 =  ( n3051 ) ? ( n47651 ) : ( VREG_3_11 ) ;
assign n47653 =  ( n3040 ) ? ( n47645 ) : ( n47652 ) ;
assign n47654 =  ( n192 ) ? ( VREG_3_11 ) : ( VREG_3_11 ) ;
assign n47655 =  ( n157 ) ? ( n47653 ) : ( n47654 ) ;
assign n47656 =  ( n6 ) ? ( n47640 ) : ( n47655 ) ;
assign n47657 =  ( n681 ) ? ( n47656 ) : ( VREG_3_11 ) ;
assign n47658 =  ( n148 ) ? ( n10470 ) : ( VREG_3_12 ) ;
assign n47659 =  ( n146 ) ? ( n10469 ) : ( n47658 ) ;
assign n47660 =  ( n144 ) ? ( n10468 ) : ( n47659 ) ;
assign n47661 =  ( n142 ) ? ( n10467 ) : ( n47660 ) ;
assign n47662 =  ( n10 ) ? ( n10466 ) : ( n47661 ) ;
assign n47663 =  ( n148 ) ? ( n11504 ) : ( VREG_3_12 ) ;
assign n47664 =  ( n146 ) ? ( n11503 ) : ( n47663 ) ;
assign n47665 =  ( n144 ) ? ( n11502 ) : ( n47664 ) ;
assign n47666 =  ( n142 ) ? ( n11501 ) : ( n47665 ) ;
assign n47667 =  ( n10 ) ? ( n11500 ) : ( n47666 ) ;
assign n47668 =  ( n11511 ) ? ( VREG_3_12 ) : ( n47662 ) ;
assign n47669 =  ( n11511 ) ? ( VREG_3_12 ) : ( n47667 ) ;
assign n47670 =  ( n3034 ) ? ( n47669 ) : ( VREG_3_12 ) ;
assign n47671 =  ( n2965 ) ? ( n47668 ) : ( n47670 ) ;
assign n47672 =  ( n1930 ) ? ( n47667 ) : ( n47671 ) ;
assign n47673 =  ( n879 ) ? ( n47662 ) : ( n47672 ) ;
assign n47674 =  ( n172 ) ? ( n11522 ) : ( VREG_3_12 ) ;
assign n47675 =  ( n170 ) ? ( n11521 ) : ( n47674 ) ;
assign n47676 =  ( n168 ) ? ( n11520 ) : ( n47675 ) ;
assign n47677 =  ( n166 ) ? ( n11519 ) : ( n47676 ) ;
assign n47678 =  ( n162 ) ? ( n11518 ) : ( n47677 ) ;
assign n47679 =  ( n172 ) ? ( n11532 ) : ( VREG_3_12 ) ;
assign n47680 =  ( n170 ) ? ( n11531 ) : ( n47679 ) ;
assign n47681 =  ( n168 ) ? ( n11530 ) : ( n47680 ) ;
assign n47682 =  ( n166 ) ? ( n11529 ) : ( n47681 ) ;
assign n47683 =  ( n162 ) ? ( n11528 ) : ( n47682 ) ;
assign n47684 =  ( n11511 ) ? ( VREG_3_12 ) : ( n47683 ) ;
assign n47685 =  ( n3051 ) ? ( n47684 ) : ( VREG_3_12 ) ;
assign n47686 =  ( n3040 ) ? ( n47678 ) : ( n47685 ) ;
assign n47687 =  ( n192 ) ? ( VREG_3_12 ) : ( VREG_3_12 ) ;
assign n47688 =  ( n157 ) ? ( n47686 ) : ( n47687 ) ;
assign n47689 =  ( n6 ) ? ( n47673 ) : ( n47688 ) ;
assign n47690 =  ( n681 ) ? ( n47689 ) : ( VREG_3_12 ) ;
assign n47691 =  ( n148 ) ? ( n12589 ) : ( VREG_3_13 ) ;
assign n47692 =  ( n146 ) ? ( n12588 ) : ( n47691 ) ;
assign n47693 =  ( n144 ) ? ( n12587 ) : ( n47692 ) ;
assign n47694 =  ( n142 ) ? ( n12586 ) : ( n47693 ) ;
assign n47695 =  ( n10 ) ? ( n12585 ) : ( n47694 ) ;
assign n47696 =  ( n148 ) ? ( n13623 ) : ( VREG_3_13 ) ;
assign n47697 =  ( n146 ) ? ( n13622 ) : ( n47696 ) ;
assign n47698 =  ( n144 ) ? ( n13621 ) : ( n47697 ) ;
assign n47699 =  ( n142 ) ? ( n13620 ) : ( n47698 ) ;
assign n47700 =  ( n10 ) ? ( n13619 ) : ( n47699 ) ;
assign n47701 =  ( n13630 ) ? ( VREG_3_13 ) : ( n47695 ) ;
assign n47702 =  ( n13630 ) ? ( VREG_3_13 ) : ( n47700 ) ;
assign n47703 =  ( n3034 ) ? ( n47702 ) : ( VREG_3_13 ) ;
assign n47704 =  ( n2965 ) ? ( n47701 ) : ( n47703 ) ;
assign n47705 =  ( n1930 ) ? ( n47700 ) : ( n47704 ) ;
assign n47706 =  ( n879 ) ? ( n47695 ) : ( n47705 ) ;
assign n47707 =  ( n172 ) ? ( n13641 ) : ( VREG_3_13 ) ;
assign n47708 =  ( n170 ) ? ( n13640 ) : ( n47707 ) ;
assign n47709 =  ( n168 ) ? ( n13639 ) : ( n47708 ) ;
assign n47710 =  ( n166 ) ? ( n13638 ) : ( n47709 ) ;
assign n47711 =  ( n162 ) ? ( n13637 ) : ( n47710 ) ;
assign n47712 =  ( n172 ) ? ( n13651 ) : ( VREG_3_13 ) ;
assign n47713 =  ( n170 ) ? ( n13650 ) : ( n47712 ) ;
assign n47714 =  ( n168 ) ? ( n13649 ) : ( n47713 ) ;
assign n47715 =  ( n166 ) ? ( n13648 ) : ( n47714 ) ;
assign n47716 =  ( n162 ) ? ( n13647 ) : ( n47715 ) ;
assign n47717 =  ( n13630 ) ? ( VREG_3_13 ) : ( n47716 ) ;
assign n47718 =  ( n3051 ) ? ( n47717 ) : ( VREG_3_13 ) ;
assign n47719 =  ( n3040 ) ? ( n47711 ) : ( n47718 ) ;
assign n47720 =  ( n192 ) ? ( VREG_3_13 ) : ( VREG_3_13 ) ;
assign n47721 =  ( n157 ) ? ( n47719 ) : ( n47720 ) ;
assign n47722 =  ( n6 ) ? ( n47706 ) : ( n47721 ) ;
assign n47723 =  ( n681 ) ? ( n47722 ) : ( VREG_3_13 ) ;
assign n47724 =  ( n148 ) ? ( n14708 ) : ( VREG_3_14 ) ;
assign n47725 =  ( n146 ) ? ( n14707 ) : ( n47724 ) ;
assign n47726 =  ( n144 ) ? ( n14706 ) : ( n47725 ) ;
assign n47727 =  ( n142 ) ? ( n14705 ) : ( n47726 ) ;
assign n47728 =  ( n10 ) ? ( n14704 ) : ( n47727 ) ;
assign n47729 =  ( n148 ) ? ( n15742 ) : ( VREG_3_14 ) ;
assign n47730 =  ( n146 ) ? ( n15741 ) : ( n47729 ) ;
assign n47731 =  ( n144 ) ? ( n15740 ) : ( n47730 ) ;
assign n47732 =  ( n142 ) ? ( n15739 ) : ( n47731 ) ;
assign n47733 =  ( n10 ) ? ( n15738 ) : ( n47732 ) ;
assign n47734 =  ( n15749 ) ? ( VREG_3_14 ) : ( n47728 ) ;
assign n47735 =  ( n15749 ) ? ( VREG_3_14 ) : ( n47733 ) ;
assign n47736 =  ( n3034 ) ? ( n47735 ) : ( VREG_3_14 ) ;
assign n47737 =  ( n2965 ) ? ( n47734 ) : ( n47736 ) ;
assign n47738 =  ( n1930 ) ? ( n47733 ) : ( n47737 ) ;
assign n47739 =  ( n879 ) ? ( n47728 ) : ( n47738 ) ;
assign n47740 =  ( n172 ) ? ( n15760 ) : ( VREG_3_14 ) ;
assign n47741 =  ( n170 ) ? ( n15759 ) : ( n47740 ) ;
assign n47742 =  ( n168 ) ? ( n15758 ) : ( n47741 ) ;
assign n47743 =  ( n166 ) ? ( n15757 ) : ( n47742 ) ;
assign n47744 =  ( n162 ) ? ( n15756 ) : ( n47743 ) ;
assign n47745 =  ( n172 ) ? ( n15770 ) : ( VREG_3_14 ) ;
assign n47746 =  ( n170 ) ? ( n15769 ) : ( n47745 ) ;
assign n47747 =  ( n168 ) ? ( n15768 ) : ( n47746 ) ;
assign n47748 =  ( n166 ) ? ( n15767 ) : ( n47747 ) ;
assign n47749 =  ( n162 ) ? ( n15766 ) : ( n47748 ) ;
assign n47750 =  ( n15749 ) ? ( VREG_3_14 ) : ( n47749 ) ;
assign n47751 =  ( n3051 ) ? ( n47750 ) : ( VREG_3_14 ) ;
assign n47752 =  ( n3040 ) ? ( n47744 ) : ( n47751 ) ;
assign n47753 =  ( n192 ) ? ( VREG_3_14 ) : ( VREG_3_14 ) ;
assign n47754 =  ( n157 ) ? ( n47752 ) : ( n47753 ) ;
assign n47755 =  ( n6 ) ? ( n47739 ) : ( n47754 ) ;
assign n47756 =  ( n681 ) ? ( n47755 ) : ( VREG_3_14 ) ;
assign n47757 =  ( n148 ) ? ( n16827 ) : ( VREG_3_15 ) ;
assign n47758 =  ( n146 ) ? ( n16826 ) : ( n47757 ) ;
assign n47759 =  ( n144 ) ? ( n16825 ) : ( n47758 ) ;
assign n47760 =  ( n142 ) ? ( n16824 ) : ( n47759 ) ;
assign n47761 =  ( n10 ) ? ( n16823 ) : ( n47760 ) ;
assign n47762 =  ( n148 ) ? ( n17861 ) : ( VREG_3_15 ) ;
assign n47763 =  ( n146 ) ? ( n17860 ) : ( n47762 ) ;
assign n47764 =  ( n144 ) ? ( n17859 ) : ( n47763 ) ;
assign n47765 =  ( n142 ) ? ( n17858 ) : ( n47764 ) ;
assign n47766 =  ( n10 ) ? ( n17857 ) : ( n47765 ) ;
assign n47767 =  ( n17868 ) ? ( VREG_3_15 ) : ( n47761 ) ;
assign n47768 =  ( n17868 ) ? ( VREG_3_15 ) : ( n47766 ) ;
assign n47769 =  ( n3034 ) ? ( n47768 ) : ( VREG_3_15 ) ;
assign n47770 =  ( n2965 ) ? ( n47767 ) : ( n47769 ) ;
assign n47771 =  ( n1930 ) ? ( n47766 ) : ( n47770 ) ;
assign n47772 =  ( n879 ) ? ( n47761 ) : ( n47771 ) ;
assign n47773 =  ( n172 ) ? ( n17879 ) : ( VREG_3_15 ) ;
assign n47774 =  ( n170 ) ? ( n17878 ) : ( n47773 ) ;
assign n47775 =  ( n168 ) ? ( n17877 ) : ( n47774 ) ;
assign n47776 =  ( n166 ) ? ( n17876 ) : ( n47775 ) ;
assign n47777 =  ( n162 ) ? ( n17875 ) : ( n47776 ) ;
assign n47778 =  ( n172 ) ? ( n17889 ) : ( VREG_3_15 ) ;
assign n47779 =  ( n170 ) ? ( n17888 ) : ( n47778 ) ;
assign n47780 =  ( n168 ) ? ( n17887 ) : ( n47779 ) ;
assign n47781 =  ( n166 ) ? ( n17886 ) : ( n47780 ) ;
assign n47782 =  ( n162 ) ? ( n17885 ) : ( n47781 ) ;
assign n47783 =  ( n17868 ) ? ( VREG_3_15 ) : ( n47782 ) ;
assign n47784 =  ( n3051 ) ? ( n47783 ) : ( VREG_3_15 ) ;
assign n47785 =  ( n3040 ) ? ( n47777 ) : ( n47784 ) ;
assign n47786 =  ( n192 ) ? ( VREG_3_15 ) : ( VREG_3_15 ) ;
assign n47787 =  ( n157 ) ? ( n47785 ) : ( n47786 ) ;
assign n47788 =  ( n6 ) ? ( n47772 ) : ( n47787 ) ;
assign n47789 =  ( n681 ) ? ( n47788 ) : ( VREG_3_15 ) ;
assign n47790 =  ( n148 ) ? ( n18946 ) : ( VREG_3_2 ) ;
assign n47791 =  ( n146 ) ? ( n18945 ) : ( n47790 ) ;
assign n47792 =  ( n144 ) ? ( n18944 ) : ( n47791 ) ;
assign n47793 =  ( n142 ) ? ( n18943 ) : ( n47792 ) ;
assign n47794 =  ( n10 ) ? ( n18942 ) : ( n47793 ) ;
assign n47795 =  ( n148 ) ? ( n19980 ) : ( VREG_3_2 ) ;
assign n47796 =  ( n146 ) ? ( n19979 ) : ( n47795 ) ;
assign n47797 =  ( n144 ) ? ( n19978 ) : ( n47796 ) ;
assign n47798 =  ( n142 ) ? ( n19977 ) : ( n47797 ) ;
assign n47799 =  ( n10 ) ? ( n19976 ) : ( n47798 ) ;
assign n47800 =  ( n19987 ) ? ( VREG_3_2 ) : ( n47794 ) ;
assign n47801 =  ( n19987 ) ? ( VREG_3_2 ) : ( n47799 ) ;
assign n47802 =  ( n3034 ) ? ( n47801 ) : ( VREG_3_2 ) ;
assign n47803 =  ( n2965 ) ? ( n47800 ) : ( n47802 ) ;
assign n47804 =  ( n1930 ) ? ( n47799 ) : ( n47803 ) ;
assign n47805 =  ( n879 ) ? ( n47794 ) : ( n47804 ) ;
assign n47806 =  ( n172 ) ? ( n19998 ) : ( VREG_3_2 ) ;
assign n47807 =  ( n170 ) ? ( n19997 ) : ( n47806 ) ;
assign n47808 =  ( n168 ) ? ( n19996 ) : ( n47807 ) ;
assign n47809 =  ( n166 ) ? ( n19995 ) : ( n47808 ) ;
assign n47810 =  ( n162 ) ? ( n19994 ) : ( n47809 ) ;
assign n47811 =  ( n172 ) ? ( n20008 ) : ( VREG_3_2 ) ;
assign n47812 =  ( n170 ) ? ( n20007 ) : ( n47811 ) ;
assign n47813 =  ( n168 ) ? ( n20006 ) : ( n47812 ) ;
assign n47814 =  ( n166 ) ? ( n20005 ) : ( n47813 ) ;
assign n47815 =  ( n162 ) ? ( n20004 ) : ( n47814 ) ;
assign n47816 =  ( n19987 ) ? ( VREG_3_2 ) : ( n47815 ) ;
assign n47817 =  ( n3051 ) ? ( n47816 ) : ( VREG_3_2 ) ;
assign n47818 =  ( n3040 ) ? ( n47810 ) : ( n47817 ) ;
assign n47819 =  ( n192 ) ? ( VREG_3_2 ) : ( VREG_3_2 ) ;
assign n47820 =  ( n157 ) ? ( n47818 ) : ( n47819 ) ;
assign n47821 =  ( n6 ) ? ( n47805 ) : ( n47820 ) ;
assign n47822 =  ( n681 ) ? ( n47821 ) : ( VREG_3_2 ) ;
assign n47823 =  ( n148 ) ? ( n21065 ) : ( VREG_3_3 ) ;
assign n47824 =  ( n146 ) ? ( n21064 ) : ( n47823 ) ;
assign n47825 =  ( n144 ) ? ( n21063 ) : ( n47824 ) ;
assign n47826 =  ( n142 ) ? ( n21062 ) : ( n47825 ) ;
assign n47827 =  ( n10 ) ? ( n21061 ) : ( n47826 ) ;
assign n47828 =  ( n148 ) ? ( n22099 ) : ( VREG_3_3 ) ;
assign n47829 =  ( n146 ) ? ( n22098 ) : ( n47828 ) ;
assign n47830 =  ( n144 ) ? ( n22097 ) : ( n47829 ) ;
assign n47831 =  ( n142 ) ? ( n22096 ) : ( n47830 ) ;
assign n47832 =  ( n10 ) ? ( n22095 ) : ( n47831 ) ;
assign n47833 =  ( n22106 ) ? ( VREG_3_3 ) : ( n47827 ) ;
assign n47834 =  ( n22106 ) ? ( VREG_3_3 ) : ( n47832 ) ;
assign n47835 =  ( n3034 ) ? ( n47834 ) : ( VREG_3_3 ) ;
assign n47836 =  ( n2965 ) ? ( n47833 ) : ( n47835 ) ;
assign n47837 =  ( n1930 ) ? ( n47832 ) : ( n47836 ) ;
assign n47838 =  ( n879 ) ? ( n47827 ) : ( n47837 ) ;
assign n47839 =  ( n172 ) ? ( n22117 ) : ( VREG_3_3 ) ;
assign n47840 =  ( n170 ) ? ( n22116 ) : ( n47839 ) ;
assign n47841 =  ( n168 ) ? ( n22115 ) : ( n47840 ) ;
assign n47842 =  ( n166 ) ? ( n22114 ) : ( n47841 ) ;
assign n47843 =  ( n162 ) ? ( n22113 ) : ( n47842 ) ;
assign n47844 =  ( n172 ) ? ( n22127 ) : ( VREG_3_3 ) ;
assign n47845 =  ( n170 ) ? ( n22126 ) : ( n47844 ) ;
assign n47846 =  ( n168 ) ? ( n22125 ) : ( n47845 ) ;
assign n47847 =  ( n166 ) ? ( n22124 ) : ( n47846 ) ;
assign n47848 =  ( n162 ) ? ( n22123 ) : ( n47847 ) ;
assign n47849 =  ( n22106 ) ? ( VREG_3_3 ) : ( n47848 ) ;
assign n47850 =  ( n3051 ) ? ( n47849 ) : ( VREG_3_3 ) ;
assign n47851 =  ( n3040 ) ? ( n47843 ) : ( n47850 ) ;
assign n47852 =  ( n192 ) ? ( VREG_3_3 ) : ( VREG_3_3 ) ;
assign n47853 =  ( n157 ) ? ( n47851 ) : ( n47852 ) ;
assign n47854 =  ( n6 ) ? ( n47838 ) : ( n47853 ) ;
assign n47855 =  ( n681 ) ? ( n47854 ) : ( VREG_3_3 ) ;
assign n47856 =  ( n148 ) ? ( n23184 ) : ( VREG_3_4 ) ;
assign n47857 =  ( n146 ) ? ( n23183 ) : ( n47856 ) ;
assign n47858 =  ( n144 ) ? ( n23182 ) : ( n47857 ) ;
assign n47859 =  ( n142 ) ? ( n23181 ) : ( n47858 ) ;
assign n47860 =  ( n10 ) ? ( n23180 ) : ( n47859 ) ;
assign n47861 =  ( n148 ) ? ( n24218 ) : ( VREG_3_4 ) ;
assign n47862 =  ( n146 ) ? ( n24217 ) : ( n47861 ) ;
assign n47863 =  ( n144 ) ? ( n24216 ) : ( n47862 ) ;
assign n47864 =  ( n142 ) ? ( n24215 ) : ( n47863 ) ;
assign n47865 =  ( n10 ) ? ( n24214 ) : ( n47864 ) ;
assign n47866 =  ( n24225 ) ? ( VREG_3_4 ) : ( n47860 ) ;
assign n47867 =  ( n24225 ) ? ( VREG_3_4 ) : ( n47865 ) ;
assign n47868 =  ( n3034 ) ? ( n47867 ) : ( VREG_3_4 ) ;
assign n47869 =  ( n2965 ) ? ( n47866 ) : ( n47868 ) ;
assign n47870 =  ( n1930 ) ? ( n47865 ) : ( n47869 ) ;
assign n47871 =  ( n879 ) ? ( n47860 ) : ( n47870 ) ;
assign n47872 =  ( n172 ) ? ( n24236 ) : ( VREG_3_4 ) ;
assign n47873 =  ( n170 ) ? ( n24235 ) : ( n47872 ) ;
assign n47874 =  ( n168 ) ? ( n24234 ) : ( n47873 ) ;
assign n47875 =  ( n166 ) ? ( n24233 ) : ( n47874 ) ;
assign n47876 =  ( n162 ) ? ( n24232 ) : ( n47875 ) ;
assign n47877 =  ( n172 ) ? ( n24246 ) : ( VREG_3_4 ) ;
assign n47878 =  ( n170 ) ? ( n24245 ) : ( n47877 ) ;
assign n47879 =  ( n168 ) ? ( n24244 ) : ( n47878 ) ;
assign n47880 =  ( n166 ) ? ( n24243 ) : ( n47879 ) ;
assign n47881 =  ( n162 ) ? ( n24242 ) : ( n47880 ) ;
assign n47882 =  ( n24225 ) ? ( VREG_3_4 ) : ( n47881 ) ;
assign n47883 =  ( n3051 ) ? ( n47882 ) : ( VREG_3_4 ) ;
assign n47884 =  ( n3040 ) ? ( n47876 ) : ( n47883 ) ;
assign n47885 =  ( n192 ) ? ( VREG_3_4 ) : ( VREG_3_4 ) ;
assign n47886 =  ( n157 ) ? ( n47884 ) : ( n47885 ) ;
assign n47887 =  ( n6 ) ? ( n47871 ) : ( n47886 ) ;
assign n47888 =  ( n681 ) ? ( n47887 ) : ( VREG_3_4 ) ;
assign n47889 =  ( n148 ) ? ( n25303 ) : ( VREG_3_5 ) ;
assign n47890 =  ( n146 ) ? ( n25302 ) : ( n47889 ) ;
assign n47891 =  ( n144 ) ? ( n25301 ) : ( n47890 ) ;
assign n47892 =  ( n142 ) ? ( n25300 ) : ( n47891 ) ;
assign n47893 =  ( n10 ) ? ( n25299 ) : ( n47892 ) ;
assign n47894 =  ( n148 ) ? ( n26337 ) : ( VREG_3_5 ) ;
assign n47895 =  ( n146 ) ? ( n26336 ) : ( n47894 ) ;
assign n47896 =  ( n144 ) ? ( n26335 ) : ( n47895 ) ;
assign n47897 =  ( n142 ) ? ( n26334 ) : ( n47896 ) ;
assign n47898 =  ( n10 ) ? ( n26333 ) : ( n47897 ) ;
assign n47899 =  ( n26344 ) ? ( VREG_3_5 ) : ( n47893 ) ;
assign n47900 =  ( n26344 ) ? ( VREG_3_5 ) : ( n47898 ) ;
assign n47901 =  ( n3034 ) ? ( n47900 ) : ( VREG_3_5 ) ;
assign n47902 =  ( n2965 ) ? ( n47899 ) : ( n47901 ) ;
assign n47903 =  ( n1930 ) ? ( n47898 ) : ( n47902 ) ;
assign n47904 =  ( n879 ) ? ( n47893 ) : ( n47903 ) ;
assign n47905 =  ( n172 ) ? ( n26355 ) : ( VREG_3_5 ) ;
assign n47906 =  ( n170 ) ? ( n26354 ) : ( n47905 ) ;
assign n47907 =  ( n168 ) ? ( n26353 ) : ( n47906 ) ;
assign n47908 =  ( n166 ) ? ( n26352 ) : ( n47907 ) ;
assign n47909 =  ( n162 ) ? ( n26351 ) : ( n47908 ) ;
assign n47910 =  ( n172 ) ? ( n26365 ) : ( VREG_3_5 ) ;
assign n47911 =  ( n170 ) ? ( n26364 ) : ( n47910 ) ;
assign n47912 =  ( n168 ) ? ( n26363 ) : ( n47911 ) ;
assign n47913 =  ( n166 ) ? ( n26362 ) : ( n47912 ) ;
assign n47914 =  ( n162 ) ? ( n26361 ) : ( n47913 ) ;
assign n47915 =  ( n26344 ) ? ( VREG_3_5 ) : ( n47914 ) ;
assign n47916 =  ( n3051 ) ? ( n47915 ) : ( VREG_3_5 ) ;
assign n47917 =  ( n3040 ) ? ( n47909 ) : ( n47916 ) ;
assign n47918 =  ( n192 ) ? ( VREG_3_5 ) : ( VREG_3_5 ) ;
assign n47919 =  ( n157 ) ? ( n47917 ) : ( n47918 ) ;
assign n47920 =  ( n6 ) ? ( n47904 ) : ( n47919 ) ;
assign n47921 =  ( n681 ) ? ( n47920 ) : ( VREG_3_5 ) ;
assign n47922 =  ( n148 ) ? ( n27422 ) : ( VREG_3_6 ) ;
assign n47923 =  ( n146 ) ? ( n27421 ) : ( n47922 ) ;
assign n47924 =  ( n144 ) ? ( n27420 ) : ( n47923 ) ;
assign n47925 =  ( n142 ) ? ( n27419 ) : ( n47924 ) ;
assign n47926 =  ( n10 ) ? ( n27418 ) : ( n47925 ) ;
assign n47927 =  ( n148 ) ? ( n28456 ) : ( VREG_3_6 ) ;
assign n47928 =  ( n146 ) ? ( n28455 ) : ( n47927 ) ;
assign n47929 =  ( n144 ) ? ( n28454 ) : ( n47928 ) ;
assign n47930 =  ( n142 ) ? ( n28453 ) : ( n47929 ) ;
assign n47931 =  ( n10 ) ? ( n28452 ) : ( n47930 ) ;
assign n47932 =  ( n28463 ) ? ( VREG_3_6 ) : ( n47926 ) ;
assign n47933 =  ( n28463 ) ? ( VREG_3_6 ) : ( n47931 ) ;
assign n47934 =  ( n3034 ) ? ( n47933 ) : ( VREG_3_6 ) ;
assign n47935 =  ( n2965 ) ? ( n47932 ) : ( n47934 ) ;
assign n47936 =  ( n1930 ) ? ( n47931 ) : ( n47935 ) ;
assign n47937 =  ( n879 ) ? ( n47926 ) : ( n47936 ) ;
assign n47938 =  ( n172 ) ? ( n28474 ) : ( VREG_3_6 ) ;
assign n47939 =  ( n170 ) ? ( n28473 ) : ( n47938 ) ;
assign n47940 =  ( n168 ) ? ( n28472 ) : ( n47939 ) ;
assign n47941 =  ( n166 ) ? ( n28471 ) : ( n47940 ) ;
assign n47942 =  ( n162 ) ? ( n28470 ) : ( n47941 ) ;
assign n47943 =  ( n172 ) ? ( n28484 ) : ( VREG_3_6 ) ;
assign n47944 =  ( n170 ) ? ( n28483 ) : ( n47943 ) ;
assign n47945 =  ( n168 ) ? ( n28482 ) : ( n47944 ) ;
assign n47946 =  ( n166 ) ? ( n28481 ) : ( n47945 ) ;
assign n47947 =  ( n162 ) ? ( n28480 ) : ( n47946 ) ;
assign n47948 =  ( n28463 ) ? ( VREG_3_6 ) : ( n47947 ) ;
assign n47949 =  ( n3051 ) ? ( n47948 ) : ( VREG_3_6 ) ;
assign n47950 =  ( n3040 ) ? ( n47942 ) : ( n47949 ) ;
assign n47951 =  ( n192 ) ? ( VREG_3_6 ) : ( VREG_3_6 ) ;
assign n47952 =  ( n157 ) ? ( n47950 ) : ( n47951 ) ;
assign n47953 =  ( n6 ) ? ( n47937 ) : ( n47952 ) ;
assign n47954 =  ( n681 ) ? ( n47953 ) : ( VREG_3_6 ) ;
assign n47955 =  ( n148 ) ? ( n29541 ) : ( VREG_3_7 ) ;
assign n47956 =  ( n146 ) ? ( n29540 ) : ( n47955 ) ;
assign n47957 =  ( n144 ) ? ( n29539 ) : ( n47956 ) ;
assign n47958 =  ( n142 ) ? ( n29538 ) : ( n47957 ) ;
assign n47959 =  ( n10 ) ? ( n29537 ) : ( n47958 ) ;
assign n47960 =  ( n148 ) ? ( n30575 ) : ( VREG_3_7 ) ;
assign n47961 =  ( n146 ) ? ( n30574 ) : ( n47960 ) ;
assign n47962 =  ( n144 ) ? ( n30573 ) : ( n47961 ) ;
assign n47963 =  ( n142 ) ? ( n30572 ) : ( n47962 ) ;
assign n47964 =  ( n10 ) ? ( n30571 ) : ( n47963 ) ;
assign n47965 =  ( n30582 ) ? ( VREG_3_7 ) : ( n47959 ) ;
assign n47966 =  ( n30582 ) ? ( VREG_3_7 ) : ( n47964 ) ;
assign n47967 =  ( n3034 ) ? ( n47966 ) : ( VREG_3_7 ) ;
assign n47968 =  ( n2965 ) ? ( n47965 ) : ( n47967 ) ;
assign n47969 =  ( n1930 ) ? ( n47964 ) : ( n47968 ) ;
assign n47970 =  ( n879 ) ? ( n47959 ) : ( n47969 ) ;
assign n47971 =  ( n172 ) ? ( n30593 ) : ( VREG_3_7 ) ;
assign n47972 =  ( n170 ) ? ( n30592 ) : ( n47971 ) ;
assign n47973 =  ( n168 ) ? ( n30591 ) : ( n47972 ) ;
assign n47974 =  ( n166 ) ? ( n30590 ) : ( n47973 ) ;
assign n47975 =  ( n162 ) ? ( n30589 ) : ( n47974 ) ;
assign n47976 =  ( n172 ) ? ( n30603 ) : ( VREG_3_7 ) ;
assign n47977 =  ( n170 ) ? ( n30602 ) : ( n47976 ) ;
assign n47978 =  ( n168 ) ? ( n30601 ) : ( n47977 ) ;
assign n47979 =  ( n166 ) ? ( n30600 ) : ( n47978 ) ;
assign n47980 =  ( n162 ) ? ( n30599 ) : ( n47979 ) ;
assign n47981 =  ( n30582 ) ? ( VREG_3_7 ) : ( n47980 ) ;
assign n47982 =  ( n3051 ) ? ( n47981 ) : ( VREG_3_7 ) ;
assign n47983 =  ( n3040 ) ? ( n47975 ) : ( n47982 ) ;
assign n47984 =  ( n192 ) ? ( VREG_3_7 ) : ( VREG_3_7 ) ;
assign n47985 =  ( n157 ) ? ( n47983 ) : ( n47984 ) ;
assign n47986 =  ( n6 ) ? ( n47970 ) : ( n47985 ) ;
assign n47987 =  ( n681 ) ? ( n47986 ) : ( VREG_3_7 ) ;
assign n47988 =  ( n148 ) ? ( n31660 ) : ( VREG_3_8 ) ;
assign n47989 =  ( n146 ) ? ( n31659 ) : ( n47988 ) ;
assign n47990 =  ( n144 ) ? ( n31658 ) : ( n47989 ) ;
assign n47991 =  ( n142 ) ? ( n31657 ) : ( n47990 ) ;
assign n47992 =  ( n10 ) ? ( n31656 ) : ( n47991 ) ;
assign n47993 =  ( n148 ) ? ( n32694 ) : ( VREG_3_8 ) ;
assign n47994 =  ( n146 ) ? ( n32693 ) : ( n47993 ) ;
assign n47995 =  ( n144 ) ? ( n32692 ) : ( n47994 ) ;
assign n47996 =  ( n142 ) ? ( n32691 ) : ( n47995 ) ;
assign n47997 =  ( n10 ) ? ( n32690 ) : ( n47996 ) ;
assign n47998 =  ( n32701 ) ? ( VREG_3_8 ) : ( n47992 ) ;
assign n47999 =  ( n32701 ) ? ( VREG_3_8 ) : ( n47997 ) ;
assign n48000 =  ( n3034 ) ? ( n47999 ) : ( VREG_3_8 ) ;
assign n48001 =  ( n2965 ) ? ( n47998 ) : ( n48000 ) ;
assign n48002 =  ( n1930 ) ? ( n47997 ) : ( n48001 ) ;
assign n48003 =  ( n879 ) ? ( n47992 ) : ( n48002 ) ;
assign n48004 =  ( n172 ) ? ( n32712 ) : ( VREG_3_8 ) ;
assign n48005 =  ( n170 ) ? ( n32711 ) : ( n48004 ) ;
assign n48006 =  ( n168 ) ? ( n32710 ) : ( n48005 ) ;
assign n48007 =  ( n166 ) ? ( n32709 ) : ( n48006 ) ;
assign n48008 =  ( n162 ) ? ( n32708 ) : ( n48007 ) ;
assign n48009 =  ( n172 ) ? ( n32722 ) : ( VREG_3_8 ) ;
assign n48010 =  ( n170 ) ? ( n32721 ) : ( n48009 ) ;
assign n48011 =  ( n168 ) ? ( n32720 ) : ( n48010 ) ;
assign n48012 =  ( n166 ) ? ( n32719 ) : ( n48011 ) ;
assign n48013 =  ( n162 ) ? ( n32718 ) : ( n48012 ) ;
assign n48014 =  ( n32701 ) ? ( VREG_3_8 ) : ( n48013 ) ;
assign n48015 =  ( n3051 ) ? ( n48014 ) : ( VREG_3_8 ) ;
assign n48016 =  ( n3040 ) ? ( n48008 ) : ( n48015 ) ;
assign n48017 =  ( n192 ) ? ( VREG_3_8 ) : ( VREG_3_8 ) ;
assign n48018 =  ( n157 ) ? ( n48016 ) : ( n48017 ) ;
assign n48019 =  ( n6 ) ? ( n48003 ) : ( n48018 ) ;
assign n48020 =  ( n681 ) ? ( n48019 ) : ( VREG_3_8 ) ;
assign n48021 =  ( n148 ) ? ( n33779 ) : ( VREG_3_9 ) ;
assign n48022 =  ( n146 ) ? ( n33778 ) : ( n48021 ) ;
assign n48023 =  ( n144 ) ? ( n33777 ) : ( n48022 ) ;
assign n48024 =  ( n142 ) ? ( n33776 ) : ( n48023 ) ;
assign n48025 =  ( n10 ) ? ( n33775 ) : ( n48024 ) ;
assign n48026 =  ( n148 ) ? ( n34813 ) : ( VREG_3_9 ) ;
assign n48027 =  ( n146 ) ? ( n34812 ) : ( n48026 ) ;
assign n48028 =  ( n144 ) ? ( n34811 ) : ( n48027 ) ;
assign n48029 =  ( n142 ) ? ( n34810 ) : ( n48028 ) ;
assign n48030 =  ( n10 ) ? ( n34809 ) : ( n48029 ) ;
assign n48031 =  ( n34820 ) ? ( VREG_3_9 ) : ( n48025 ) ;
assign n48032 =  ( n34820 ) ? ( VREG_3_9 ) : ( n48030 ) ;
assign n48033 =  ( n3034 ) ? ( n48032 ) : ( VREG_3_9 ) ;
assign n48034 =  ( n2965 ) ? ( n48031 ) : ( n48033 ) ;
assign n48035 =  ( n1930 ) ? ( n48030 ) : ( n48034 ) ;
assign n48036 =  ( n879 ) ? ( n48025 ) : ( n48035 ) ;
assign n48037 =  ( n172 ) ? ( n34831 ) : ( VREG_3_9 ) ;
assign n48038 =  ( n170 ) ? ( n34830 ) : ( n48037 ) ;
assign n48039 =  ( n168 ) ? ( n34829 ) : ( n48038 ) ;
assign n48040 =  ( n166 ) ? ( n34828 ) : ( n48039 ) ;
assign n48041 =  ( n162 ) ? ( n34827 ) : ( n48040 ) ;
assign n48042 =  ( n172 ) ? ( n34841 ) : ( VREG_3_9 ) ;
assign n48043 =  ( n170 ) ? ( n34840 ) : ( n48042 ) ;
assign n48044 =  ( n168 ) ? ( n34839 ) : ( n48043 ) ;
assign n48045 =  ( n166 ) ? ( n34838 ) : ( n48044 ) ;
assign n48046 =  ( n162 ) ? ( n34837 ) : ( n48045 ) ;
assign n48047 =  ( n34820 ) ? ( VREG_3_9 ) : ( n48046 ) ;
assign n48048 =  ( n3051 ) ? ( n48047 ) : ( VREG_3_9 ) ;
assign n48049 =  ( n3040 ) ? ( n48041 ) : ( n48048 ) ;
assign n48050 =  ( n192 ) ? ( VREG_3_9 ) : ( VREG_3_9 ) ;
assign n48051 =  ( n157 ) ? ( n48049 ) : ( n48050 ) ;
assign n48052 =  ( n6 ) ? ( n48036 ) : ( n48051 ) ;
assign n48053 =  ( n681 ) ? ( n48052 ) : ( VREG_3_9 ) ;
assign n48054 =  ( n148 ) ? ( n1924 ) : ( VREG_4_0 ) ;
assign n48055 =  ( n146 ) ? ( n1923 ) : ( n48054 ) ;
assign n48056 =  ( n144 ) ? ( n1922 ) : ( n48055 ) ;
assign n48057 =  ( n142 ) ? ( n1921 ) : ( n48056 ) ;
assign n48058 =  ( n10 ) ? ( n1920 ) : ( n48057 ) ;
assign n48059 =  ( n148 ) ? ( n2959 ) : ( VREG_4_0 ) ;
assign n48060 =  ( n146 ) ? ( n2958 ) : ( n48059 ) ;
assign n48061 =  ( n144 ) ? ( n2957 ) : ( n48060 ) ;
assign n48062 =  ( n142 ) ? ( n2956 ) : ( n48061 ) ;
assign n48063 =  ( n10 ) ? ( n2955 ) : ( n48062 ) ;
assign n48064 =  ( n3032 ) ? ( VREG_4_0 ) : ( n48058 ) ;
assign n48065 =  ( n3032 ) ? ( VREG_4_0 ) : ( n48063 ) ;
assign n48066 =  ( n3034 ) ? ( n48065 ) : ( VREG_4_0 ) ;
assign n48067 =  ( n2965 ) ? ( n48064 ) : ( n48066 ) ;
assign n48068 =  ( n1930 ) ? ( n48063 ) : ( n48067 ) ;
assign n48069 =  ( n879 ) ? ( n48058 ) : ( n48068 ) ;
assign n48070 =  ( n172 ) ? ( n3045 ) : ( VREG_4_0 ) ;
assign n48071 =  ( n170 ) ? ( n3044 ) : ( n48070 ) ;
assign n48072 =  ( n168 ) ? ( n3043 ) : ( n48071 ) ;
assign n48073 =  ( n166 ) ? ( n3042 ) : ( n48072 ) ;
assign n48074 =  ( n162 ) ? ( n3041 ) : ( n48073 ) ;
assign n48075 =  ( n172 ) ? ( n3056 ) : ( VREG_4_0 ) ;
assign n48076 =  ( n170 ) ? ( n3055 ) : ( n48075 ) ;
assign n48077 =  ( n168 ) ? ( n3054 ) : ( n48076 ) ;
assign n48078 =  ( n166 ) ? ( n3053 ) : ( n48077 ) ;
assign n48079 =  ( n162 ) ? ( n3052 ) : ( n48078 ) ;
assign n48080 =  ( n3032 ) ? ( VREG_4_0 ) : ( n48079 ) ;
assign n48081 =  ( n3051 ) ? ( n48080 ) : ( VREG_4_0 ) ;
assign n48082 =  ( n3040 ) ? ( n48074 ) : ( n48081 ) ;
assign n48083 =  ( n192 ) ? ( VREG_4_0 ) : ( VREG_4_0 ) ;
assign n48084 =  ( n157 ) ? ( n48082 ) : ( n48083 ) ;
assign n48085 =  ( n6 ) ? ( n48069 ) : ( n48084 ) ;
assign n48086 =  ( n747 ) ? ( n48085 ) : ( VREG_4_0 ) ;
assign n48087 =  ( n148 ) ? ( n4113 ) : ( VREG_4_1 ) ;
assign n48088 =  ( n146 ) ? ( n4112 ) : ( n48087 ) ;
assign n48089 =  ( n144 ) ? ( n4111 ) : ( n48088 ) ;
assign n48090 =  ( n142 ) ? ( n4110 ) : ( n48089 ) ;
assign n48091 =  ( n10 ) ? ( n4109 ) : ( n48090 ) ;
assign n48092 =  ( n148 ) ? ( n5147 ) : ( VREG_4_1 ) ;
assign n48093 =  ( n146 ) ? ( n5146 ) : ( n48092 ) ;
assign n48094 =  ( n144 ) ? ( n5145 ) : ( n48093 ) ;
assign n48095 =  ( n142 ) ? ( n5144 ) : ( n48094 ) ;
assign n48096 =  ( n10 ) ? ( n5143 ) : ( n48095 ) ;
assign n48097 =  ( n5154 ) ? ( VREG_4_1 ) : ( n48091 ) ;
assign n48098 =  ( n5154 ) ? ( VREG_4_1 ) : ( n48096 ) ;
assign n48099 =  ( n3034 ) ? ( n48098 ) : ( VREG_4_1 ) ;
assign n48100 =  ( n2965 ) ? ( n48097 ) : ( n48099 ) ;
assign n48101 =  ( n1930 ) ? ( n48096 ) : ( n48100 ) ;
assign n48102 =  ( n879 ) ? ( n48091 ) : ( n48101 ) ;
assign n48103 =  ( n172 ) ? ( n5165 ) : ( VREG_4_1 ) ;
assign n48104 =  ( n170 ) ? ( n5164 ) : ( n48103 ) ;
assign n48105 =  ( n168 ) ? ( n5163 ) : ( n48104 ) ;
assign n48106 =  ( n166 ) ? ( n5162 ) : ( n48105 ) ;
assign n48107 =  ( n162 ) ? ( n5161 ) : ( n48106 ) ;
assign n48108 =  ( n172 ) ? ( n5175 ) : ( VREG_4_1 ) ;
assign n48109 =  ( n170 ) ? ( n5174 ) : ( n48108 ) ;
assign n48110 =  ( n168 ) ? ( n5173 ) : ( n48109 ) ;
assign n48111 =  ( n166 ) ? ( n5172 ) : ( n48110 ) ;
assign n48112 =  ( n162 ) ? ( n5171 ) : ( n48111 ) ;
assign n48113 =  ( n5154 ) ? ( VREG_4_1 ) : ( n48112 ) ;
assign n48114 =  ( n3051 ) ? ( n48113 ) : ( VREG_4_1 ) ;
assign n48115 =  ( n3040 ) ? ( n48107 ) : ( n48114 ) ;
assign n48116 =  ( n192 ) ? ( VREG_4_1 ) : ( VREG_4_1 ) ;
assign n48117 =  ( n157 ) ? ( n48115 ) : ( n48116 ) ;
assign n48118 =  ( n6 ) ? ( n48102 ) : ( n48117 ) ;
assign n48119 =  ( n747 ) ? ( n48118 ) : ( VREG_4_1 ) ;
assign n48120 =  ( n148 ) ? ( n6232 ) : ( VREG_4_10 ) ;
assign n48121 =  ( n146 ) ? ( n6231 ) : ( n48120 ) ;
assign n48122 =  ( n144 ) ? ( n6230 ) : ( n48121 ) ;
assign n48123 =  ( n142 ) ? ( n6229 ) : ( n48122 ) ;
assign n48124 =  ( n10 ) ? ( n6228 ) : ( n48123 ) ;
assign n48125 =  ( n148 ) ? ( n7266 ) : ( VREG_4_10 ) ;
assign n48126 =  ( n146 ) ? ( n7265 ) : ( n48125 ) ;
assign n48127 =  ( n144 ) ? ( n7264 ) : ( n48126 ) ;
assign n48128 =  ( n142 ) ? ( n7263 ) : ( n48127 ) ;
assign n48129 =  ( n10 ) ? ( n7262 ) : ( n48128 ) ;
assign n48130 =  ( n7273 ) ? ( VREG_4_10 ) : ( n48124 ) ;
assign n48131 =  ( n7273 ) ? ( VREG_4_10 ) : ( n48129 ) ;
assign n48132 =  ( n3034 ) ? ( n48131 ) : ( VREG_4_10 ) ;
assign n48133 =  ( n2965 ) ? ( n48130 ) : ( n48132 ) ;
assign n48134 =  ( n1930 ) ? ( n48129 ) : ( n48133 ) ;
assign n48135 =  ( n879 ) ? ( n48124 ) : ( n48134 ) ;
assign n48136 =  ( n172 ) ? ( n7284 ) : ( VREG_4_10 ) ;
assign n48137 =  ( n170 ) ? ( n7283 ) : ( n48136 ) ;
assign n48138 =  ( n168 ) ? ( n7282 ) : ( n48137 ) ;
assign n48139 =  ( n166 ) ? ( n7281 ) : ( n48138 ) ;
assign n48140 =  ( n162 ) ? ( n7280 ) : ( n48139 ) ;
assign n48141 =  ( n172 ) ? ( n7294 ) : ( VREG_4_10 ) ;
assign n48142 =  ( n170 ) ? ( n7293 ) : ( n48141 ) ;
assign n48143 =  ( n168 ) ? ( n7292 ) : ( n48142 ) ;
assign n48144 =  ( n166 ) ? ( n7291 ) : ( n48143 ) ;
assign n48145 =  ( n162 ) ? ( n7290 ) : ( n48144 ) ;
assign n48146 =  ( n7273 ) ? ( VREG_4_10 ) : ( n48145 ) ;
assign n48147 =  ( n3051 ) ? ( n48146 ) : ( VREG_4_10 ) ;
assign n48148 =  ( n3040 ) ? ( n48140 ) : ( n48147 ) ;
assign n48149 =  ( n192 ) ? ( VREG_4_10 ) : ( VREG_4_10 ) ;
assign n48150 =  ( n157 ) ? ( n48148 ) : ( n48149 ) ;
assign n48151 =  ( n6 ) ? ( n48135 ) : ( n48150 ) ;
assign n48152 =  ( n747 ) ? ( n48151 ) : ( VREG_4_10 ) ;
assign n48153 =  ( n148 ) ? ( n8351 ) : ( VREG_4_11 ) ;
assign n48154 =  ( n146 ) ? ( n8350 ) : ( n48153 ) ;
assign n48155 =  ( n144 ) ? ( n8349 ) : ( n48154 ) ;
assign n48156 =  ( n142 ) ? ( n8348 ) : ( n48155 ) ;
assign n48157 =  ( n10 ) ? ( n8347 ) : ( n48156 ) ;
assign n48158 =  ( n148 ) ? ( n9385 ) : ( VREG_4_11 ) ;
assign n48159 =  ( n146 ) ? ( n9384 ) : ( n48158 ) ;
assign n48160 =  ( n144 ) ? ( n9383 ) : ( n48159 ) ;
assign n48161 =  ( n142 ) ? ( n9382 ) : ( n48160 ) ;
assign n48162 =  ( n10 ) ? ( n9381 ) : ( n48161 ) ;
assign n48163 =  ( n9392 ) ? ( VREG_4_11 ) : ( n48157 ) ;
assign n48164 =  ( n9392 ) ? ( VREG_4_11 ) : ( n48162 ) ;
assign n48165 =  ( n3034 ) ? ( n48164 ) : ( VREG_4_11 ) ;
assign n48166 =  ( n2965 ) ? ( n48163 ) : ( n48165 ) ;
assign n48167 =  ( n1930 ) ? ( n48162 ) : ( n48166 ) ;
assign n48168 =  ( n879 ) ? ( n48157 ) : ( n48167 ) ;
assign n48169 =  ( n172 ) ? ( n9403 ) : ( VREG_4_11 ) ;
assign n48170 =  ( n170 ) ? ( n9402 ) : ( n48169 ) ;
assign n48171 =  ( n168 ) ? ( n9401 ) : ( n48170 ) ;
assign n48172 =  ( n166 ) ? ( n9400 ) : ( n48171 ) ;
assign n48173 =  ( n162 ) ? ( n9399 ) : ( n48172 ) ;
assign n48174 =  ( n172 ) ? ( n9413 ) : ( VREG_4_11 ) ;
assign n48175 =  ( n170 ) ? ( n9412 ) : ( n48174 ) ;
assign n48176 =  ( n168 ) ? ( n9411 ) : ( n48175 ) ;
assign n48177 =  ( n166 ) ? ( n9410 ) : ( n48176 ) ;
assign n48178 =  ( n162 ) ? ( n9409 ) : ( n48177 ) ;
assign n48179 =  ( n9392 ) ? ( VREG_4_11 ) : ( n48178 ) ;
assign n48180 =  ( n3051 ) ? ( n48179 ) : ( VREG_4_11 ) ;
assign n48181 =  ( n3040 ) ? ( n48173 ) : ( n48180 ) ;
assign n48182 =  ( n192 ) ? ( VREG_4_11 ) : ( VREG_4_11 ) ;
assign n48183 =  ( n157 ) ? ( n48181 ) : ( n48182 ) ;
assign n48184 =  ( n6 ) ? ( n48168 ) : ( n48183 ) ;
assign n48185 =  ( n747 ) ? ( n48184 ) : ( VREG_4_11 ) ;
assign n48186 =  ( n148 ) ? ( n10470 ) : ( VREG_4_12 ) ;
assign n48187 =  ( n146 ) ? ( n10469 ) : ( n48186 ) ;
assign n48188 =  ( n144 ) ? ( n10468 ) : ( n48187 ) ;
assign n48189 =  ( n142 ) ? ( n10467 ) : ( n48188 ) ;
assign n48190 =  ( n10 ) ? ( n10466 ) : ( n48189 ) ;
assign n48191 =  ( n148 ) ? ( n11504 ) : ( VREG_4_12 ) ;
assign n48192 =  ( n146 ) ? ( n11503 ) : ( n48191 ) ;
assign n48193 =  ( n144 ) ? ( n11502 ) : ( n48192 ) ;
assign n48194 =  ( n142 ) ? ( n11501 ) : ( n48193 ) ;
assign n48195 =  ( n10 ) ? ( n11500 ) : ( n48194 ) ;
assign n48196 =  ( n11511 ) ? ( VREG_4_12 ) : ( n48190 ) ;
assign n48197 =  ( n11511 ) ? ( VREG_4_12 ) : ( n48195 ) ;
assign n48198 =  ( n3034 ) ? ( n48197 ) : ( VREG_4_12 ) ;
assign n48199 =  ( n2965 ) ? ( n48196 ) : ( n48198 ) ;
assign n48200 =  ( n1930 ) ? ( n48195 ) : ( n48199 ) ;
assign n48201 =  ( n879 ) ? ( n48190 ) : ( n48200 ) ;
assign n48202 =  ( n172 ) ? ( n11522 ) : ( VREG_4_12 ) ;
assign n48203 =  ( n170 ) ? ( n11521 ) : ( n48202 ) ;
assign n48204 =  ( n168 ) ? ( n11520 ) : ( n48203 ) ;
assign n48205 =  ( n166 ) ? ( n11519 ) : ( n48204 ) ;
assign n48206 =  ( n162 ) ? ( n11518 ) : ( n48205 ) ;
assign n48207 =  ( n172 ) ? ( n11532 ) : ( VREG_4_12 ) ;
assign n48208 =  ( n170 ) ? ( n11531 ) : ( n48207 ) ;
assign n48209 =  ( n168 ) ? ( n11530 ) : ( n48208 ) ;
assign n48210 =  ( n166 ) ? ( n11529 ) : ( n48209 ) ;
assign n48211 =  ( n162 ) ? ( n11528 ) : ( n48210 ) ;
assign n48212 =  ( n11511 ) ? ( VREG_4_12 ) : ( n48211 ) ;
assign n48213 =  ( n3051 ) ? ( n48212 ) : ( VREG_4_12 ) ;
assign n48214 =  ( n3040 ) ? ( n48206 ) : ( n48213 ) ;
assign n48215 =  ( n192 ) ? ( VREG_4_12 ) : ( VREG_4_12 ) ;
assign n48216 =  ( n157 ) ? ( n48214 ) : ( n48215 ) ;
assign n48217 =  ( n6 ) ? ( n48201 ) : ( n48216 ) ;
assign n48218 =  ( n747 ) ? ( n48217 ) : ( VREG_4_12 ) ;
assign n48219 =  ( n148 ) ? ( n12589 ) : ( VREG_4_13 ) ;
assign n48220 =  ( n146 ) ? ( n12588 ) : ( n48219 ) ;
assign n48221 =  ( n144 ) ? ( n12587 ) : ( n48220 ) ;
assign n48222 =  ( n142 ) ? ( n12586 ) : ( n48221 ) ;
assign n48223 =  ( n10 ) ? ( n12585 ) : ( n48222 ) ;
assign n48224 =  ( n148 ) ? ( n13623 ) : ( VREG_4_13 ) ;
assign n48225 =  ( n146 ) ? ( n13622 ) : ( n48224 ) ;
assign n48226 =  ( n144 ) ? ( n13621 ) : ( n48225 ) ;
assign n48227 =  ( n142 ) ? ( n13620 ) : ( n48226 ) ;
assign n48228 =  ( n10 ) ? ( n13619 ) : ( n48227 ) ;
assign n48229 =  ( n13630 ) ? ( VREG_4_13 ) : ( n48223 ) ;
assign n48230 =  ( n13630 ) ? ( VREG_4_13 ) : ( n48228 ) ;
assign n48231 =  ( n3034 ) ? ( n48230 ) : ( VREG_4_13 ) ;
assign n48232 =  ( n2965 ) ? ( n48229 ) : ( n48231 ) ;
assign n48233 =  ( n1930 ) ? ( n48228 ) : ( n48232 ) ;
assign n48234 =  ( n879 ) ? ( n48223 ) : ( n48233 ) ;
assign n48235 =  ( n172 ) ? ( n13641 ) : ( VREG_4_13 ) ;
assign n48236 =  ( n170 ) ? ( n13640 ) : ( n48235 ) ;
assign n48237 =  ( n168 ) ? ( n13639 ) : ( n48236 ) ;
assign n48238 =  ( n166 ) ? ( n13638 ) : ( n48237 ) ;
assign n48239 =  ( n162 ) ? ( n13637 ) : ( n48238 ) ;
assign n48240 =  ( n172 ) ? ( n13651 ) : ( VREG_4_13 ) ;
assign n48241 =  ( n170 ) ? ( n13650 ) : ( n48240 ) ;
assign n48242 =  ( n168 ) ? ( n13649 ) : ( n48241 ) ;
assign n48243 =  ( n166 ) ? ( n13648 ) : ( n48242 ) ;
assign n48244 =  ( n162 ) ? ( n13647 ) : ( n48243 ) ;
assign n48245 =  ( n13630 ) ? ( VREG_4_13 ) : ( n48244 ) ;
assign n48246 =  ( n3051 ) ? ( n48245 ) : ( VREG_4_13 ) ;
assign n48247 =  ( n3040 ) ? ( n48239 ) : ( n48246 ) ;
assign n48248 =  ( n192 ) ? ( VREG_4_13 ) : ( VREG_4_13 ) ;
assign n48249 =  ( n157 ) ? ( n48247 ) : ( n48248 ) ;
assign n48250 =  ( n6 ) ? ( n48234 ) : ( n48249 ) ;
assign n48251 =  ( n747 ) ? ( n48250 ) : ( VREG_4_13 ) ;
assign n48252 =  ( n148 ) ? ( n14708 ) : ( VREG_4_14 ) ;
assign n48253 =  ( n146 ) ? ( n14707 ) : ( n48252 ) ;
assign n48254 =  ( n144 ) ? ( n14706 ) : ( n48253 ) ;
assign n48255 =  ( n142 ) ? ( n14705 ) : ( n48254 ) ;
assign n48256 =  ( n10 ) ? ( n14704 ) : ( n48255 ) ;
assign n48257 =  ( n148 ) ? ( n15742 ) : ( VREG_4_14 ) ;
assign n48258 =  ( n146 ) ? ( n15741 ) : ( n48257 ) ;
assign n48259 =  ( n144 ) ? ( n15740 ) : ( n48258 ) ;
assign n48260 =  ( n142 ) ? ( n15739 ) : ( n48259 ) ;
assign n48261 =  ( n10 ) ? ( n15738 ) : ( n48260 ) ;
assign n48262 =  ( n15749 ) ? ( VREG_4_14 ) : ( n48256 ) ;
assign n48263 =  ( n15749 ) ? ( VREG_4_14 ) : ( n48261 ) ;
assign n48264 =  ( n3034 ) ? ( n48263 ) : ( VREG_4_14 ) ;
assign n48265 =  ( n2965 ) ? ( n48262 ) : ( n48264 ) ;
assign n48266 =  ( n1930 ) ? ( n48261 ) : ( n48265 ) ;
assign n48267 =  ( n879 ) ? ( n48256 ) : ( n48266 ) ;
assign n48268 =  ( n172 ) ? ( n15760 ) : ( VREG_4_14 ) ;
assign n48269 =  ( n170 ) ? ( n15759 ) : ( n48268 ) ;
assign n48270 =  ( n168 ) ? ( n15758 ) : ( n48269 ) ;
assign n48271 =  ( n166 ) ? ( n15757 ) : ( n48270 ) ;
assign n48272 =  ( n162 ) ? ( n15756 ) : ( n48271 ) ;
assign n48273 =  ( n172 ) ? ( n15770 ) : ( VREG_4_14 ) ;
assign n48274 =  ( n170 ) ? ( n15769 ) : ( n48273 ) ;
assign n48275 =  ( n168 ) ? ( n15768 ) : ( n48274 ) ;
assign n48276 =  ( n166 ) ? ( n15767 ) : ( n48275 ) ;
assign n48277 =  ( n162 ) ? ( n15766 ) : ( n48276 ) ;
assign n48278 =  ( n15749 ) ? ( VREG_4_14 ) : ( n48277 ) ;
assign n48279 =  ( n3051 ) ? ( n48278 ) : ( VREG_4_14 ) ;
assign n48280 =  ( n3040 ) ? ( n48272 ) : ( n48279 ) ;
assign n48281 =  ( n192 ) ? ( VREG_4_14 ) : ( VREG_4_14 ) ;
assign n48282 =  ( n157 ) ? ( n48280 ) : ( n48281 ) ;
assign n48283 =  ( n6 ) ? ( n48267 ) : ( n48282 ) ;
assign n48284 =  ( n747 ) ? ( n48283 ) : ( VREG_4_14 ) ;
assign n48285 =  ( n148 ) ? ( n16827 ) : ( VREG_4_15 ) ;
assign n48286 =  ( n146 ) ? ( n16826 ) : ( n48285 ) ;
assign n48287 =  ( n144 ) ? ( n16825 ) : ( n48286 ) ;
assign n48288 =  ( n142 ) ? ( n16824 ) : ( n48287 ) ;
assign n48289 =  ( n10 ) ? ( n16823 ) : ( n48288 ) ;
assign n48290 =  ( n148 ) ? ( n17861 ) : ( VREG_4_15 ) ;
assign n48291 =  ( n146 ) ? ( n17860 ) : ( n48290 ) ;
assign n48292 =  ( n144 ) ? ( n17859 ) : ( n48291 ) ;
assign n48293 =  ( n142 ) ? ( n17858 ) : ( n48292 ) ;
assign n48294 =  ( n10 ) ? ( n17857 ) : ( n48293 ) ;
assign n48295 =  ( n17868 ) ? ( VREG_4_15 ) : ( n48289 ) ;
assign n48296 =  ( n17868 ) ? ( VREG_4_15 ) : ( n48294 ) ;
assign n48297 =  ( n3034 ) ? ( n48296 ) : ( VREG_4_15 ) ;
assign n48298 =  ( n2965 ) ? ( n48295 ) : ( n48297 ) ;
assign n48299 =  ( n1930 ) ? ( n48294 ) : ( n48298 ) ;
assign n48300 =  ( n879 ) ? ( n48289 ) : ( n48299 ) ;
assign n48301 =  ( n172 ) ? ( n17879 ) : ( VREG_4_15 ) ;
assign n48302 =  ( n170 ) ? ( n17878 ) : ( n48301 ) ;
assign n48303 =  ( n168 ) ? ( n17877 ) : ( n48302 ) ;
assign n48304 =  ( n166 ) ? ( n17876 ) : ( n48303 ) ;
assign n48305 =  ( n162 ) ? ( n17875 ) : ( n48304 ) ;
assign n48306 =  ( n172 ) ? ( n17889 ) : ( VREG_4_15 ) ;
assign n48307 =  ( n170 ) ? ( n17888 ) : ( n48306 ) ;
assign n48308 =  ( n168 ) ? ( n17887 ) : ( n48307 ) ;
assign n48309 =  ( n166 ) ? ( n17886 ) : ( n48308 ) ;
assign n48310 =  ( n162 ) ? ( n17885 ) : ( n48309 ) ;
assign n48311 =  ( n17868 ) ? ( VREG_4_15 ) : ( n48310 ) ;
assign n48312 =  ( n3051 ) ? ( n48311 ) : ( VREG_4_15 ) ;
assign n48313 =  ( n3040 ) ? ( n48305 ) : ( n48312 ) ;
assign n48314 =  ( n192 ) ? ( VREG_4_15 ) : ( VREG_4_15 ) ;
assign n48315 =  ( n157 ) ? ( n48313 ) : ( n48314 ) ;
assign n48316 =  ( n6 ) ? ( n48300 ) : ( n48315 ) ;
assign n48317 =  ( n747 ) ? ( n48316 ) : ( VREG_4_15 ) ;
assign n48318 =  ( n148 ) ? ( n18946 ) : ( VREG_4_2 ) ;
assign n48319 =  ( n146 ) ? ( n18945 ) : ( n48318 ) ;
assign n48320 =  ( n144 ) ? ( n18944 ) : ( n48319 ) ;
assign n48321 =  ( n142 ) ? ( n18943 ) : ( n48320 ) ;
assign n48322 =  ( n10 ) ? ( n18942 ) : ( n48321 ) ;
assign n48323 =  ( n148 ) ? ( n19980 ) : ( VREG_4_2 ) ;
assign n48324 =  ( n146 ) ? ( n19979 ) : ( n48323 ) ;
assign n48325 =  ( n144 ) ? ( n19978 ) : ( n48324 ) ;
assign n48326 =  ( n142 ) ? ( n19977 ) : ( n48325 ) ;
assign n48327 =  ( n10 ) ? ( n19976 ) : ( n48326 ) ;
assign n48328 =  ( n19987 ) ? ( VREG_4_2 ) : ( n48322 ) ;
assign n48329 =  ( n19987 ) ? ( VREG_4_2 ) : ( n48327 ) ;
assign n48330 =  ( n3034 ) ? ( n48329 ) : ( VREG_4_2 ) ;
assign n48331 =  ( n2965 ) ? ( n48328 ) : ( n48330 ) ;
assign n48332 =  ( n1930 ) ? ( n48327 ) : ( n48331 ) ;
assign n48333 =  ( n879 ) ? ( n48322 ) : ( n48332 ) ;
assign n48334 =  ( n172 ) ? ( n19998 ) : ( VREG_4_2 ) ;
assign n48335 =  ( n170 ) ? ( n19997 ) : ( n48334 ) ;
assign n48336 =  ( n168 ) ? ( n19996 ) : ( n48335 ) ;
assign n48337 =  ( n166 ) ? ( n19995 ) : ( n48336 ) ;
assign n48338 =  ( n162 ) ? ( n19994 ) : ( n48337 ) ;
assign n48339 =  ( n172 ) ? ( n20008 ) : ( VREG_4_2 ) ;
assign n48340 =  ( n170 ) ? ( n20007 ) : ( n48339 ) ;
assign n48341 =  ( n168 ) ? ( n20006 ) : ( n48340 ) ;
assign n48342 =  ( n166 ) ? ( n20005 ) : ( n48341 ) ;
assign n48343 =  ( n162 ) ? ( n20004 ) : ( n48342 ) ;
assign n48344 =  ( n19987 ) ? ( VREG_4_2 ) : ( n48343 ) ;
assign n48345 =  ( n3051 ) ? ( n48344 ) : ( VREG_4_2 ) ;
assign n48346 =  ( n3040 ) ? ( n48338 ) : ( n48345 ) ;
assign n48347 =  ( n192 ) ? ( VREG_4_2 ) : ( VREG_4_2 ) ;
assign n48348 =  ( n157 ) ? ( n48346 ) : ( n48347 ) ;
assign n48349 =  ( n6 ) ? ( n48333 ) : ( n48348 ) ;
assign n48350 =  ( n747 ) ? ( n48349 ) : ( VREG_4_2 ) ;
assign n48351 =  ( n148 ) ? ( n21065 ) : ( VREG_4_3 ) ;
assign n48352 =  ( n146 ) ? ( n21064 ) : ( n48351 ) ;
assign n48353 =  ( n144 ) ? ( n21063 ) : ( n48352 ) ;
assign n48354 =  ( n142 ) ? ( n21062 ) : ( n48353 ) ;
assign n48355 =  ( n10 ) ? ( n21061 ) : ( n48354 ) ;
assign n48356 =  ( n148 ) ? ( n22099 ) : ( VREG_4_3 ) ;
assign n48357 =  ( n146 ) ? ( n22098 ) : ( n48356 ) ;
assign n48358 =  ( n144 ) ? ( n22097 ) : ( n48357 ) ;
assign n48359 =  ( n142 ) ? ( n22096 ) : ( n48358 ) ;
assign n48360 =  ( n10 ) ? ( n22095 ) : ( n48359 ) ;
assign n48361 =  ( n22106 ) ? ( VREG_4_3 ) : ( n48355 ) ;
assign n48362 =  ( n22106 ) ? ( VREG_4_3 ) : ( n48360 ) ;
assign n48363 =  ( n3034 ) ? ( n48362 ) : ( VREG_4_3 ) ;
assign n48364 =  ( n2965 ) ? ( n48361 ) : ( n48363 ) ;
assign n48365 =  ( n1930 ) ? ( n48360 ) : ( n48364 ) ;
assign n48366 =  ( n879 ) ? ( n48355 ) : ( n48365 ) ;
assign n48367 =  ( n172 ) ? ( n22117 ) : ( VREG_4_3 ) ;
assign n48368 =  ( n170 ) ? ( n22116 ) : ( n48367 ) ;
assign n48369 =  ( n168 ) ? ( n22115 ) : ( n48368 ) ;
assign n48370 =  ( n166 ) ? ( n22114 ) : ( n48369 ) ;
assign n48371 =  ( n162 ) ? ( n22113 ) : ( n48370 ) ;
assign n48372 =  ( n172 ) ? ( n22127 ) : ( VREG_4_3 ) ;
assign n48373 =  ( n170 ) ? ( n22126 ) : ( n48372 ) ;
assign n48374 =  ( n168 ) ? ( n22125 ) : ( n48373 ) ;
assign n48375 =  ( n166 ) ? ( n22124 ) : ( n48374 ) ;
assign n48376 =  ( n162 ) ? ( n22123 ) : ( n48375 ) ;
assign n48377 =  ( n22106 ) ? ( VREG_4_3 ) : ( n48376 ) ;
assign n48378 =  ( n3051 ) ? ( n48377 ) : ( VREG_4_3 ) ;
assign n48379 =  ( n3040 ) ? ( n48371 ) : ( n48378 ) ;
assign n48380 =  ( n192 ) ? ( VREG_4_3 ) : ( VREG_4_3 ) ;
assign n48381 =  ( n157 ) ? ( n48379 ) : ( n48380 ) ;
assign n48382 =  ( n6 ) ? ( n48366 ) : ( n48381 ) ;
assign n48383 =  ( n747 ) ? ( n48382 ) : ( VREG_4_3 ) ;
assign n48384 =  ( n148 ) ? ( n23184 ) : ( VREG_4_4 ) ;
assign n48385 =  ( n146 ) ? ( n23183 ) : ( n48384 ) ;
assign n48386 =  ( n144 ) ? ( n23182 ) : ( n48385 ) ;
assign n48387 =  ( n142 ) ? ( n23181 ) : ( n48386 ) ;
assign n48388 =  ( n10 ) ? ( n23180 ) : ( n48387 ) ;
assign n48389 =  ( n148 ) ? ( n24218 ) : ( VREG_4_4 ) ;
assign n48390 =  ( n146 ) ? ( n24217 ) : ( n48389 ) ;
assign n48391 =  ( n144 ) ? ( n24216 ) : ( n48390 ) ;
assign n48392 =  ( n142 ) ? ( n24215 ) : ( n48391 ) ;
assign n48393 =  ( n10 ) ? ( n24214 ) : ( n48392 ) ;
assign n48394 =  ( n24225 ) ? ( VREG_4_4 ) : ( n48388 ) ;
assign n48395 =  ( n24225 ) ? ( VREG_4_4 ) : ( n48393 ) ;
assign n48396 =  ( n3034 ) ? ( n48395 ) : ( VREG_4_4 ) ;
assign n48397 =  ( n2965 ) ? ( n48394 ) : ( n48396 ) ;
assign n48398 =  ( n1930 ) ? ( n48393 ) : ( n48397 ) ;
assign n48399 =  ( n879 ) ? ( n48388 ) : ( n48398 ) ;
assign n48400 =  ( n172 ) ? ( n24236 ) : ( VREG_4_4 ) ;
assign n48401 =  ( n170 ) ? ( n24235 ) : ( n48400 ) ;
assign n48402 =  ( n168 ) ? ( n24234 ) : ( n48401 ) ;
assign n48403 =  ( n166 ) ? ( n24233 ) : ( n48402 ) ;
assign n48404 =  ( n162 ) ? ( n24232 ) : ( n48403 ) ;
assign n48405 =  ( n172 ) ? ( n24246 ) : ( VREG_4_4 ) ;
assign n48406 =  ( n170 ) ? ( n24245 ) : ( n48405 ) ;
assign n48407 =  ( n168 ) ? ( n24244 ) : ( n48406 ) ;
assign n48408 =  ( n166 ) ? ( n24243 ) : ( n48407 ) ;
assign n48409 =  ( n162 ) ? ( n24242 ) : ( n48408 ) ;
assign n48410 =  ( n24225 ) ? ( VREG_4_4 ) : ( n48409 ) ;
assign n48411 =  ( n3051 ) ? ( n48410 ) : ( VREG_4_4 ) ;
assign n48412 =  ( n3040 ) ? ( n48404 ) : ( n48411 ) ;
assign n48413 =  ( n192 ) ? ( VREG_4_4 ) : ( VREG_4_4 ) ;
assign n48414 =  ( n157 ) ? ( n48412 ) : ( n48413 ) ;
assign n48415 =  ( n6 ) ? ( n48399 ) : ( n48414 ) ;
assign n48416 =  ( n747 ) ? ( n48415 ) : ( VREG_4_4 ) ;
assign n48417 =  ( n148 ) ? ( n25303 ) : ( VREG_4_5 ) ;
assign n48418 =  ( n146 ) ? ( n25302 ) : ( n48417 ) ;
assign n48419 =  ( n144 ) ? ( n25301 ) : ( n48418 ) ;
assign n48420 =  ( n142 ) ? ( n25300 ) : ( n48419 ) ;
assign n48421 =  ( n10 ) ? ( n25299 ) : ( n48420 ) ;
assign n48422 =  ( n148 ) ? ( n26337 ) : ( VREG_4_5 ) ;
assign n48423 =  ( n146 ) ? ( n26336 ) : ( n48422 ) ;
assign n48424 =  ( n144 ) ? ( n26335 ) : ( n48423 ) ;
assign n48425 =  ( n142 ) ? ( n26334 ) : ( n48424 ) ;
assign n48426 =  ( n10 ) ? ( n26333 ) : ( n48425 ) ;
assign n48427 =  ( n26344 ) ? ( VREG_4_5 ) : ( n48421 ) ;
assign n48428 =  ( n26344 ) ? ( VREG_4_5 ) : ( n48426 ) ;
assign n48429 =  ( n3034 ) ? ( n48428 ) : ( VREG_4_5 ) ;
assign n48430 =  ( n2965 ) ? ( n48427 ) : ( n48429 ) ;
assign n48431 =  ( n1930 ) ? ( n48426 ) : ( n48430 ) ;
assign n48432 =  ( n879 ) ? ( n48421 ) : ( n48431 ) ;
assign n48433 =  ( n172 ) ? ( n26355 ) : ( VREG_4_5 ) ;
assign n48434 =  ( n170 ) ? ( n26354 ) : ( n48433 ) ;
assign n48435 =  ( n168 ) ? ( n26353 ) : ( n48434 ) ;
assign n48436 =  ( n166 ) ? ( n26352 ) : ( n48435 ) ;
assign n48437 =  ( n162 ) ? ( n26351 ) : ( n48436 ) ;
assign n48438 =  ( n172 ) ? ( n26365 ) : ( VREG_4_5 ) ;
assign n48439 =  ( n170 ) ? ( n26364 ) : ( n48438 ) ;
assign n48440 =  ( n168 ) ? ( n26363 ) : ( n48439 ) ;
assign n48441 =  ( n166 ) ? ( n26362 ) : ( n48440 ) ;
assign n48442 =  ( n162 ) ? ( n26361 ) : ( n48441 ) ;
assign n48443 =  ( n26344 ) ? ( VREG_4_5 ) : ( n48442 ) ;
assign n48444 =  ( n3051 ) ? ( n48443 ) : ( VREG_4_5 ) ;
assign n48445 =  ( n3040 ) ? ( n48437 ) : ( n48444 ) ;
assign n48446 =  ( n192 ) ? ( VREG_4_5 ) : ( VREG_4_5 ) ;
assign n48447 =  ( n157 ) ? ( n48445 ) : ( n48446 ) ;
assign n48448 =  ( n6 ) ? ( n48432 ) : ( n48447 ) ;
assign n48449 =  ( n747 ) ? ( n48448 ) : ( VREG_4_5 ) ;
assign n48450 =  ( n148 ) ? ( n27422 ) : ( VREG_4_6 ) ;
assign n48451 =  ( n146 ) ? ( n27421 ) : ( n48450 ) ;
assign n48452 =  ( n144 ) ? ( n27420 ) : ( n48451 ) ;
assign n48453 =  ( n142 ) ? ( n27419 ) : ( n48452 ) ;
assign n48454 =  ( n10 ) ? ( n27418 ) : ( n48453 ) ;
assign n48455 =  ( n148 ) ? ( n28456 ) : ( VREG_4_6 ) ;
assign n48456 =  ( n146 ) ? ( n28455 ) : ( n48455 ) ;
assign n48457 =  ( n144 ) ? ( n28454 ) : ( n48456 ) ;
assign n48458 =  ( n142 ) ? ( n28453 ) : ( n48457 ) ;
assign n48459 =  ( n10 ) ? ( n28452 ) : ( n48458 ) ;
assign n48460 =  ( n28463 ) ? ( VREG_4_6 ) : ( n48454 ) ;
assign n48461 =  ( n28463 ) ? ( VREG_4_6 ) : ( n48459 ) ;
assign n48462 =  ( n3034 ) ? ( n48461 ) : ( VREG_4_6 ) ;
assign n48463 =  ( n2965 ) ? ( n48460 ) : ( n48462 ) ;
assign n48464 =  ( n1930 ) ? ( n48459 ) : ( n48463 ) ;
assign n48465 =  ( n879 ) ? ( n48454 ) : ( n48464 ) ;
assign n48466 =  ( n172 ) ? ( n28474 ) : ( VREG_4_6 ) ;
assign n48467 =  ( n170 ) ? ( n28473 ) : ( n48466 ) ;
assign n48468 =  ( n168 ) ? ( n28472 ) : ( n48467 ) ;
assign n48469 =  ( n166 ) ? ( n28471 ) : ( n48468 ) ;
assign n48470 =  ( n162 ) ? ( n28470 ) : ( n48469 ) ;
assign n48471 =  ( n172 ) ? ( n28484 ) : ( VREG_4_6 ) ;
assign n48472 =  ( n170 ) ? ( n28483 ) : ( n48471 ) ;
assign n48473 =  ( n168 ) ? ( n28482 ) : ( n48472 ) ;
assign n48474 =  ( n166 ) ? ( n28481 ) : ( n48473 ) ;
assign n48475 =  ( n162 ) ? ( n28480 ) : ( n48474 ) ;
assign n48476 =  ( n28463 ) ? ( VREG_4_6 ) : ( n48475 ) ;
assign n48477 =  ( n3051 ) ? ( n48476 ) : ( VREG_4_6 ) ;
assign n48478 =  ( n3040 ) ? ( n48470 ) : ( n48477 ) ;
assign n48479 =  ( n192 ) ? ( VREG_4_6 ) : ( VREG_4_6 ) ;
assign n48480 =  ( n157 ) ? ( n48478 ) : ( n48479 ) ;
assign n48481 =  ( n6 ) ? ( n48465 ) : ( n48480 ) ;
assign n48482 =  ( n747 ) ? ( n48481 ) : ( VREG_4_6 ) ;
assign n48483 =  ( n148 ) ? ( n29541 ) : ( VREG_4_7 ) ;
assign n48484 =  ( n146 ) ? ( n29540 ) : ( n48483 ) ;
assign n48485 =  ( n144 ) ? ( n29539 ) : ( n48484 ) ;
assign n48486 =  ( n142 ) ? ( n29538 ) : ( n48485 ) ;
assign n48487 =  ( n10 ) ? ( n29537 ) : ( n48486 ) ;
assign n48488 =  ( n148 ) ? ( n30575 ) : ( VREG_4_7 ) ;
assign n48489 =  ( n146 ) ? ( n30574 ) : ( n48488 ) ;
assign n48490 =  ( n144 ) ? ( n30573 ) : ( n48489 ) ;
assign n48491 =  ( n142 ) ? ( n30572 ) : ( n48490 ) ;
assign n48492 =  ( n10 ) ? ( n30571 ) : ( n48491 ) ;
assign n48493 =  ( n30582 ) ? ( VREG_4_7 ) : ( n48487 ) ;
assign n48494 =  ( n30582 ) ? ( VREG_4_7 ) : ( n48492 ) ;
assign n48495 =  ( n3034 ) ? ( n48494 ) : ( VREG_4_7 ) ;
assign n48496 =  ( n2965 ) ? ( n48493 ) : ( n48495 ) ;
assign n48497 =  ( n1930 ) ? ( n48492 ) : ( n48496 ) ;
assign n48498 =  ( n879 ) ? ( n48487 ) : ( n48497 ) ;
assign n48499 =  ( n172 ) ? ( n30593 ) : ( VREG_4_7 ) ;
assign n48500 =  ( n170 ) ? ( n30592 ) : ( n48499 ) ;
assign n48501 =  ( n168 ) ? ( n30591 ) : ( n48500 ) ;
assign n48502 =  ( n166 ) ? ( n30590 ) : ( n48501 ) ;
assign n48503 =  ( n162 ) ? ( n30589 ) : ( n48502 ) ;
assign n48504 =  ( n172 ) ? ( n30603 ) : ( VREG_4_7 ) ;
assign n48505 =  ( n170 ) ? ( n30602 ) : ( n48504 ) ;
assign n48506 =  ( n168 ) ? ( n30601 ) : ( n48505 ) ;
assign n48507 =  ( n166 ) ? ( n30600 ) : ( n48506 ) ;
assign n48508 =  ( n162 ) ? ( n30599 ) : ( n48507 ) ;
assign n48509 =  ( n30582 ) ? ( VREG_4_7 ) : ( n48508 ) ;
assign n48510 =  ( n3051 ) ? ( n48509 ) : ( VREG_4_7 ) ;
assign n48511 =  ( n3040 ) ? ( n48503 ) : ( n48510 ) ;
assign n48512 =  ( n192 ) ? ( VREG_4_7 ) : ( VREG_4_7 ) ;
assign n48513 =  ( n157 ) ? ( n48511 ) : ( n48512 ) ;
assign n48514 =  ( n6 ) ? ( n48498 ) : ( n48513 ) ;
assign n48515 =  ( n747 ) ? ( n48514 ) : ( VREG_4_7 ) ;
assign n48516 =  ( n148 ) ? ( n31660 ) : ( VREG_4_8 ) ;
assign n48517 =  ( n146 ) ? ( n31659 ) : ( n48516 ) ;
assign n48518 =  ( n144 ) ? ( n31658 ) : ( n48517 ) ;
assign n48519 =  ( n142 ) ? ( n31657 ) : ( n48518 ) ;
assign n48520 =  ( n10 ) ? ( n31656 ) : ( n48519 ) ;
assign n48521 =  ( n148 ) ? ( n32694 ) : ( VREG_4_8 ) ;
assign n48522 =  ( n146 ) ? ( n32693 ) : ( n48521 ) ;
assign n48523 =  ( n144 ) ? ( n32692 ) : ( n48522 ) ;
assign n48524 =  ( n142 ) ? ( n32691 ) : ( n48523 ) ;
assign n48525 =  ( n10 ) ? ( n32690 ) : ( n48524 ) ;
assign n48526 =  ( n32701 ) ? ( VREG_4_8 ) : ( n48520 ) ;
assign n48527 =  ( n32701 ) ? ( VREG_4_8 ) : ( n48525 ) ;
assign n48528 =  ( n3034 ) ? ( n48527 ) : ( VREG_4_8 ) ;
assign n48529 =  ( n2965 ) ? ( n48526 ) : ( n48528 ) ;
assign n48530 =  ( n1930 ) ? ( n48525 ) : ( n48529 ) ;
assign n48531 =  ( n879 ) ? ( n48520 ) : ( n48530 ) ;
assign n48532 =  ( n172 ) ? ( n32712 ) : ( VREG_4_8 ) ;
assign n48533 =  ( n170 ) ? ( n32711 ) : ( n48532 ) ;
assign n48534 =  ( n168 ) ? ( n32710 ) : ( n48533 ) ;
assign n48535 =  ( n166 ) ? ( n32709 ) : ( n48534 ) ;
assign n48536 =  ( n162 ) ? ( n32708 ) : ( n48535 ) ;
assign n48537 =  ( n172 ) ? ( n32722 ) : ( VREG_4_8 ) ;
assign n48538 =  ( n170 ) ? ( n32721 ) : ( n48537 ) ;
assign n48539 =  ( n168 ) ? ( n32720 ) : ( n48538 ) ;
assign n48540 =  ( n166 ) ? ( n32719 ) : ( n48539 ) ;
assign n48541 =  ( n162 ) ? ( n32718 ) : ( n48540 ) ;
assign n48542 =  ( n32701 ) ? ( VREG_4_8 ) : ( n48541 ) ;
assign n48543 =  ( n3051 ) ? ( n48542 ) : ( VREG_4_8 ) ;
assign n48544 =  ( n3040 ) ? ( n48536 ) : ( n48543 ) ;
assign n48545 =  ( n192 ) ? ( VREG_4_8 ) : ( VREG_4_8 ) ;
assign n48546 =  ( n157 ) ? ( n48544 ) : ( n48545 ) ;
assign n48547 =  ( n6 ) ? ( n48531 ) : ( n48546 ) ;
assign n48548 =  ( n747 ) ? ( n48547 ) : ( VREG_4_8 ) ;
assign n48549 =  ( n148 ) ? ( n33779 ) : ( VREG_4_9 ) ;
assign n48550 =  ( n146 ) ? ( n33778 ) : ( n48549 ) ;
assign n48551 =  ( n144 ) ? ( n33777 ) : ( n48550 ) ;
assign n48552 =  ( n142 ) ? ( n33776 ) : ( n48551 ) ;
assign n48553 =  ( n10 ) ? ( n33775 ) : ( n48552 ) ;
assign n48554 =  ( n148 ) ? ( n34813 ) : ( VREG_4_9 ) ;
assign n48555 =  ( n146 ) ? ( n34812 ) : ( n48554 ) ;
assign n48556 =  ( n144 ) ? ( n34811 ) : ( n48555 ) ;
assign n48557 =  ( n142 ) ? ( n34810 ) : ( n48556 ) ;
assign n48558 =  ( n10 ) ? ( n34809 ) : ( n48557 ) ;
assign n48559 =  ( n34820 ) ? ( VREG_4_9 ) : ( n48553 ) ;
assign n48560 =  ( n34820 ) ? ( VREG_4_9 ) : ( n48558 ) ;
assign n48561 =  ( n3034 ) ? ( n48560 ) : ( VREG_4_9 ) ;
assign n48562 =  ( n2965 ) ? ( n48559 ) : ( n48561 ) ;
assign n48563 =  ( n1930 ) ? ( n48558 ) : ( n48562 ) ;
assign n48564 =  ( n879 ) ? ( n48553 ) : ( n48563 ) ;
assign n48565 =  ( n172 ) ? ( n34831 ) : ( VREG_4_9 ) ;
assign n48566 =  ( n170 ) ? ( n34830 ) : ( n48565 ) ;
assign n48567 =  ( n168 ) ? ( n34829 ) : ( n48566 ) ;
assign n48568 =  ( n166 ) ? ( n34828 ) : ( n48567 ) ;
assign n48569 =  ( n162 ) ? ( n34827 ) : ( n48568 ) ;
assign n48570 =  ( n172 ) ? ( n34841 ) : ( VREG_4_9 ) ;
assign n48571 =  ( n170 ) ? ( n34840 ) : ( n48570 ) ;
assign n48572 =  ( n168 ) ? ( n34839 ) : ( n48571 ) ;
assign n48573 =  ( n166 ) ? ( n34838 ) : ( n48572 ) ;
assign n48574 =  ( n162 ) ? ( n34837 ) : ( n48573 ) ;
assign n48575 =  ( n34820 ) ? ( VREG_4_9 ) : ( n48574 ) ;
assign n48576 =  ( n3051 ) ? ( n48575 ) : ( VREG_4_9 ) ;
assign n48577 =  ( n3040 ) ? ( n48569 ) : ( n48576 ) ;
assign n48578 =  ( n192 ) ? ( VREG_4_9 ) : ( VREG_4_9 ) ;
assign n48579 =  ( n157 ) ? ( n48577 ) : ( n48578 ) ;
assign n48580 =  ( n6 ) ? ( n48564 ) : ( n48579 ) ;
assign n48581 =  ( n747 ) ? ( n48580 ) : ( VREG_4_9 ) ;
assign n48582 =  ( n148 ) ? ( n1924 ) : ( VREG_5_0 ) ;
assign n48583 =  ( n146 ) ? ( n1923 ) : ( n48582 ) ;
assign n48584 =  ( n144 ) ? ( n1922 ) : ( n48583 ) ;
assign n48585 =  ( n142 ) ? ( n1921 ) : ( n48584 ) ;
assign n48586 =  ( n10 ) ? ( n1920 ) : ( n48585 ) ;
assign n48587 =  ( n148 ) ? ( n2959 ) : ( VREG_5_0 ) ;
assign n48588 =  ( n146 ) ? ( n2958 ) : ( n48587 ) ;
assign n48589 =  ( n144 ) ? ( n2957 ) : ( n48588 ) ;
assign n48590 =  ( n142 ) ? ( n2956 ) : ( n48589 ) ;
assign n48591 =  ( n10 ) ? ( n2955 ) : ( n48590 ) ;
assign n48592 =  ( n3032 ) ? ( VREG_5_0 ) : ( n48586 ) ;
assign n48593 =  ( n3032 ) ? ( VREG_5_0 ) : ( n48591 ) ;
assign n48594 =  ( n3034 ) ? ( n48593 ) : ( VREG_5_0 ) ;
assign n48595 =  ( n2965 ) ? ( n48592 ) : ( n48594 ) ;
assign n48596 =  ( n1930 ) ? ( n48591 ) : ( n48595 ) ;
assign n48597 =  ( n879 ) ? ( n48586 ) : ( n48596 ) ;
assign n48598 =  ( n172 ) ? ( n3045 ) : ( VREG_5_0 ) ;
assign n48599 =  ( n170 ) ? ( n3044 ) : ( n48598 ) ;
assign n48600 =  ( n168 ) ? ( n3043 ) : ( n48599 ) ;
assign n48601 =  ( n166 ) ? ( n3042 ) : ( n48600 ) ;
assign n48602 =  ( n162 ) ? ( n3041 ) : ( n48601 ) ;
assign n48603 =  ( n172 ) ? ( n3056 ) : ( VREG_5_0 ) ;
assign n48604 =  ( n170 ) ? ( n3055 ) : ( n48603 ) ;
assign n48605 =  ( n168 ) ? ( n3054 ) : ( n48604 ) ;
assign n48606 =  ( n166 ) ? ( n3053 ) : ( n48605 ) ;
assign n48607 =  ( n162 ) ? ( n3052 ) : ( n48606 ) ;
assign n48608 =  ( n3032 ) ? ( VREG_5_0 ) : ( n48607 ) ;
assign n48609 =  ( n3051 ) ? ( n48608 ) : ( VREG_5_0 ) ;
assign n48610 =  ( n3040 ) ? ( n48602 ) : ( n48609 ) ;
assign n48611 =  ( n192 ) ? ( VREG_5_0 ) : ( VREG_5_0 ) ;
assign n48612 =  ( n157 ) ? ( n48610 ) : ( n48611 ) ;
assign n48613 =  ( n6 ) ? ( n48597 ) : ( n48612 ) ;
assign n48614 =  ( n769 ) ? ( n48613 ) : ( VREG_5_0 ) ;
assign n48615 =  ( n148 ) ? ( n4113 ) : ( VREG_5_1 ) ;
assign n48616 =  ( n146 ) ? ( n4112 ) : ( n48615 ) ;
assign n48617 =  ( n144 ) ? ( n4111 ) : ( n48616 ) ;
assign n48618 =  ( n142 ) ? ( n4110 ) : ( n48617 ) ;
assign n48619 =  ( n10 ) ? ( n4109 ) : ( n48618 ) ;
assign n48620 =  ( n148 ) ? ( n5147 ) : ( VREG_5_1 ) ;
assign n48621 =  ( n146 ) ? ( n5146 ) : ( n48620 ) ;
assign n48622 =  ( n144 ) ? ( n5145 ) : ( n48621 ) ;
assign n48623 =  ( n142 ) ? ( n5144 ) : ( n48622 ) ;
assign n48624 =  ( n10 ) ? ( n5143 ) : ( n48623 ) ;
assign n48625 =  ( n5154 ) ? ( VREG_5_1 ) : ( n48619 ) ;
assign n48626 =  ( n5154 ) ? ( VREG_5_1 ) : ( n48624 ) ;
assign n48627 =  ( n3034 ) ? ( n48626 ) : ( VREG_5_1 ) ;
assign n48628 =  ( n2965 ) ? ( n48625 ) : ( n48627 ) ;
assign n48629 =  ( n1930 ) ? ( n48624 ) : ( n48628 ) ;
assign n48630 =  ( n879 ) ? ( n48619 ) : ( n48629 ) ;
assign n48631 =  ( n172 ) ? ( n5165 ) : ( VREG_5_1 ) ;
assign n48632 =  ( n170 ) ? ( n5164 ) : ( n48631 ) ;
assign n48633 =  ( n168 ) ? ( n5163 ) : ( n48632 ) ;
assign n48634 =  ( n166 ) ? ( n5162 ) : ( n48633 ) ;
assign n48635 =  ( n162 ) ? ( n5161 ) : ( n48634 ) ;
assign n48636 =  ( n172 ) ? ( n5175 ) : ( VREG_5_1 ) ;
assign n48637 =  ( n170 ) ? ( n5174 ) : ( n48636 ) ;
assign n48638 =  ( n168 ) ? ( n5173 ) : ( n48637 ) ;
assign n48639 =  ( n166 ) ? ( n5172 ) : ( n48638 ) ;
assign n48640 =  ( n162 ) ? ( n5171 ) : ( n48639 ) ;
assign n48641 =  ( n5154 ) ? ( VREG_5_1 ) : ( n48640 ) ;
assign n48642 =  ( n3051 ) ? ( n48641 ) : ( VREG_5_1 ) ;
assign n48643 =  ( n3040 ) ? ( n48635 ) : ( n48642 ) ;
assign n48644 =  ( n192 ) ? ( VREG_5_1 ) : ( VREG_5_1 ) ;
assign n48645 =  ( n157 ) ? ( n48643 ) : ( n48644 ) ;
assign n48646 =  ( n6 ) ? ( n48630 ) : ( n48645 ) ;
assign n48647 =  ( n769 ) ? ( n48646 ) : ( VREG_5_1 ) ;
assign n48648 =  ( n148 ) ? ( n6232 ) : ( VREG_5_10 ) ;
assign n48649 =  ( n146 ) ? ( n6231 ) : ( n48648 ) ;
assign n48650 =  ( n144 ) ? ( n6230 ) : ( n48649 ) ;
assign n48651 =  ( n142 ) ? ( n6229 ) : ( n48650 ) ;
assign n48652 =  ( n10 ) ? ( n6228 ) : ( n48651 ) ;
assign n48653 =  ( n148 ) ? ( n7266 ) : ( VREG_5_10 ) ;
assign n48654 =  ( n146 ) ? ( n7265 ) : ( n48653 ) ;
assign n48655 =  ( n144 ) ? ( n7264 ) : ( n48654 ) ;
assign n48656 =  ( n142 ) ? ( n7263 ) : ( n48655 ) ;
assign n48657 =  ( n10 ) ? ( n7262 ) : ( n48656 ) ;
assign n48658 =  ( n7273 ) ? ( VREG_5_10 ) : ( n48652 ) ;
assign n48659 =  ( n7273 ) ? ( VREG_5_10 ) : ( n48657 ) ;
assign n48660 =  ( n3034 ) ? ( n48659 ) : ( VREG_5_10 ) ;
assign n48661 =  ( n2965 ) ? ( n48658 ) : ( n48660 ) ;
assign n48662 =  ( n1930 ) ? ( n48657 ) : ( n48661 ) ;
assign n48663 =  ( n879 ) ? ( n48652 ) : ( n48662 ) ;
assign n48664 =  ( n172 ) ? ( n7284 ) : ( VREG_5_10 ) ;
assign n48665 =  ( n170 ) ? ( n7283 ) : ( n48664 ) ;
assign n48666 =  ( n168 ) ? ( n7282 ) : ( n48665 ) ;
assign n48667 =  ( n166 ) ? ( n7281 ) : ( n48666 ) ;
assign n48668 =  ( n162 ) ? ( n7280 ) : ( n48667 ) ;
assign n48669 =  ( n172 ) ? ( n7294 ) : ( VREG_5_10 ) ;
assign n48670 =  ( n170 ) ? ( n7293 ) : ( n48669 ) ;
assign n48671 =  ( n168 ) ? ( n7292 ) : ( n48670 ) ;
assign n48672 =  ( n166 ) ? ( n7291 ) : ( n48671 ) ;
assign n48673 =  ( n162 ) ? ( n7290 ) : ( n48672 ) ;
assign n48674 =  ( n7273 ) ? ( VREG_5_10 ) : ( n48673 ) ;
assign n48675 =  ( n3051 ) ? ( n48674 ) : ( VREG_5_10 ) ;
assign n48676 =  ( n3040 ) ? ( n48668 ) : ( n48675 ) ;
assign n48677 =  ( n192 ) ? ( VREG_5_10 ) : ( VREG_5_10 ) ;
assign n48678 =  ( n157 ) ? ( n48676 ) : ( n48677 ) ;
assign n48679 =  ( n6 ) ? ( n48663 ) : ( n48678 ) ;
assign n48680 =  ( n769 ) ? ( n48679 ) : ( VREG_5_10 ) ;
assign n48681 =  ( n148 ) ? ( n8351 ) : ( VREG_5_11 ) ;
assign n48682 =  ( n146 ) ? ( n8350 ) : ( n48681 ) ;
assign n48683 =  ( n144 ) ? ( n8349 ) : ( n48682 ) ;
assign n48684 =  ( n142 ) ? ( n8348 ) : ( n48683 ) ;
assign n48685 =  ( n10 ) ? ( n8347 ) : ( n48684 ) ;
assign n48686 =  ( n148 ) ? ( n9385 ) : ( VREG_5_11 ) ;
assign n48687 =  ( n146 ) ? ( n9384 ) : ( n48686 ) ;
assign n48688 =  ( n144 ) ? ( n9383 ) : ( n48687 ) ;
assign n48689 =  ( n142 ) ? ( n9382 ) : ( n48688 ) ;
assign n48690 =  ( n10 ) ? ( n9381 ) : ( n48689 ) ;
assign n48691 =  ( n9392 ) ? ( VREG_5_11 ) : ( n48685 ) ;
assign n48692 =  ( n9392 ) ? ( VREG_5_11 ) : ( n48690 ) ;
assign n48693 =  ( n3034 ) ? ( n48692 ) : ( VREG_5_11 ) ;
assign n48694 =  ( n2965 ) ? ( n48691 ) : ( n48693 ) ;
assign n48695 =  ( n1930 ) ? ( n48690 ) : ( n48694 ) ;
assign n48696 =  ( n879 ) ? ( n48685 ) : ( n48695 ) ;
assign n48697 =  ( n172 ) ? ( n9403 ) : ( VREG_5_11 ) ;
assign n48698 =  ( n170 ) ? ( n9402 ) : ( n48697 ) ;
assign n48699 =  ( n168 ) ? ( n9401 ) : ( n48698 ) ;
assign n48700 =  ( n166 ) ? ( n9400 ) : ( n48699 ) ;
assign n48701 =  ( n162 ) ? ( n9399 ) : ( n48700 ) ;
assign n48702 =  ( n172 ) ? ( n9413 ) : ( VREG_5_11 ) ;
assign n48703 =  ( n170 ) ? ( n9412 ) : ( n48702 ) ;
assign n48704 =  ( n168 ) ? ( n9411 ) : ( n48703 ) ;
assign n48705 =  ( n166 ) ? ( n9410 ) : ( n48704 ) ;
assign n48706 =  ( n162 ) ? ( n9409 ) : ( n48705 ) ;
assign n48707 =  ( n9392 ) ? ( VREG_5_11 ) : ( n48706 ) ;
assign n48708 =  ( n3051 ) ? ( n48707 ) : ( VREG_5_11 ) ;
assign n48709 =  ( n3040 ) ? ( n48701 ) : ( n48708 ) ;
assign n48710 =  ( n192 ) ? ( VREG_5_11 ) : ( VREG_5_11 ) ;
assign n48711 =  ( n157 ) ? ( n48709 ) : ( n48710 ) ;
assign n48712 =  ( n6 ) ? ( n48696 ) : ( n48711 ) ;
assign n48713 =  ( n769 ) ? ( n48712 ) : ( VREG_5_11 ) ;
assign n48714 =  ( n148 ) ? ( n10470 ) : ( VREG_5_12 ) ;
assign n48715 =  ( n146 ) ? ( n10469 ) : ( n48714 ) ;
assign n48716 =  ( n144 ) ? ( n10468 ) : ( n48715 ) ;
assign n48717 =  ( n142 ) ? ( n10467 ) : ( n48716 ) ;
assign n48718 =  ( n10 ) ? ( n10466 ) : ( n48717 ) ;
assign n48719 =  ( n148 ) ? ( n11504 ) : ( VREG_5_12 ) ;
assign n48720 =  ( n146 ) ? ( n11503 ) : ( n48719 ) ;
assign n48721 =  ( n144 ) ? ( n11502 ) : ( n48720 ) ;
assign n48722 =  ( n142 ) ? ( n11501 ) : ( n48721 ) ;
assign n48723 =  ( n10 ) ? ( n11500 ) : ( n48722 ) ;
assign n48724 =  ( n11511 ) ? ( VREG_5_12 ) : ( n48718 ) ;
assign n48725 =  ( n11511 ) ? ( VREG_5_12 ) : ( n48723 ) ;
assign n48726 =  ( n3034 ) ? ( n48725 ) : ( VREG_5_12 ) ;
assign n48727 =  ( n2965 ) ? ( n48724 ) : ( n48726 ) ;
assign n48728 =  ( n1930 ) ? ( n48723 ) : ( n48727 ) ;
assign n48729 =  ( n879 ) ? ( n48718 ) : ( n48728 ) ;
assign n48730 =  ( n172 ) ? ( n11522 ) : ( VREG_5_12 ) ;
assign n48731 =  ( n170 ) ? ( n11521 ) : ( n48730 ) ;
assign n48732 =  ( n168 ) ? ( n11520 ) : ( n48731 ) ;
assign n48733 =  ( n166 ) ? ( n11519 ) : ( n48732 ) ;
assign n48734 =  ( n162 ) ? ( n11518 ) : ( n48733 ) ;
assign n48735 =  ( n172 ) ? ( n11532 ) : ( VREG_5_12 ) ;
assign n48736 =  ( n170 ) ? ( n11531 ) : ( n48735 ) ;
assign n48737 =  ( n168 ) ? ( n11530 ) : ( n48736 ) ;
assign n48738 =  ( n166 ) ? ( n11529 ) : ( n48737 ) ;
assign n48739 =  ( n162 ) ? ( n11528 ) : ( n48738 ) ;
assign n48740 =  ( n11511 ) ? ( VREG_5_12 ) : ( n48739 ) ;
assign n48741 =  ( n3051 ) ? ( n48740 ) : ( VREG_5_12 ) ;
assign n48742 =  ( n3040 ) ? ( n48734 ) : ( n48741 ) ;
assign n48743 =  ( n192 ) ? ( VREG_5_12 ) : ( VREG_5_12 ) ;
assign n48744 =  ( n157 ) ? ( n48742 ) : ( n48743 ) ;
assign n48745 =  ( n6 ) ? ( n48729 ) : ( n48744 ) ;
assign n48746 =  ( n769 ) ? ( n48745 ) : ( VREG_5_12 ) ;
assign n48747 =  ( n148 ) ? ( n12589 ) : ( VREG_5_13 ) ;
assign n48748 =  ( n146 ) ? ( n12588 ) : ( n48747 ) ;
assign n48749 =  ( n144 ) ? ( n12587 ) : ( n48748 ) ;
assign n48750 =  ( n142 ) ? ( n12586 ) : ( n48749 ) ;
assign n48751 =  ( n10 ) ? ( n12585 ) : ( n48750 ) ;
assign n48752 =  ( n148 ) ? ( n13623 ) : ( VREG_5_13 ) ;
assign n48753 =  ( n146 ) ? ( n13622 ) : ( n48752 ) ;
assign n48754 =  ( n144 ) ? ( n13621 ) : ( n48753 ) ;
assign n48755 =  ( n142 ) ? ( n13620 ) : ( n48754 ) ;
assign n48756 =  ( n10 ) ? ( n13619 ) : ( n48755 ) ;
assign n48757 =  ( n13630 ) ? ( VREG_5_13 ) : ( n48751 ) ;
assign n48758 =  ( n13630 ) ? ( VREG_5_13 ) : ( n48756 ) ;
assign n48759 =  ( n3034 ) ? ( n48758 ) : ( VREG_5_13 ) ;
assign n48760 =  ( n2965 ) ? ( n48757 ) : ( n48759 ) ;
assign n48761 =  ( n1930 ) ? ( n48756 ) : ( n48760 ) ;
assign n48762 =  ( n879 ) ? ( n48751 ) : ( n48761 ) ;
assign n48763 =  ( n172 ) ? ( n13641 ) : ( VREG_5_13 ) ;
assign n48764 =  ( n170 ) ? ( n13640 ) : ( n48763 ) ;
assign n48765 =  ( n168 ) ? ( n13639 ) : ( n48764 ) ;
assign n48766 =  ( n166 ) ? ( n13638 ) : ( n48765 ) ;
assign n48767 =  ( n162 ) ? ( n13637 ) : ( n48766 ) ;
assign n48768 =  ( n172 ) ? ( n13651 ) : ( VREG_5_13 ) ;
assign n48769 =  ( n170 ) ? ( n13650 ) : ( n48768 ) ;
assign n48770 =  ( n168 ) ? ( n13649 ) : ( n48769 ) ;
assign n48771 =  ( n166 ) ? ( n13648 ) : ( n48770 ) ;
assign n48772 =  ( n162 ) ? ( n13647 ) : ( n48771 ) ;
assign n48773 =  ( n13630 ) ? ( VREG_5_13 ) : ( n48772 ) ;
assign n48774 =  ( n3051 ) ? ( n48773 ) : ( VREG_5_13 ) ;
assign n48775 =  ( n3040 ) ? ( n48767 ) : ( n48774 ) ;
assign n48776 =  ( n192 ) ? ( VREG_5_13 ) : ( VREG_5_13 ) ;
assign n48777 =  ( n157 ) ? ( n48775 ) : ( n48776 ) ;
assign n48778 =  ( n6 ) ? ( n48762 ) : ( n48777 ) ;
assign n48779 =  ( n769 ) ? ( n48778 ) : ( VREG_5_13 ) ;
assign n48780 =  ( n148 ) ? ( n14708 ) : ( VREG_5_14 ) ;
assign n48781 =  ( n146 ) ? ( n14707 ) : ( n48780 ) ;
assign n48782 =  ( n144 ) ? ( n14706 ) : ( n48781 ) ;
assign n48783 =  ( n142 ) ? ( n14705 ) : ( n48782 ) ;
assign n48784 =  ( n10 ) ? ( n14704 ) : ( n48783 ) ;
assign n48785 =  ( n148 ) ? ( n15742 ) : ( VREG_5_14 ) ;
assign n48786 =  ( n146 ) ? ( n15741 ) : ( n48785 ) ;
assign n48787 =  ( n144 ) ? ( n15740 ) : ( n48786 ) ;
assign n48788 =  ( n142 ) ? ( n15739 ) : ( n48787 ) ;
assign n48789 =  ( n10 ) ? ( n15738 ) : ( n48788 ) ;
assign n48790 =  ( n15749 ) ? ( VREG_5_14 ) : ( n48784 ) ;
assign n48791 =  ( n15749 ) ? ( VREG_5_14 ) : ( n48789 ) ;
assign n48792 =  ( n3034 ) ? ( n48791 ) : ( VREG_5_14 ) ;
assign n48793 =  ( n2965 ) ? ( n48790 ) : ( n48792 ) ;
assign n48794 =  ( n1930 ) ? ( n48789 ) : ( n48793 ) ;
assign n48795 =  ( n879 ) ? ( n48784 ) : ( n48794 ) ;
assign n48796 =  ( n172 ) ? ( n15760 ) : ( VREG_5_14 ) ;
assign n48797 =  ( n170 ) ? ( n15759 ) : ( n48796 ) ;
assign n48798 =  ( n168 ) ? ( n15758 ) : ( n48797 ) ;
assign n48799 =  ( n166 ) ? ( n15757 ) : ( n48798 ) ;
assign n48800 =  ( n162 ) ? ( n15756 ) : ( n48799 ) ;
assign n48801 =  ( n172 ) ? ( n15770 ) : ( VREG_5_14 ) ;
assign n48802 =  ( n170 ) ? ( n15769 ) : ( n48801 ) ;
assign n48803 =  ( n168 ) ? ( n15768 ) : ( n48802 ) ;
assign n48804 =  ( n166 ) ? ( n15767 ) : ( n48803 ) ;
assign n48805 =  ( n162 ) ? ( n15766 ) : ( n48804 ) ;
assign n48806 =  ( n15749 ) ? ( VREG_5_14 ) : ( n48805 ) ;
assign n48807 =  ( n3051 ) ? ( n48806 ) : ( VREG_5_14 ) ;
assign n48808 =  ( n3040 ) ? ( n48800 ) : ( n48807 ) ;
assign n48809 =  ( n192 ) ? ( VREG_5_14 ) : ( VREG_5_14 ) ;
assign n48810 =  ( n157 ) ? ( n48808 ) : ( n48809 ) ;
assign n48811 =  ( n6 ) ? ( n48795 ) : ( n48810 ) ;
assign n48812 =  ( n769 ) ? ( n48811 ) : ( VREG_5_14 ) ;
assign n48813 =  ( n148 ) ? ( n16827 ) : ( VREG_5_15 ) ;
assign n48814 =  ( n146 ) ? ( n16826 ) : ( n48813 ) ;
assign n48815 =  ( n144 ) ? ( n16825 ) : ( n48814 ) ;
assign n48816 =  ( n142 ) ? ( n16824 ) : ( n48815 ) ;
assign n48817 =  ( n10 ) ? ( n16823 ) : ( n48816 ) ;
assign n48818 =  ( n148 ) ? ( n17861 ) : ( VREG_5_15 ) ;
assign n48819 =  ( n146 ) ? ( n17860 ) : ( n48818 ) ;
assign n48820 =  ( n144 ) ? ( n17859 ) : ( n48819 ) ;
assign n48821 =  ( n142 ) ? ( n17858 ) : ( n48820 ) ;
assign n48822 =  ( n10 ) ? ( n17857 ) : ( n48821 ) ;
assign n48823 =  ( n17868 ) ? ( VREG_5_15 ) : ( n48817 ) ;
assign n48824 =  ( n17868 ) ? ( VREG_5_15 ) : ( n48822 ) ;
assign n48825 =  ( n3034 ) ? ( n48824 ) : ( VREG_5_15 ) ;
assign n48826 =  ( n2965 ) ? ( n48823 ) : ( n48825 ) ;
assign n48827 =  ( n1930 ) ? ( n48822 ) : ( n48826 ) ;
assign n48828 =  ( n879 ) ? ( n48817 ) : ( n48827 ) ;
assign n48829 =  ( n172 ) ? ( n17879 ) : ( VREG_5_15 ) ;
assign n48830 =  ( n170 ) ? ( n17878 ) : ( n48829 ) ;
assign n48831 =  ( n168 ) ? ( n17877 ) : ( n48830 ) ;
assign n48832 =  ( n166 ) ? ( n17876 ) : ( n48831 ) ;
assign n48833 =  ( n162 ) ? ( n17875 ) : ( n48832 ) ;
assign n48834 =  ( n172 ) ? ( n17889 ) : ( VREG_5_15 ) ;
assign n48835 =  ( n170 ) ? ( n17888 ) : ( n48834 ) ;
assign n48836 =  ( n168 ) ? ( n17887 ) : ( n48835 ) ;
assign n48837 =  ( n166 ) ? ( n17886 ) : ( n48836 ) ;
assign n48838 =  ( n162 ) ? ( n17885 ) : ( n48837 ) ;
assign n48839 =  ( n17868 ) ? ( VREG_5_15 ) : ( n48838 ) ;
assign n48840 =  ( n3051 ) ? ( n48839 ) : ( VREG_5_15 ) ;
assign n48841 =  ( n3040 ) ? ( n48833 ) : ( n48840 ) ;
assign n48842 =  ( n192 ) ? ( VREG_5_15 ) : ( VREG_5_15 ) ;
assign n48843 =  ( n157 ) ? ( n48841 ) : ( n48842 ) ;
assign n48844 =  ( n6 ) ? ( n48828 ) : ( n48843 ) ;
assign n48845 =  ( n769 ) ? ( n48844 ) : ( VREG_5_15 ) ;
assign n48846 =  ( n148 ) ? ( n18946 ) : ( VREG_5_2 ) ;
assign n48847 =  ( n146 ) ? ( n18945 ) : ( n48846 ) ;
assign n48848 =  ( n144 ) ? ( n18944 ) : ( n48847 ) ;
assign n48849 =  ( n142 ) ? ( n18943 ) : ( n48848 ) ;
assign n48850 =  ( n10 ) ? ( n18942 ) : ( n48849 ) ;
assign n48851 =  ( n148 ) ? ( n19980 ) : ( VREG_5_2 ) ;
assign n48852 =  ( n146 ) ? ( n19979 ) : ( n48851 ) ;
assign n48853 =  ( n144 ) ? ( n19978 ) : ( n48852 ) ;
assign n48854 =  ( n142 ) ? ( n19977 ) : ( n48853 ) ;
assign n48855 =  ( n10 ) ? ( n19976 ) : ( n48854 ) ;
assign n48856 =  ( n19987 ) ? ( VREG_5_2 ) : ( n48850 ) ;
assign n48857 =  ( n19987 ) ? ( VREG_5_2 ) : ( n48855 ) ;
assign n48858 =  ( n3034 ) ? ( n48857 ) : ( VREG_5_2 ) ;
assign n48859 =  ( n2965 ) ? ( n48856 ) : ( n48858 ) ;
assign n48860 =  ( n1930 ) ? ( n48855 ) : ( n48859 ) ;
assign n48861 =  ( n879 ) ? ( n48850 ) : ( n48860 ) ;
assign n48862 =  ( n172 ) ? ( n19998 ) : ( VREG_5_2 ) ;
assign n48863 =  ( n170 ) ? ( n19997 ) : ( n48862 ) ;
assign n48864 =  ( n168 ) ? ( n19996 ) : ( n48863 ) ;
assign n48865 =  ( n166 ) ? ( n19995 ) : ( n48864 ) ;
assign n48866 =  ( n162 ) ? ( n19994 ) : ( n48865 ) ;
assign n48867 =  ( n172 ) ? ( n20008 ) : ( VREG_5_2 ) ;
assign n48868 =  ( n170 ) ? ( n20007 ) : ( n48867 ) ;
assign n48869 =  ( n168 ) ? ( n20006 ) : ( n48868 ) ;
assign n48870 =  ( n166 ) ? ( n20005 ) : ( n48869 ) ;
assign n48871 =  ( n162 ) ? ( n20004 ) : ( n48870 ) ;
assign n48872 =  ( n19987 ) ? ( VREG_5_2 ) : ( n48871 ) ;
assign n48873 =  ( n3051 ) ? ( n48872 ) : ( VREG_5_2 ) ;
assign n48874 =  ( n3040 ) ? ( n48866 ) : ( n48873 ) ;
assign n48875 =  ( n192 ) ? ( VREG_5_2 ) : ( VREG_5_2 ) ;
assign n48876 =  ( n157 ) ? ( n48874 ) : ( n48875 ) ;
assign n48877 =  ( n6 ) ? ( n48861 ) : ( n48876 ) ;
assign n48878 =  ( n769 ) ? ( n48877 ) : ( VREG_5_2 ) ;
assign n48879 =  ( n148 ) ? ( n21065 ) : ( VREG_5_3 ) ;
assign n48880 =  ( n146 ) ? ( n21064 ) : ( n48879 ) ;
assign n48881 =  ( n144 ) ? ( n21063 ) : ( n48880 ) ;
assign n48882 =  ( n142 ) ? ( n21062 ) : ( n48881 ) ;
assign n48883 =  ( n10 ) ? ( n21061 ) : ( n48882 ) ;
assign n48884 =  ( n148 ) ? ( n22099 ) : ( VREG_5_3 ) ;
assign n48885 =  ( n146 ) ? ( n22098 ) : ( n48884 ) ;
assign n48886 =  ( n144 ) ? ( n22097 ) : ( n48885 ) ;
assign n48887 =  ( n142 ) ? ( n22096 ) : ( n48886 ) ;
assign n48888 =  ( n10 ) ? ( n22095 ) : ( n48887 ) ;
assign n48889 =  ( n22106 ) ? ( VREG_5_3 ) : ( n48883 ) ;
assign n48890 =  ( n22106 ) ? ( VREG_5_3 ) : ( n48888 ) ;
assign n48891 =  ( n3034 ) ? ( n48890 ) : ( VREG_5_3 ) ;
assign n48892 =  ( n2965 ) ? ( n48889 ) : ( n48891 ) ;
assign n48893 =  ( n1930 ) ? ( n48888 ) : ( n48892 ) ;
assign n48894 =  ( n879 ) ? ( n48883 ) : ( n48893 ) ;
assign n48895 =  ( n172 ) ? ( n22117 ) : ( VREG_5_3 ) ;
assign n48896 =  ( n170 ) ? ( n22116 ) : ( n48895 ) ;
assign n48897 =  ( n168 ) ? ( n22115 ) : ( n48896 ) ;
assign n48898 =  ( n166 ) ? ( n22114 ) : ( n48897 ) ;
assign n48899 =  ( n162 ) ? ( n22113 ) : ( n48898 ) ;
assign n48900 =  ( n172 ) ? ( n22127 ) : ( VREG_5_3 ) ;
assign n48901 =  ( n170 ) ? ( n22126 ) : ( n48900 ) ;
assign n48902 =  ( n168 ) ? ( n22125 ) : ( n48901 ) ;
assign n48903 =  ( n166 ) ? ( n22124 ) : ( n48902 ) ;
assign n48904 =  ( n162 ) ? ( n22123 ) : ( n48903 ) ;
assign n48905 =  ( n22106 ) ? ( VREG_5_3 ) : ( n48904 ) ;
assign n48906 =  ( n3051 ) ? ( n48905 ) : ( VREG_5_3 ) ;
assign n48907 =  ( n3040 ) ? ( n48899 ) : ( n48906 ) ;
assign n48908 =  ( n192 ) ? ( VREG_5_3 ) : ( VREG_5_3 ) ;
assign n48909 =  ( n157 ) ? ( n48907 ) : ( n48908 ) ;
assign n48910 =  ( n6 ) ? ( n48894 ) : ( n48909 ) ;
assign n48911 =  ( n769 ) ? ( n48910 ) : ( VREG_5_3 ) ;
assign n48912 =  ( n148 ) ? ( n23184 ) : ( VREG_5_4 ) ;
assign n48913 =  ( n146 ) ? ( n23183 ) : ( n48912 ) ;
assign n48914 =  ( n144 ) ? ( n23182 ) : ( n48913 ) ;
assign n48915 =  ( n142 ) ? ( n23181 ) : ( n48914 ) ;
assign n48916 =  ( n10 ) ? ( n23180 ) : ( n48915 ) ;
assign n48917 =  ( n148 ) ? ( n24218 ) : ( VREG_5_4 ) ;
assign n48918 =  ( n146 ) ? ( n24217 ) : ( n48917 ) ;
assign n48919 =  ( n144 ) ? ( n24216 ) : ( n48918 ) ;
assign n48920 =  ( n142 ) ? ( n24215 ) : ( n48919 ) ;
assign n48921 =  ( n10 ) ? ( n24214 ) : ( n48920 ) ;
assign n48922 =  ( n24225 ) ? ( VREG_5_4 ) : ( n48916 ) ;
assign n48923 =  ( n24225 ) ? ( VREG_5_4 ) : ( n48921 ) ;
assign n48924 =  ( n3034 ) ? ( n48923 ) : ( VREG_5_4 ) ;
assign n48925 =  ( n2965 ) ? ( n48922 ) : ( n48924 ) ;
assign n48926 =  ( n1930 ) ? ( n48921 ) : ( n48925 ) ;
assign n48927 =  ( n879 ) ? ( n48916 ) : ( n48926 ) ;
assign n48928 =  ( n172 ) ? ( n24236 ) : ( VREG_5_4 ) ;
assign n48929 =  ( n170 ) ? ( n24235 ) : ( n48928 ) ;
assign n48930 =  ( n168 ) ? ( n24234 ) : ( n48929 ) ;
assign n48931 =  ( n166 ) ? ( n24233 ) : ( n48930 ) ;
assign n48932 =  ( n162 ) ? ( n24232 ) : ( n48931 ) ;
assign n48933 =  ( n172 ) ? ( n24246 ) : ( VREG_5_4 ) ;
assign n48934 =  ( n170 ) ? ( n24245 ) : ( n48933 ) ;
assign n48935 =  ( n168 ) ? ( n24244 ) : ( n48934 ) ;
assign n48936 =  ( n166 ) ? ( n24243 ) : ( n48935 ) ;
assign n48937 =  ( n162 ) ? ( n24242 ) : ( n48936 ) ;
assign n48938 =  ( n24225 ) ? ( VREG_5_4 ) : ( n48937 ) ;
assign n48939 =  ( n3051 ) ? ( n48938 ) : ( VREG_5_4 ) ;
assign n48940 =  ( n3040 ) ? ( n48932 ) : ( n48939 ) ;
assign n48941 =  ( n192 ) ? ( VREG_5_4 ) : ( VREG_5_4 ) ;
assign n48942 =  ( n157 ) ? ( n48940 ) : ( n48941 ) ;
assign n48943 =  ( n6 ) ? ( n48927 ) : ( n48942 ) ;
assign n48944 =  ( n769 ) ? ( n48943 ) : ( VREG_5_4 ) ;
assign n48945 =  ( n148 ) ? ( n25303 ) : ( VREG_5_5 ) ;
assign n48946 =  ( n146 ) ? ( n25302 ) : ( n48945 ) ;
assign n48947 =  ( n144 ) ? ( n25301 ) : ( n48946 ) ;
assign n48948 =  ( n142 ) ? ( n25300 ) : ( n48947 ) ;
assign n48949 =  ( n10 ) ? ( n25299 ) : ( n48948 ) ;
assign n48950 =  ( n148 ) ? ( n26337 ) : ( VREG_5_5 ) ;
assign n48951 =  ( n146 ) ? ( n26336 ) : ( n48950 ) ;
assign n48952 =  ( n144 ) ? ( n26335 ) : ( n48951 ) ;
assign n48953 =  ( n142 ) ? ( n26334 ) : ( n48952 ) ;
assign n48954 =  ( n10 ) ? ( n26333 ) : ( n48953 ) ;
assign n48955 =  ( n26344 ) ? ( VREG_5_5 ) : ( n48949 ) ;
assign n48956 =  ( n26344 ) ? ( VREG_5_5 ) : ( n48954 ) ;
assign n48957 =  ( n3034 ) ? ( n48956 ) : ( VREG_5_5 ) ;
assign n48958 =  ( n2965 ) ? ( n48955 ) : ( n48957 ) ;
assign n48959 =  ( n1930 ) ? ( n48954 ) : ( n48958 ) ;
assign n48960 =  ( n879 ) ? ( n48949 ) : ( n48959 ) ;
assign n48961 =  ( n172 ) ? ( n26355 ) : ( VREG_5_5 ) ;
assign n48962 =  ( n170 ) ? ( n26354 ) : ( n48961 ) ;
assign n48963 =  ( n168 ) ? ( n26353 ) : ( n48962 ) ;
assign n48964 =  ( n166 ) ? ( n26352 ) : ( n48963 ) ;
assign n48965 =  ( n162 ) ? ( n26351 ) : ( n48964 ) ;
assign n48966 =  ( n172 ) ? ( n26365 ) : ( VREG_5_5 ) ;
assign n48967 =  ( n170 ) ? ( n26364 ) : ( n48966 ) ;
assign n48968 =  ( n168 ) ? ( n26363 ) : ( n48967 ) ;
assign n48969 =  ( n166 ) ? ( n26362 ) : ( n48968 ) ;
assign n48970 =  ( n162 ) ? ( n26361 ) : ( n48969 ) ;
assign n48971 =  ( n26344 ) ? ( VREG_5_5 ) : ( n48970 ) ;
assign n48972 =  ( n3051 ) ? ( n48971 ) : ( VREG_5_5 ) ;
assign n48973 =  ( n3040 ) ? ( n48965 ) : ( n48972 ) ;
assign n48974 =  ( n192 ) ? ( VREG_5_5 ) : ( VREG_5_5 ) ;
assign n48975 =  ( n157 ) ? ( n48973 ) : ( n48974 ) ;
assign n48976 =  ( n6 ) ? ( n48960 ) : ( n48975 ) ;
assign n48977 =  ( n769 ) ? ( n48976 ) : ( VREG_5_5 ) ;
assign n48978 =  ( n148 ) ? ( n27422 ) : ( VREG_5_6 ) ;
assign n48979 =  ( n146 ) ? ( n27421 ) : ( n48978 ) ;
assign n48980 =  ( n144 ) ? ( n27420 ) : ( n48979 ) ;
assign n48981 =  ( n142 ) ? ( n27419 ) : ( n48980 ) ;
assign n48982 =  ( n10 ) ? ( n27418 ) : ( n48981 ) ;
assign n48983 =  ( n148 ) ? ( n28456 ) : ( VREG_5_6 ) ;
assign n48984 =  ( n146 ) ? ( n28455 ) : ( n48983 ) ;
assign n48985 =  ( n144 ) ? ( n28454 ) : ( n48984 ) ;
assign n48986 =  ( n142 ) ? ( n28453 ) : ( n48985 ) ;
assign n48987 =  ( n10 ) ? ( n28452 ) : ( n48986 ) ;
assign n48988 =  ( n28463 ) ? ( VREG_5_6 ) : ( n48982 ) ;
assign n48989 =  ( n28463 ) ? ( VREG_5_6 ) : ( n48987 ) ;
assign n48990 =  ( n3034 ) ? ( n48989 ) : ( VREG_5_6 ) ;
assign n48991 =  ( n2965 ) ? ( n48988 ) : ( n48990 ) ;
assign n48992 =  ( n1930 ) ? ( n48987 ) : ( n48991 ) ;
assign n48993 =  ( n879 ) ? ( n48982 ) : ( n48992 ) ;
assign n48994 =  ( n172 ) ? ( n28474 ) : ( VREG_5_6 ) ;
assign n48995 =  ( n170 ) ? ( n28473 ) : ( n48994 ) ;
assign n48996 =  ( n168 ) ? ( n28472 ) : ( n48995 ) ;
assign n48997 =  ( n166 ) ? ( n28471 ) : ( n48996 ) ;
assign n48998 =  ( n162 ) ? ( n28470 ) : ( n48997 ) ;
assign n48999 =  ( n172 ) ? ( n28484 ) : ( VREG_5_6 ) ;
assign n49000 =  ( n170 ) ? ( n28483 ) : ( n48999 ) ;
assign n49001 =  ( n168 ) ? ( n28482 ) : ( n49000 ) ;
assign n49002 =  ( n166 ) ? ( n28481 ) : ( n49001 ) ;
assign n49003 =  ( n162 ) ? ( n28480 ) : ( n49002 ) ;
assign n49004 =  ( n28463 ) ? ( VREG_5_6 ) : ( n49003 ) ;
assign n49005 =  ( n3051 ) ? ( n49004 ) : ( VREG_5_6 ) ;
assign n49006 =  ( n3040 ) ? ( n48998 ) : ( n49005 ) ;
assign n49007 =  ( n192 ) ? ( VREG_5_6 ) : ( VREG_5_6 ) ;
assign n49008 =  ( n157 ) ? ( n49006 ) : ( n49007 ) ;
assign n49009 =  ( n6 ) ? ( n48993 ) : ( n49008 ) ;
assign n49010 =  ( n769 ) ? ( n49009 ) : ( VREG_5_6 ) ;
assign n49011 =  ( n148 ) ? ( n29541 ) : ( VREG_5_7 ) ;
assign n49012 =  ( n146 ) ? ( n29540 ) : ( n49011 ) ;
assign n49013 =  ( n144 ) ? ( n29539 ) : ( n49012 ) ;
assign n49014 =  ( n142 ) ? ( n29538 ) : ( n49013 ) ;
assign n49015 =  ( n10 ) ? ( n29537 ) : ( n49014 ) ;
assign n49016 =  ( n148 ) ? ( n30575 ) : ( VREG_5_7 ) ;
assign n49017 =  ( n146 ) ? ( n30574 ) : ( n49016 ) ;
assign n49018 =  ( n144 ) ? ( n30573 ) : ( n49017 ) ;
assign n49019 =  ( n142 ) ? ( n30572 ) : ( n49018 ) ;
assign n49020 =  ( n10 ) ? ( n30571 ) : ( n49019 ) ;
assign n49021 =  ( n30582 ) ? ( VREG_5_7 ) : ( n49015 ) ;
assign n49022 =  ( n30582 ) ? ( VREG_5_7 ) : ( n49020 ) ;
assign n49023 =  ( n3034 ) ? ( n49022 ) : ( VREG_5_7 ) ;
assign n49024 =  ( n2965 ) ? ( n49021 ) : ( n49023 ) ;
assign n49025 =  ( n1930 ) ? ( n49020 ) : ( n49024 ) ;
assign n49026 =  ( n879 ) ? ( n49015 ) : ( n49025 ) ;
assign n49027 =  ( n172 ) ? ( n30593 ) : ( VREG_5_7 ) ;
assign n49028 =  ( n170 ) ? ( n30592 ) : ( n49027 ) ;
assign n49029 =  ( n168 ) ? ( n30591 ) : ( n49028 ) ;
assign n49030 =  ( n166 ) ? ( n30590 ) : ( n49029 ) ;
assign n49031 =  ( n162 ) ? ( n30589 ) : ( n49030 ) ;
assign n49032 =  ( n172 ) ? ( n30603 ) : ( VREG_5_7 ) ;
assign n49033 =  ( n170 ) ? ( n30602 ) : ( n49032 ) ;
assign n49034 =  ( n168 ) ? ( n30601 ) : ( n49033 ) ;
assign n49035 =  ( n166 ) ? ( n30600 ) : ( n49034 ) ;
assign n49036 =  ( n162 ) ? ( n30599 ) : ( n49035 ) ;
assign n49037 =  ( n30582 ) ? ( VREG_5_7 ) : ( n49036 ) ;
assign n49038 =  ( n3051 ) ? ( n49037 ) : ( VREG_5_7 ) ;
assign n49039 =  ( n3040 ) ? ( n49031 ) : ( n49038 ) ;
assign n49040 =  ( n192 ) ? ( VREG_5_7 ) : ( VREG_5_7 ) ;
assign n49041 =  ( n157 ) ? ( n49039 ) : ( n49040 ) ;
assign n49042 =  ( n6 ) ? ( n49026 ) : ( n49041 ) ;
assign n49043 =  ( n769 ) ? ( n49042 ) : ( VREG_5_7 ) ;
assign n49044 =  ( n148 ) ? ( n31660 ) : ( VREG_5_8 ) ;
assign n49045 =  ( n146 ) ? ( n31659 ) : ( n49044 ) ;
assign n49046 =  ( n144 ) ? ( n31658 ) : ( n49045 ) ;
assign n49047 =  ( n142 ) ? ( n31657 ) : ( n49046 ) ;
assign n49048 =  ( n10 ) ? ( n31656 ) : ( n49047 ) ;
assign n49049 =  ( n148 ) ? ( n32694 ) : ( VREG_5_8 ) ;
assign n49050 =  ( n146 ) ? ( n32693 ) : ( n49049 ) ;
assign n49051 =  ( n144 ) ? ( n32692 ) : ( n49050 ) ;
assign n49052 =  ( n142 ) ? ( n32691 ) : ( n49051 ) ;
assign n49053 =  ( n10 ) ? ( n32690 ) : ( n49052 ) ;
assign n49054 =  ( n32701 ) ? ( VREG_5_8 ) : ( n49048 ) ;
assign n49055 =  ( n32701 ) ? ( VREG_5_8 ) : ( n49053 ) ;
assign n49056 =  ( n3034 ) ? ( n49055 ) : ( VREG_5_8 ) ;
assign n49057 =  ( n2965 ) ? ( n49054 ) : ( n49056 ) ;
assign n49058 =  ( n1930 ) ? ( n49053 ) : ( n49057 ) ;
assign n49059 =  ( n879 ) ? ( n49048 ) : ( n49058 ) ;
assign n49060 =  ( n172 ) ? ( n32712 ) : ( VREG_5_8 ) ;
assign n49061 =  ( n170 ) ? ( n32711 ) : ( n49060 ) ;
assign n49062 =  ( n168 ) ? ( n32710 ) : ( n49061 ) ;
assign n49063 =  ( n166 ) ? ( n32709 ) : ( n49062 ) ;
assign n49064 =  ( n162 ) ? ( n32708 ) : ( n49063 ) ;
assign n49065 =  ( n172 ) ? ( n32722 ) : ( VREG_5_8 ) ;
assign n49066 =  ( n170 ) ? ( n32721 ) : ( n49065 ) ;
assign n49067 =  ( n168 ) ? ( n32720 ) : ( n49066 ) ;
assign n49068 =  ( n166 ) ? ( n32719 ) : ( n49067 ) ;
assign n49069 =  ( n162 ) ? ( n32718 ) : ( n49068 ) ;
assign n49070 =  ( n32701 ) ? ( VREG_5_8 ) : ( n49069 ) ;
assign n49071 =  ( n3051 ) ? ( n49070 ) : ( VREG_5_8 ) ;
assign n49072 =  ( n3040 ) ? ( n49064 ) : ( n49071 ) ;
assign n49073 =  ( n192 ) ? ( VREG_5_8 ) : ( VREG_5_8 ) ;
assign n49074 =  ( n157 ) ? ( n49072 ) : ( n49073 ) ;
assign n49075 =  ( n6 ) ? ( n49059 ) : ( n49074 ) ;
assign n49076 =  ( n769 ) ? ( n49075 ) : ( VREG_5_8 ) ;
assign n49077 =  ( n148 ) ? ( n33779 ) : ( VREG_5_9 ) ;
assign n49078 =  ( n146 ) ? ( n33778 ) : ( n49077 ) ;
assign n49079 =  ( n144 ) ? ( n33777 ) : ( n49078 ) ;
assign n49080 =  ( n142 ) ? ( n33776 ) : ( n49079 ) ;
assign n49081 =  ( n10 ) ? ( n33775 ) : ( n49080 ) ;
assign n49082 =  ( n148 ) ? ( n34813 ) : ( VREG_5_9 ) ;
assign n49083 =  ( n146 ) ? ( n34812 ) : ( n49082 ) ;
assign n49084 =  ( n144 ) ? ( n34811 ) : ( n49083 ) ;
assign n49085 =  ( n142 ) ? ( n34810 ) : ( n49084 ) ;
assign n49086 =  ( n10 ) ? ( n34809 ) : ( n49085 ) ;
assign n49087 =  ( n34820 ) ? ( VREG_5_9 ) : ( n49081 ) ;
assign n49088 =  ( n34820 ) ? ( VREG_5_9 ) : ( n49086 ) ;
assign n49089 =  ( n3034 ) ? ( n49088 ) : ( VREG_5_9 ) ;
assign n49090 =  ( n2965 ) ? ( n49087 ) : ( n49089 ) ;
assign n49091 =  ( n1930 ) ? ( n49086 ) : ( n49090 ) ;
assign n49092 =  ( n879 ) ? ( n49081 ) : ( n49091 ) ;
assign n49093 =  ( n172 ) ? ( n34831 ) : ( VREG_5_9 ) ;
assign n49094 =  ( n170 ) ? ( n34830 ) : ( n49093 ) ;
assign n49095 =  ( n168 ) ? ( n34829 ) : ( n49094 ) ;
assign n49096 =  ( n166 ) ? ( n34828 ) : ( n49095 ) ;
assign n49097 =  ( n162 ) ? ( n34827 ) : ( n49096 ) ;
assign n49098 =  ( n172 ) ? ( n34841 ) : ( VREG_5_9 ) ;
assign n49099 =  ( n170 ) ? ( n34840 ) : ( n49098 ) ;
assign n49100 =  ( n168 ) ? ( n34839 ) : ( n49099 ) ;
assign n49101 =  ( n166 ) ? ( n34838 ) : ( n49100 ) ;
assign n49102 =  ( n162 ) ? ( n34837 ) : ( n49101 ) ;
assign n49103 =  ( n34820 ) ? ( VREG_5_9 ) : ( n49102 ) ;
assign n49104 =  ( n3051 ) ? ( n49103 ) : ( VREG_5_9 ) ;
assign n49105 =  ( n3040 ) ? ( n49097 ) : ( n49104 ) ;
assign n49106 =  ( n192 ) ? ( VREG_5_9 ) : ( VREG_5_9 ) ;
assign n49107 =  ( n157 ) ? ( n49105 ) : ( n49106 ) ;
assign n49108 =  ( n6 ) ? ( n49092 ) : ( n49107 ) ;
assign n49109 =  ( n769 ) ? ( n49108 ) : ( VREG_5_9 ) ;
assign n49110 =  ( n148 ) ? ( n1924 ) : ( VREG_6_0 ) ;
assign n49111 =  ( n146 ) ? ( n1923 ) : ( n49110 ) ;
assign n49112 =  ( n144 ) ? ( n1922 ) : ( n49111 ) ;
assign n49113 =  ( n142 ) ? ( n1921 ) : ( n49112 ) ;
assign n49114 =  ( n10 ) ? ( n1920 ) : ( n49113 ) ;
assign n49115 =  ( n148 ) ? ( n2959 ) : ( VREG_6_0 ) ;
assign n49116 =  ( n146 ) ? ( n2958 ) : ( n49115 ) ;
assign n49117 =  ( n144 ) ? ( n2957 ) : ( n49116 ) ;
assign n49118 =  ( n142 ) ? ( n2956 ) : ( n49117 ) ;
assign n49119 =  ( n10 ) ? ( n2955 ) : ( n49118 ) ;
assign n49120 =  ( n3032 ) ? ( VREG_6_0 ) : ( n49114 ) ;
assign n49121 =  ( n3032 ) ? ( VREG_6_0 ) : ( n49119 ) ;
assign n49122 =  ( n3034 ) ? ( n49121 ) : ( VREG_6_0 ) ;
assign n49123 =  ( n2965 ) ? ( n49120 ) : ( n49122 ) ;
assign n49124 =  ( n1930 ) ? ( n49119 ) : ( n49123 ) ;
assign n49125 =  ( n879 ) ? ( n49114 ) : ( n49124 ) ;
assign n49126 =  ( n172 ) ? ( n3045 ) : ( VREG_6_0 ) ;
assign n49127 =  ( n170 ) ? ( n3044 ) : ( n49126 ) ;
assign n49128 =  ( n168 ) ? ( n3043 ) : ( n49127 ) ;
assign n49129 =  ( n166 ) ? ( n3042 ) : ( n49128 ) ;
assign n49130 =  ( n162 ) ? ( n3041 ) : ( n49129 ) ;
assign n49131 =  ( n172 ) ? ( n3056 ) : ( VREG_6_0 ) ;
assign n49132 =  ( n170 ) ? ( n3055 ) : ( n49131 ) ;
assign n49133 =  ( n168 ) ? ( n3054 ) : ( n49132 ) ;
assign n49134 =  ( n166 ) ? ( n3053 ) : ( n49133 ) ;
assign n49135 =  ( n162 ) ? ( n3052 ) : ( n49134 ) ;
assign n49136 =  ( n3032 ) ? ( VREG_6_0 ) : ( n49135 ) ;
assign n49137 =  ( n3051 ) ? ( n49136 ) : ( VREG_6_0 ) ;
assign n49138 =  ( n3040 ) ? ( n49130 ) : ( n49137 ) ;
assign n49139 =  ( n192 ) ? ( VREG_6_0 ) : ( VREG_6_0 ) ;
assign n49140 =  ( n157 ) ? ( n49138 ) : ( n49139 ) ;
assign n49141 =  ( n6 ) ? ( n49125 ) : ( n49140 ) ;
assign n49142 =  ( n791 ) ? ( n49141 ) : ( VREG_6_0 ) ;
assign n49143 =  ( n148 ) ? ( n4113 ) : ( VREG_6_1 ) ;
assign n49144 =  ( n146 ) ? ( n4112 ) : ( n49143 ) ;
assign n49145 =  ( n144 ) ? ( n4111 ) : ( n49144 ) ;
assign n49146 =  ( n142 ) ? ( n4110 ) : ( n49145 ) ;
assign n49147 =  ( n10 ) ? ( n4109 ) : ( n49146 ) ;
assign n49148 =  ( n148 ) ? ( n5147 ) : ( VREG_6_1 ) ;
assign n49149 =  ( n146 ) ? ( n5146 ) : ( n49148 ) ;
assign n49150 =  ( n144 ) ? ( n5145 ) : ( n49149 ) ;
assign n49151 =  ( n142 ) ? ( n5144 ) : ( n49150 ) ;
assign n49152 =  ( n10 ) ? ( n5143 ) : ( n49151 ) ;
assign n49153 =  ( n5154 ) ? ( VREG_6_1 ) : ( n49147 ) ;
assign n49154 =  ( n5154 ) ? ( VREG_6_1 ) : ( n49152 ) ;
assign n49155 =  ( n3034 ) ? ( n49154 ) : ( VREG_6_1 ) ;
assign n49156 =  ( n2965 ) ? ( n49153 ) : ( n49155 ) ;
assign n49157 =  ( n1930 ) ? ( n49152 ) : ( n49156 ) ;
assign n49158 =  ( n879 ) ? ( n49147 ) : ( n49157 ) ;
assign n49159 =  ( n172 ) ? ( n5165 ) : ( VREG_6_1 ) ;
assign n49160 =  ( n170 ) ? ( n5164 ) : ( n49159 ) ;
assign n49161 =  ( n168 ) ? ( n5163 ) : ( n49160 ) ;
assign n49162 =  ( n166 ) ? ( n5162 ) : ( n49161 ) ;
assign n49163 =  ( n162 ) ? ( n5161 ) : ( n49162 ) ;
assign n49164 =  ( n172 ) ? ( n5175 ) : ( VREG_6_1 ) ;
assign n49165 =  ( n170 ) ? ( n5174 ) : ( n49164 ) ;
assign n49166 =  ( n168 ) ? ( n5173 ) : ( n49165 ) ;
assign n49167 =  ( n166 ) ? ( n5172 ) : ( n49166 ) ;
assign n49168 =  ( n162 ) ? ( n5171 ) : ( n49167 ) ;
assign n49169 =  ( n5154 ) ? ( VREG_6_1 ) : ( n49168 ) ;
assign n49170 =  ( n3051 ) ? ( n49169 ) : ( VREG_6_1 ) ;
assign n49171 =  ( n3040 ) ? ( n49163 ) : ( n49170 ) ;
assign n49172 =  ( n192 ) ? ( VREG_6_1 ) : ( VREG_6_1 ) ;
assign n49173 =  ( n157 ) ? ( n49171 ) : ( n49172 ) ;
assign n49174 =  ( n6 ) ? ( n49158 ) : ( n49173 ) ;
assign n49175 =  ( n791 ) ? ( n49174 ) : ( VREG_6_1 ) ;
assign n49176 =  ( n148 ) ? ( n6232 ) : ( VREG_6_10 ) ;
assign n49177 =  ( n146 ) ? ( n6231 ) : ( n49176 ) ;
assign n49178 =  ( n144 ) ? ( n6230 ) : ( n49177 ) ;
assign n49179 =  ( n142 ) ? ( n6229 ) : ( n49178 ) ;
assign n49180 =  ( n10 ) ? ( n6228 ) : ( n49179 ) ;
assign n49181 =  ( n148 ) ? ( n7266 ) : ( VREG_6_10 ) ;
assign n49182 =  ( n146 ) ? ( n7265 ) : ( n49181 ) ;
assign n49183 =  ( n144 ) ? ( n7264 ) : ( n49182 ) ;
assign n49184 =  ( n142 ) ? ( n7263 ) : ( n49183 ) ;
assign n49185 =  ( n10 ) ? ( n7262 ) : ( n49184 ) ;
assign n49186 =  ( n7273 ) ? ( VREG_6_10 ) : ( n49180 ) ;
assign n49187 =  ( n7273 ) ? ( VREG_6_10 ) : ( n49185 ) ;
assign n49188 =  ( n3034 ) ? ( n49187 ) : ( VREG_6_10 ) ;
assign n49189 =  ( n2965 ) ? ( n49186 ) : ( n49188 ) ;
assign n49190 =  ( n1930 ) ? ( n49185 ) : ( n49189 ) ;
assign n49191 =  ( n879 ) ? ( n49180 ) : ( n49190 ) ;
assign n49192 =  ( n172 ) ? ( n7284 ) : ( VREG_6_10 ) ;
assign n49193 =  ( n170 ) ? ( n7283 ) : ( n49192 ) ;
assign n49194 =  ( n168 ) ? ( n7282 ) : ( n49193 ) ;
assign n49195 =  ( n166 ) ? ( n7281 ) : ( n49194 ) ;
assign n49196 =  ( n162 ) ? ( n7280 ) : ( n49195 ) ;
assign n49197 =  ( n172 ) ? ( n7294 ) : ( VREG_6_10 ) ;
assign n49198 =  ( n170 ) ? ( n7293 ) : ( n49197 ) ;
assign n49199 =  ( n168 ) ? ( n7292 ) : ( n49198 ) ;
assign n49200 =  ( n166 ) ? ( n7291 ) : ( n49199 ) ;
assign n49201 =  ( n162 ) ? ( n7290 ) : ( n49200 ) ;
assign n49202 =  ( n7273 ) ? ( VREG_6_10 ) : ( n49201 ) ;
assign n49203 =  ( n3051 ) ? ( n49202 ) : ( VREG_6_10 ) ;
assign n49204 =  ( n3040 ) ? ( n49196 ) : ( n49203 ) ;
assign n49205 =  ( n192 ) ? ( VREG_6_10 ) : ( VREG_6_10 ) ;
assign n49206 =  ( n157 ) ? ( n49204 ) : ( n49205 ) ;
assign n49207 =  ( n6 ) ? ( n49191 ) : ( n49206 ) ;
assign n49208 =  ( n791 ) ? ( n49207 ) : ( VREG_6_10 ) ;
assign n49209 =  ( n148 ) ? ( n8351 ) : ( VREG_6_11 ) ;
assign n49210 =  ( n146 ) ? ( n8350 ) : ( n49209 ) ;
assign n49211 =  ( n144 ) ? ( n8349 ) : ( n49210 ) ;
assign n49212 =  ( n142 ) ? ( n8348 ) : ( n49211 ) ;
assign n49213 =  ( n10 ) ? ( n8347 ) : ( n49212 ) ;
assign n49214 =  ( n148 ) ? ( n9385 ) : ( VREG_6_11 ) ;
assign n49215 =  ( n146 ) ? ( n9384 ) : ( n49214 ) ;
assign n49216 =  ( n144 ) ? ( n9383 ) : ( n49215 ) ;
assign n49217 =  ( n142 ) ? ( n9382 ) : ( n49216 ) ;
assign n49218 =  ( n10 ) ? ( n9381 ) : ( n49217 ) ;
assign n49219 =  ( n9392 ) ? ( VREG_6_11 ) : ( n49213 ) ;
assign n49220 =  ( n9392 ) ? ( VREG_6_11 ) : ( n49218 ) ;
assign n49221 =  ( n3034 ) ? ( n49220 ) : ( VREG_6_11 ) ;
assign n49222 =  ( n2965 ) ? ( n49219 ) : ( n49221 ) ;
assign n49223 =  ( n1930 ) ? ( n49218 ) : ( n49222 ) ;
assign n49224 =  ( n879 ) ? ( n49213 ) : ( n49223 ) ;
assign n49225 =  ( n172 ) ? ( n9403 ) : ( VREG_6_11 ) ;
assign n49226 =  ( n170 ) ? ( n9402 ) : ( n49225 ) ;
assign n49227 =  ( n168 ) ? ( n9401 ) : ( n49226 ) ;
assign n49228 =  ( n166 ) ? ( n9400 ) : ( n49227 ) ;
assign n49229 =  ( n162 ) ? ( n9399 ) : ( n49228 ) ;
assign n49230 =  ( n172 ) ? ( n9413 ) : ( VREG_6_11 ) ;
assign n49231 =  ( n170 ) ? ( n9412 ) : ( n49230 ) ;
assign n49232 =  ( n168 ) ? ( n9411 ) : ( n49231 ) ;
assign n49233 =  ( n166 ) ? ( n9410 ) : ( n49232 ) ;
assign n49234 =  ( n162 ) ? ( n9409 ) : ( n49233 ) ;
assign n49235 =  ( n9392 ) ? ( VREG_6_11 ) : ( n49234 ) ;
assign n49236 =  ( n3051 ) ? ( n49235 ) : ( VREG_6_11 ) ;
assign n49237 =  ( n3040 ) ? ( n49229 ) : ( n49236 ) ;
assign n49238 =  ( n192 ) ? ( VREG_6_11 ) : ( VREG_6_11 ) ;
assign n49239 =  ( n157 ) ? ( n49237 ) : ( n49238 ) ;
assign n49240 =  ( n6 ) ? ( n49224 ) : ( n49239 ) ;
assign n49241 =  ( n791 ) ? ( n49240 ) : ( VREG_6_11 ) ;
assign n49242 =  ( n148 ) ? ( n10470 ) : ( VREG_6_12 ) ;
assign n49243 =  ( n146 ) ? ( n10469 ) : ( n49242 ) ;
assign n49244 =  ( n144 ) ? ( n10468 ) : ( n49243 ) ;
assign n49245 =  ( n142 ) ? ( n10467 ) : ( n49244 ) ;
assign n49246 =  ( n10 ) ? ( n10466 ) : ( n49245 ) ;
assign n49247 =  ( n148 ) ? ( n11504 ) : ( VREG_6_12 ) ;
assign n49248 =  ( n146 ) ? ( n11503 ) : ( n49247 ) ;
assign n49249 =  ( n144 ) ? ( n11502 ) : ( n49248 ) ;
assign n49250 =  ( n142 ) ? ( n11501 ) : ( n49249 ) ;
assign n49251 =  ( n10 ) ? ( n11500 ) : ( n49250 ) ;
assign n49252 =  ( n11511 ) ? ( VREG_6_12 ) : ( n49246 ) ;
assign n49253 =  ( n11511 ) ? ( VREG_6_12 ) : ( n49251 ) ;
assign n49254 =  ( n3034 ) ? ( n49253 ) : ( VREG_6_12 ) ;
assign n49255 =  ( n2965 ) ? ( n49252 ) : ( n49254 ) ;
assign n49256 =  ( n1930 ) ? ( n49251 ) : ( n49255 ) ;
assign n49257 =  ( n879 ) ? ( n49246 ) : ( n49256 ) ;
assign n49258 =  ( n172 ) ? ( n11522 ) : ( VREG_6_12 ) ;
assign n49259 =  ( n170 ) ? ( n11521 ) : ( n49258 ) ;
assign n49260 =  ( n168 ) ? ( n11520 ) : ( n49259 ) ;
assign n49261 =  ( n166 ) ? ( n11519 ) : ( n49260 ) ;
assign n49262 =  ( n162 ) ? ( n11518 ) : ( n49261 ) ;
assign n49263 =  ( n172 ) ? ( n11532 ) : ( VREG_6_12 ) ;
assign n49264 =  ( n170 ) ? ( n11531 ) : ( n49263 ) ;
assign n49265 =  ( n168 ) ? ( n11530 ) : ( n49264 ) ;
assign n49266 =  ( n166 ) ? ( n11529 ) : ( n49265 ) ;
assign n49267 =  ( n162 ) ? ( n11528 ) : ( n49266 ) ;
assign n49268 =  ( n11511 ) ? ( VREG_6_12 ) : ( n49267 ) ;
assign n49269 =  ( n3051 ) ? ( n49268 ) : ( VREG_6_12 ) ;
assign n49270 =  ( n3040 ) ? ( n49262 ) : ( n49269 ) ;
assign n49271 =  ( n192 ) ? ( VREG_6_12 ) : ( VREG_6_12 ) ;
assign n49272 =  ( n157 ) ? ( n49270 ) : ( n49271 ) ;
assign n49273 =  ( n6 ) ? ( n49257 ) : ( n49272 ) ;
assign n49274 =  ( n791 ) ? ( n49273 ) : ( VREG_6_12 ) ;
assign n49275 =  ( n148 ) ? ( n12589 ) : ( VREG_6_13 ) ;
assign n49276 =  ( n146 ) ? ( n12588 ) : ( n49275 ) ;
assign n49277 =  ( n144 ) ? ( n12587 ) : ( n49276 ) ;
assign n49278 =  ( n142 ) ? ( n12586 ) : ( n49277 ) ;
assign n49279 =  ( n10 ) ? ( n12585 ) : ( n49278 ) ;
assign n49280 =  ( n148 ) ? ( n13623 ) : ( VREG_6_13 ) ;
assign n49281 =  ( n146 ) ? ( n13622 ) : ( n49280 ) ;
assign n49282 =  ( n144 ) ? ( n13621 ) : ( n49281 ) ;
assign n49283 =  ( n142 ) ? ( n13620 ) : ( n49282 ) ;
assign n49284 =  ( n10 ) ? ( n13619 ) : ( n49283 ) ;
assign n49285 =  ( n13630 ) ? ( VREG_6_13 ) : ( n49279 ) ;
assign n49286 =  ( n13630 ) ? ( VREG_6_13 ) : ( n49284 ) ;
assign n49287 =  ( n3034 ) ? ( n49286 ) : ( VREG_6_13 ) ;
assign n49288 =  ( n2965 ) ? ( n49285 ) : ( n49287 ) ;
assign n49289 =  ( n1930 ) ? ( n49284 ) : ( n49288 ) ;
assign n49290 =  ( n879 ) ? ( n49279 ) : ( n49289 ) ;
assign n49291 =  ( n172 ) ? ( n13641 ) : ( VREG_6_13 ) ;
assign n49292 =  ( n170 ) ? ( n13640 ) : ( n49291 ) ;
assign n49293 =  ( n168 ) ? ( n13639 ) : ( n49292 ) ;
assign n49294 =  ( n166 ) ? ( n13638 ) : ( n49293 ) ;
assign n49295 =  ( n162 ) ? ( n13637 ) : ( n49294 ) ;
assign n49296 =  ( n172 ) ? ( n13651 ) : ( VREG_6_13 ) ;
assign n49297 =  ( n170 ) ? ( n13650 ) : ( n49296 ) ;
assign n49298 =  ( n168 ) ? ( n13649 ) : ( n49297 ) ;
assign n49299 =  ( n166 ) ? ( n13648 ) : ( n49298 ) ;
assign n49300 =  ( n162 ) ? ( n13647 ) : ( n49299 ) ;
assign n49301 =  ( n13630 ) ? ( VREG_6_13 ) : ( n49300 ) ;
assign n49302 =  ( n3051 ) ? ( n49301 ) : ( VREG_6_13 ) ;
assign n49303 =  ( n3040 ) ? ( n49295 ) : ( n49302 ) ;
assign n49304 =  ( n192 ) ? ( VREG_6_13 ) : ( VREG_6_13 ) ;
assign n49305 =  ( n157 ) ? ( n49303 ) : ( n49304 ) ;
assign n49306 =  ( n6 ) ? ( n49290 ) : ( n49305 ) ;
assign n49307 =  ( n791 ) ? ( n49306 ) : ( VREG_6_13 ) ;
assign n49308 =  ( n148 ) ? ( n14708 ) : ( VREG_6_14 ) ;
assign n49309 =  ( n146 ) ? ( n14707 ) : ( n49308 ) ;
assign n49310 =  ( n144 ) ? ( n14706 ) : ( n49309 ) ;
assign n49311 =  ( n142 ) ? ( n14705 ) : ( n49310 ) ;
assign n49312 =  ( n10 ) ? ( n14704 ) : ( n49311 ) ;
assign n49313 =  ( n148 ) ? ( n15742 ) : ( VREG_6_14 ) ;
assign n49314 =  ( n146 ) ? ( n15741 ) : ( n49313 ) ;
assign n49315 =  ( n144 ) ? ( n15740 ) : ( n49314 ) ;
assign n49316 =  ( n142 ) ? ( n15739 ) : ( n49315 ) ;
assign n49317 =  ( n10 ) ? ( n15738 ) : ( n49316 ) ;
assign n49318 =  ( n15749 ) ? ( VREG_6_14 ) : ( n49312 ) ;
assign n49319 =  ( n15749 ) ? ( VREG_6_14 ) : ( n49317 ) ;
assign n49320 =  ( n3034 ) ? ( n49319 ) : ( VREG_6_14 ) ;
assign n49321 =  ( n2965 ) ? ( n49318 ) : ( n49320 ) ;
assign n49322 =  ( n1930 ) ? ( n49317 ) : ( n49321 ) ;
assign n49323 =  ( n879 ) ? ( n49312 ) : ( n49322 ) ;
assign n49324 =  ( n172 ) ? ( n15760 ) : ( VREG_6_14 ) ;
assign n49325 =  ( n170 ) ? ( n15759 ) : ( n49324 ) ;
assign n49326 =  ( n168 ) ? ( n15758 ) : ( n49325 ) ;
assign n49327 =  ( n166 ) ? ( n15757 ) : ( n49326 ) ;
assign n49328 =  ( n162 ) ? ( n15756 ) : ( n49327 ) ;
assign n49329 =  ( n172 ) ? ( n15770 ) : ( VREG_6_14 ) ;
assign n49330 =  ( n170 ) ? ( n15769 ) : ( n49329 ) ;
assign n49331 =  ( n168 ) ? ( n15768 ) : ( n49330 ) ;
assign n49332 =  ( n166 ) ? ( n15767 ) : ( n49331 ) ;
assign n49333 =  ( n162 ) ? ( n15766 ) : ( n49332 ) ;
assign n49334 =  ( n15749 ) ? ( VREG_6_14 ) : ( n49333 ) ;
assign n49335 =  ( n3051 ) ? ( n49334 ) : ( VREG_6_14 ) ;
assign n49336 =  ( n3040 ) ? ( n49328 ) : ( n49335 ) ;
assign n49337 =  ( n192 ) ? ( VREG_6_14 ) : ( VREG_6_14 ) ;
assign n49338 =  ( n157 ) ? ( n49336 ) : ( n49337 ) ;
assign n49339 =  ( n6 ) ? ( n49323 ) : ( n49338 ) ;
assign n49340 =  ( n791 ) ? ( n49339 ) : ( VREG_6_14 ) ;
assign n49341 =  ( n148 ) ? ( n16827 ) : ( VREG_6_15 ) ;
assign n49342 =  ( n146 ) ? ( n16826 ) : ( n49341 ) ;
assign n49343 =  ( n144 ) ? ( n16825 ) : ( n49342 ) ;
assign n49344 =  ( n142 ) ? ( n16824 ) : ( n49343 ) ;
assign n49345 =  ( n10 ) ? ( n16823 ) : ( n49344 ) ;
assign n49346 =  ( n148 ) ? ( n17861 ) : ( VREG_6_15 ) ;
assign n49347 =  ( n146 ) ? ( n17860 ) : ( n49346 ) ;
assign n49348 =  ( n144 ) ? ( n17859 ) : ( n49347 ) ;
assign n49349 =  ( n142 ) ? ( n17858 ) : ( n49348 ) ;
assign n49350 =  ( n10 ) ? ( n17857 ) : ( n49349 ) ;
assign n49351 =  ( n17868 ) ? ( VREG_6_15 ) : ( n49345 ) ;
assign n49352 =  ( n17868 ) ? ( VREG_6_15 ) : ( n49350 ) ;
assign n49353 =  ( n3034 ) ? ( n49352 ) : ( VREG_6_15 ) ;
assign n49354 =  ( n2965 ) ? ( n49351 ) : ( n49353 ) ;
assign n49355 =  ( n1930 ) ? ( n49350 ) : ( n49354 ) ;
assign n49356 =  ( n879 ) ? ( n49345 ) : ( n49355 ) ;
assign n49357 =  ( n172 ) ? ( n17879 ) : ( VREG_6_15 ) ;
assign n49358 =  ( n170 ) ? ( n17878 ) : ( n49357 ) ;
assign n49359 =  ( n168 ) ? ( n17877 ) : ( n49358 ) ;
assign n49360 =  ( n166 ) ? ( n17876 ) : ( n49359 ) ;
assign n49361 =  ( n162 ) ? ( n17875 ) : ( n49360 ) ;
assign n49362 =  ( n172 ) ? ( n17889 ) : ( VREG_6_15 ) ;
assign n49363 =  ( n170 ) ? ( n17888 ) : ( n49362 ) ;
assign n49364 =  ( n168 ) ? ( n17887 ) : ( n49363 ) ;
assign n49365 =  ( n166 ) ? ( n17886 ) : ( n49364 ) ;
assign n49366 =  ( n162 ) ? ( n17885 ) : ( n49365 ) ;
assign n49367 =  ( n17868 ) ? ( VREG_6_15 ) : ( n49366 ) ;
assign n49368 =  ( n3051 ) ? ( n49367 ) : ( VREG_6_15 ) ;
assign n49369 =  ( n3040 ) ? ( n49361 ) : ( n49368 ) ;
assign n49370 =  ( n192 ) ? ( VREG_6_15 ) : ( VREG_6_15 ) ;
assign n49371 =  ( n157 ) ? ( n49369 ) : ( n49370 ) ;
assign n49372 =  ( n6 ) ? ( n49356 ) : ( n49371 ) ;
assign n49373 =  ( n791 ) ? ( n49372 ) : ( VREG_6_15 ) ;
assign n49374 =  ( n148 ) ? ( n18946 ) : ( VREG_6_2 ) ;
assign n49375 =  ( n146 ) ? ( n18945 ) : ( n49374 ) ;
assign n49376 =  ( n144 ) ? ( n18944 ) : ( n49375 ) ;
assign n49377 =  ( n142 ) ? ( n18943 ) : ( n49376 ) ;
assign n49378 =  ( n10 ) ? ( n18942 ) : ( n49377 ) ;
assign n49379 =  ( n148 ) ? ( n19980 ) : ( VREG_6_2 ) ;
assign n49380 =  ( n146 ) ? ( n19979 ) : ( n49379 ) ;
assign n49381 =  ( n144 ) ? ( n19978 ) : ( n49380 ) ;
assign n49382 =  ( n142 ) ? ( n19977 ) : ( n49381 ) ;
assign n49383 =  ( n10 ) ? ( n19976 ) : ( n49382 ) ;
assign n49384 =  ( n19987 ) ? ( VREG_6_2 ) : ( n49378 ) ;
assign n49385 =  ( n19987 ) ? ( VREG_6_2 ) : ( n49383 ) ;
assign n49386 =  ( n3034 ) ? ( n49385 ) : ( VREG_6_2 ) ;
assign n49387 =  ( n2965 ) ? ( n49384 ) : ( n49386 ) ;
assign n49388 =  ( n1930 ) ? ( n49383 ) : ( n49387 ) ;
assign n49389 =  ( n879 ) ? ( n49378 ) : ( n49388 ) ;
assign n49390 =  ( n172 ) ? ( n19998 ) : ( VREG_6_2 ) ;
assign n49391 =  ( n170 ) ? ( n19997 ) : ( n49390 ) ;
assign n49392 =  ( n168 ) ? ( n19996 ) : ( n49391 ) ;
assign n49393 =  ( n166 ) ? ( n19995 ) : ( n49392 ) ;
assign n49394 =  ( n162 ) ? ( n19994 ) : ( n49393 ) ;
assign n49395 =  ( n172 ) ? ( n20008 ) : ( VREG_6_2 ) ;
assign n49396 =  ( n170 ) ? ( n20007 ) : ( n49395 ) ;
assign n49397 =  ( n168 ) ? ( n20006 ) : ( n49396 ) ;
assign n49398 =  ( n166 ) ? ( n20005 ) : ( n49397 ) ;
assign n49399 =  ( n162 ) ? ( n20004 ) : ( n49398 ) ;
assign n49400 =  ( n19987 ) ? ( VREG_6_2 ) : ( n49399 ) ;
assign n49401 =  ( n3051 ) ? ( n49400 ) : ( VREG_6_2 ) ;
assign n49402 =  ( n3040 ) ? ( n49394 ) : ( n49401 ) ;
assign n49403 =  ( n192 ) ? ( VREG_6_2 ) : ( VREG_6_2 ) ;
assign n49404 =  ( n157 ) ? ( n49402 ) : ( n49403 ) ;
assign n49405 =  ( n6 ) ? ( n49389 ) : ( n49404 ) ;
assign n49406 =  ( n791 ) ? ( n49405 ) : ( VREG_6_2 ) ;
assign n49407 =  ( n148 ) ? ( n21065 ) : ( VREG_6_3 ) ;
assign n49408 =  ( n146 ) ? ( n21064 ) : ( n49407 ) ;
assign n49409 =  ( n144 ) ? ( n21063 ) : ( n49408 ) ;
assign n49410 =  ( n142 ) ? ( n21062 ) : ( n49409 ) ;
assign n49411 =  ( n10 ) ? ( n21061 ) : ( n49410 ) ;
assign n49412 =  ( n148 ) ? ( n22099 ) : ( VREG_6_3 ) ;
assign n49413 =  ( n146 ) ? ( n22098 ) : ( n49412 ) ;
assign n49414 =  ( n144 ) ? ( n22097 ) : ( n49413 ) ;
assign n49415 =  ( n142 ) ? ( n22096 ) : ( n49414 ) ;
assign n49416 =  ( n10 ) ? ( n22095 ) : ( n49415 ) ;
assign n49417 =  ( n22106 ) ? ( VREG_6_3 ) : ( n49411 ) ;
assign n49418 =  ( n22106 ) ? ( VREG_6_3 ) : ( n49416 ) ;
assign n49419 =  ( n3034 ) ? ( n49418 ) : ( VREG_6_3 ) ;
assign n49420 =  ( n2965 ) ? ( n49417 ) : ( n49419 ) ;
assign n49421 =  ( n1930 ) ? ( n49416 ) : ( n49420 ) ;
assign n49422 =  ( n879 ) ? ( n49411 ) : ( n49421 ) ;
assign n49423 =  ( n172 ) ? ( n22117 ) : ( VREG_6_3 ) ;
assign n49424 =  ( n170 ) ? ( n22116 ) : ( n49423 ) ;
assign n49425 =  ( n168 ) ? ( n22115 ) : ( n49424 ) ;
assign n49426 =  ( n166 ) ? ( n22114 ) : ( n49425 ) ;
assign n49427 =  ( n162 ) ? ( n22113 ) : ( n49426 ) ;
assign n49428 =  ( n172 ) ? ( n22127 ) : ( VREG_6_3 ) ;
assign n49429 =  ( n170 ) ? ( n22126 ) : ( n49428 ) ;
assign n49430 =  ( n168 ) ? ( n22125 ) : ( n49429 ) ;
assign n49431 =  ( n166 ) ? ( n22124 ) : ( n49430 ) ;
assign n49432 =  ( n162 ) ? ( n22123 ) : ( n49431 ) ;
assign n49433 =  ( n22106 ) ? ( VREG_6_3 ) : ( n49432 ) ;
assign n49434 =  ( n3051 ) ? ( n49433 ) : ( VREG_6_3 ) ;
assign n49435 =  ( n3040 ) ? ( n49427 ) : ( n49434 ) ;
assign n49436 =  ( n192 ) ? ( VREG_6_3 ) : ( VREG_6_3 ) ;
assign n49437 =  ( n157 ) ? ( n49435 ) : ( n49436 ) ;
assign n49438 =  ( n6 ) ? ( n49422 ) : ( n49437 ) ;
assign n49439 =  ( n791 ) ? ( n49438 ) : ( VREG_6_3 ) ;
assign n49440 =  ( n148 ) ? ( n23184 ) : ( VREG_6_4 ) ;
assign n49441 =  ( n146 ) ? ( n23183 ) : ( n49440 ) ;
assign n49442 =  ( n144 ) ? ( n23182 ) : ( n49441 ) ;
assign n49443 =  ( n142 ) ? ( n23181 ) : ( n49442 ) ;
assign n49444 =  ( n10 ) ? ( n23180 ) : ( n49443 ) ;
assign n49445 =  ( n148 ) ? ( n24218 ) : ( VREG_6_4 ) ;
assign n49446 =  ( n146 ) ? ( n24217 ) : ( n49445 ) ;
assign n49447 =  ( n144 ) ? ( n24216 ) : ( n49446 ) ;
assign n49448 =  ( n142 ) ? ( n24215 ) : ( n49447 ) ;
assign n49449 =  ( n10 ) ? ( n24214 ) : ( n49448 ) ;
assign n49450 =  ( n24225 ) ? ( VREG_6_4 ) : ( n49444 ) ;
assign n49451 =  ( n24225 ) ? ( VREG_6_4 ) : ( n49449 ) ;
assign n49452 =  ( n3034 ) ? ( n49451 ) : ( VREG_6_4 ) ;
assign n49453 =  ( n2965 ) ? ( n49450 ) : ( n49452 ) ;
assign n49454 =  ( n1930 ) ? ( n49449 ) : ( n49453 ) ;
assign n49455 =  ( n879 ) ? ( n49444 ) : ( n49454 ) ;
assign n49456 =  ( n172 ) ? ( n24236 ) : ( VREG_6_4 ) ;
assign n49457 =  ( n170 ) ? ( n24235 ) : ( n49456 ) ;
assign n49458 =  ( n168 ) ? ( n24234 ) : ( n49457 ) ;
assign n49459 =  ( n166 ) ? ( n24233 ) : ( n49458 ) ;
assign n49460 =  ( n162 ) ? ( n24232 ) : ( n49459 ) ;
assign n49461 =  ( n172 ) ? ( n24246 ) : ( VREG_6_4 ) ;
assign n49462 =  ( n170 ) ? ( n24245 ) : ( n49461 ) ;
assign n49463 =  ( n168 ) ? ( n24244 ) : ( n49462 ) ;
assign n49464 =  ( n166 ) ? ( n24243 ) : ( n49463 ) ;
assign n49465 =  ( n162 ) ? ( n24242 ) : ( n49464 ) ;
assign n49466 =  ( n24225 ) ? ( VREG_6_4 ) : ( n49465 ) ;
assign n49467 =  ( n3051 ) ? ( n49466 ) : ( VREG_6_4 ) ;
assign n49468 =  ( n3040 ) ? ( n49460 ) : ( n49467 ) ;
assign n49469 =  ( n192 ) ? ( VREG_6_4 ) : ( VREG_6_4 ) ;
assign n49470 =  ( n157 ) ? ( n49468 ) : ( n49469 ) ;
assign n49471 =  ( n6 ) ? ( n49455 ) : ( n49470 ) ;
assign n49472 =  ( n791 ) ? ( n49471 ) : ( VREG_6_4 ) ;
assign n49473 =  ( n148 ) ? ( n25303 ) : ( VREG_6_5 ) ;
assign n49474 =  ( n146 ) ? ( n25302 ) : ( n49473 ) ;
assign n49475 =  ( n144 ) ? ( n25301 ) : ( n49474 ) ;
assign n49476 =  ( n142 ) ? ( n25300 ) : ( n49475 ) ;
assign n49477 =  ( n10 ) ? ( n25299 ) : ( n49476 ) ;
assign n49478 =  ( n148 ) ? ( n26337 ) : ( VREG_6_5 ) ;
assign n49479 =  ( n146 ) ? ( n26336 ) : ( n49478 ) ;
assign n49480 =  ( n144 ) ? ( n26335 ) : ( n49479 ) ;
assign n49481 =  ( n142 ) ? ( n26334 ) : ( n49480 ) ;
assign n49482 =  ( n10 ) ? ( n26333 ) : ( n49481 ) ;
assign n49483 =  ( n26344 ) ? ( VREG_6_5 ) : ( n49477 ) ;
assign n49484 =  ( n26344 ) ? ( VREG_6_5 ) : ( n49482 ) ;
assign n49485 =  ( n3034 ) ? ( n49484 ) : ( VREG_6_5 ) ;
assign n49486 =  ( n2965 ) ? ( n49483 ) : ( n49485 ) ;
assign n49487 =  ( n1930 ) ? ( n49482 ) : ( n49486 ) ;
assign n49488 =  ( n879 ) ? ( n49477 ) : ( n49487 ) ;
assign n49489 =  ( n172 ) ? ( n26355 ) : ( VREG_6_5 ) ;
assign n49490 =  ( n170 ) ? ( n26354 ) : ( n49489 ) ;
assign n49491 =  ( n168 ) ? ( n26353 ) : ( n49490 ) ;
assign n49492 =  ( n166 ) ? ( n26352 ) : ( n49491 ) ;
assign n49493 =  ( n162 ) ? ( n26351 ) : ( n49492 ) ;
assign n49494 =  ( n172 ) ? ( n26365 ) : ( VREG_6_5 ) ;
assign n49495 =  ( n170 ) ? ( n26364 ) : ( n49494 ) ;
assign n49496 =  ( n168 ) ? ( n26363 ) : ( n49495 ) ;
assign n49497 =  ( n166 ) ? ( n26362 ) : ( n49496 ) ;
assign n49498 =  ( n162 ) ? ( n26361 ) : ( n49497 ) ;
assign n49499 =  ( n26344 ) ? ( VREG_6_5 ) : ( n49498 ) ;
assign n49500 =  ( n3051 ) ? ( n49499 ) : ( VREG_6_5 ) ;
assign n49501 =  ( n3040 ) ? ( n49493 ) : ( n49500 ) ;
assign n49502 =  ( n192 ) ? ( VREG_6_5 ) : ( VREG_6_5 ) ;
assign n49503 =  ( n157 ) ? ( n49501 ) : ( n49502 ) ;
assign n49504 =  ( n6 ) ? ( n49488 ) : ( n49503 ) ;
assign n49505 =  ( n791 ) ? ( n49504 ) : ( VREG_6_5 ) ;
assign n49506 =  ( n148 ) ? ( n27422 ) : ( VREG_6_6 ) ;
assign n49507 =  ( n146 ) ? ( n27421 ) : ( n49506 ) ;
assign n49508 =  ( n144 ) ? ( n27420 ) : ( n49507 ) ;
assign n49509 =  ( n142 ) ? ( n27419 ) : ( n49508 ) ;
assign n49510 =  ( n10 ) ? ( n27418 ) : ( n49509 ) ;
assign n49511 =  ( n148 ) ? ( n28456 ) : ( VREG_6_6 ) ;
assign n49512 =  ( n146 ) ? ( n28455 ) : ( n49511 ) ;
assign n49513 =  ( n144 ) ? ( n28454 ) : ( n49512 ) ;
assign n49514 =  ( n142 ) ? ( n28453 ) : ( n49513 ) ;
assign n49515 =  ( n10 ) ? ( n28452 ) : ( n49514 ) ;
assign n49516 =  ( n28463 ) ? ( VREG_6_6 ) : ( n49510 ) ;
assign n49517 =  ( n28463 ) ? ( VREG_6_6 ) : ( n49515 ) ;
assign n49518 =  ( n3034 ) ? ( n49517 ) : ( VREG_6_6 ) ;
assign n49519 =  ( n2965 ) ? ( n49516 ) : ( n49518 ) ;
assign n49520 =  ( n1930 ) ? ( n49515 ) : ( n49519 ) ;
assign n49521 =  ( n879 ) ? ( n49510 ) : ( n49520 ) ;
assign n49522 =  ( n172 ) ? ( n28474 ) : ( VREG_6_6 ) ;
assign n49523 =  ( n170 ) ? ( n28473 ) : ( n49522 ) ;
assign n49524 =  ( n168 ) ? ( n28472 ) : ( n49523 ) ;
assign n49525 =  ( n166 ) ? ( n28471 ) : ( n49524 ) ;
assign n49526 =  ( n162 ) ? ( n28470 ) : ( n49525 ) ;
assign n49527 =  ( n172 ) ? ( n28484 ) : ( VREG_6_6 ) ;
assign n49528 =  ( n170 ) ? ( n28483 ) : ( n49527 ) ;
assign n49529 =  ( n168 ) ? ( n28482 ) : ( n49528 ) ;
assign n49530 =  ( n166 ) ? ( n28481 ) : ( n49529 ) ;
assign n49531 =  ( n162 ) ? ( n28480 ) : ( n49530 ) ;
assign n49532 =  ( n28463 ) ? ( VREG_6_6 ) : ( n49531 ) ;
assign n49533 =  ( n3051 ) ? ( n49532 ) : ( VREG_6_6 ) ;
assign n49534 =  ( n3040 ) ? ( n49526 ) : ( n49533 ) ;
assign n49535 =  ( n192 ) ? ( VREG_6_6 ) : ( VREG_6_6 ) ;
assign n49536 =  ( n157 ) ? ( n49534 ) : ( n49535 ) ;
assign n49537 =  ( n6 ) ? ( n49521 ) : ( n49536 ) ;
assign n49538 =  ( n791 ) ? ( n49537 ) : ( VREG_6_6 ) ;
assign n49539 =  ( n148 ) ? ( n29541 ) : ( VREG_6_7 ) ;
assign n49540 =  ( n146 ) ? ( n29540 ) : ( n49539 ) ;
assign n49541 =  ( n144 ) ? ( n29539 ) : ( n49540 ) ;
assign n49542 =  ( n142 ) ? ( n29538 ) : ( n49541 ) ;
assign n49543 =  ( n10 ) ? ( n29537 ) : ( n49542 ) ;
assign n49544 =  ( n148 ) ? ( n30575 ) : ( VREG_6_7 ) ;
assign n49545 =  ( n146 ) ? ( n30574 ) : ( n49544 ) ;
assign n49546 =  ( n144 ) ? ( n30573 ) : ( n49545 ) ;
assign n49547 =  ( n142 ) ? ( n30572 ) : ( n49546 ) ;
assign n49548 =  ( n10 ) ? ( n30571 ) : ( n49547 ) ;
assign n49549 =  ( n30582 ) ? ( VREG_6_7 ) : ( n49543 ) ;
assign n49550 =  ( n30582 ) ? ( VREG_6_7 ) : ( n49548 ) ;
assign n49551 =  ( n3034 ) ? ( n49550 ) : ( VREG_6_7 ) ;
assign n49552 =  ( n2965 ) ? ( n49549 ) : ( n49551 ) ;
assign n49553 =  ( n1930 ) ? ( n49548 ) : ( n49552 ) ;
assign n49554 =  ( n879 ) ? ( n49543 ) : ( n49553 ) ;
assign n49555 =  ( n172 ) ? ( n30593 ) : ( VREG_6_7 ) ;
assign n49556 =  ( n170 ) ? ( n30592 ) : ( n49555 ) ;
assign n49557 =  ( n168 ) ? ( n30591 ) : ( n49556 ) ;
assign n49558 =  ( n166 ) ? ( n30590 ) : ( n49557 ) ;
assign n49559 =  ( n162 ) ? ( n30589 ) : ( n49558 ) ;
assign n49560 =  ( n172 ) ? ( n30603 ) : ( VREG_6_7 ) ;
assign n49561 =  ( n170 ) ? ( n30602 ) : ( n49560 ) ;
assign n49562 =  ( n168 ) ? ( n30601 ) : ( n49561 ) ;
assign n49563 =  ( n166 ) ? ( n30600 ) : ( n49562 ) ;
assign n49564 =  ( n162 ) ? ( n30599 ) : ( n49563 ) ;
assign n49565 =  ( n30582 ) ? ( VREG_6_7 ) : ( n49564 ) ;
assign n49566 =  ( n3051 ) ? ( n49565 ) : ( VREG_6_7 ) ;
assign n49567 =  ( n3040 ) ? ( n49559 ) : ( n49566 ) ;
assign n49568 =  ( n192 ) ? ( VREG_6_7 ) : ( VREG_6_7 ) ;
assign n49569 =  ( n157 ) ? ( n49567 ) : ( n49568 ) ;
assign n49570 =  ( n6 ) ? ( n49554 ) : ( n49569 ) ;
assign n49571 =  ( n791 ) ? ( n49570 ) : ( VREG_6_7 ) ;
assign n49572 =  ( n148 ) ? ( n31660 ) : ( VREG_6_8 ) ;
assign n49573 =  ( n146 ) ? ( n31659 ) : ( n49572 ) ;
assign n49574 =  ( n144 ) ? ( n31658 ) : ( n49573 ) ;
assign n49575 =  ( n142 ) ? ( n31657 ) : ( n49574 ) ;
assign n49576 =  ( n10 ) ? ( n31656 ) : ( n49575 ) ;
assign n49577 =  ( n148 ) ? ( n32694 ) : ( VREG_6_8 ) ;
assign n49578 =  ( n146 ) ? ( n32693 ) : ( n49577 ) ;
assign n49579 =  ( n144 ) ? ( n32692 ) : ( n49578 ) ;
assign n49580 =  ( n142 ) ? ( n32691 ) : ( n49579 ) ;
assign n49581 =  ( n10 ) ? ( n32690 ) : ( n49580 ) ;
assign n49582 =  ( n32701 ) ? ( VREG_6_8 ) : ( n49576 ) ;
assign n49583 =  ( n32701 ) ? ( VREG_6_8 ) : ( n49581 ) ;
assign n49584 =  ( n3034 ) ? ( n49583 ) : ( VREG_6_8 ) ;
assign n49585 =  ( n2965 ) ? ( n49582 ) : ( n49584 ) ;
assign n49586 =  ( n1930 ) ? ( n49581 ) : ( n49585 ) ;
assign n49587 =  ( n879 ) ? ( n49576 ) : ( n49586 ) ;
assign n49588 =  ( n172 ) ? ( n32712 ) : ( VREG_6_8 ) ;
assign n49589 =  ( n170 ) ? ( n32711 ) : ( n49588 ) ;
assign n49590 =  ( n168 ) ? ( n32710 ) : ( n49589 ) ;
assign n49591 =  ( n166 ) ? ( n32709 ) : ( n49590 ) ;
assign n49592 =  ( n162 ) ? ( n32708 ) : ( n49591 ) ;
assign n49593 =  ( n172 ) ? ( n32722 ) : ( VREG_6_8 ) ;
assign n49594 =  ( n170 ) ? ( n32721 ) : ( n49593 ) ;
assign n49595 =  ( n168 ) ? ( n32720 ) : ( n49594 ) ;
assign n49596 =  ( n166 ) ? ( n32719 ) : ( n49595 ) ;
assign n49597 =  ( n162 ) ? ( n32718 ) : ( n49596 ) ;
assign n49598 =  ( n32701 ) ? ( VREG_6_8 ) : ( n49597 ) ;
assign n49599 =  ( n3051 ) ? ( n49598 ) : ( VREG_6_8 ) ;
assign n49600 =  ( n3040 ) ? ( n49592 ) : ( n49599 ) ;
assign n49601 =  ( n192 ) ? ( VREG_6_8 ) : ( VREG_6_8 ) ;
assign n49602 =  ( n157 ) ? ( n49600 ) : ( n49601 ) ;
assign n49603 =  ( n6 ) ? ( n49587 ) : ( n49602 ) ;
assign n49604 =  ( n791 ) ? ( n49603 ) : ( VREG_6_8 ) ;
assign n49605 =  ( n148 ) ? ( n33779 ) : ( VREG_6_9 ) ;
assign n49606 =  ( n146 ) ? ( n33778 ) : ( n49605 ) ;
assign n49607 =  ( n144 ) ? ( n33777 ) : ( n49606 ) ;
assign n49608 =  ( n142 ) ? ( n33776 ) : ( n49607 ) ;
assign n49609 =  ( n10 ) ? ( n33775 ) : ( n49608 ) ;
assign n49610 =  ( n148 ) ? ( n34813 ) : ( VREG_6_9 ) ;
assign n49611 =  ( n146 ) ? ( n34812 ) : ( n49610 ) ;
assign n49612 =  ( n144 ) ? ( n34811 ) : ( n49611 ) ;
assign n49613 =  ( n142 ) ? ( n34810 ) : ( n49612 ) ;
assign n49614 =  ( n10 ) ? ( n34809 ) : ( n49613 ) ;
assign n49615 =  ( n34820 ) ? ( VREG_6_9 ) : ( n49609 ) ;
assign n49616 =  ( n34820 ) ? ( VREG_6_9 ) : ( n49614 ) ;
assign n49617 =  ( n3034 ) ? ( n49616 ) : ( VREG_6_9 ) ;
assign n49618 =  ( n2965 ) ? ( n49615 ) : ( n49617 ) ;
assign n49619 =  ( n1930 ) ? ( n49614 ) : ( n49618 ) ;
assign n49620 =  ( n879 ) ? ( n49609 ) : ( n49619 ) ;
assign n49621 =  ( n172 ) ? ( n34831 ) : ( VREG_6_9 ) ;
assign n49622 =  ( n170 ) ? ( n34830 ) : ( n49621 ) ;
assign n49623 =  ( n168 ) ? ( n34829 ) : ( n49622 ) ;
assign n49624 =  ( n166 ) ? ( n34828 ) : ( n49623 ) ;
assign n49625 =  ( n162 ) ? ( n34827 ) : ( n49624 ) ;
assign n49626 =  ( n172 ) ? ( n34841 ) : ( VREG_6_9 ) ;
assign n49627 =  ( n170 ) ? ( n34840 ) : ( n49626 ) ;
assign n49628 =  ( n168 ) ? ( n34839 ) : ( n49627 ) ;
assign n49629 =  ( n166 ) ? ( n34838 ) : ( n49628 ) ;
assign n49630 =  ( n162 ) ? ( n34837 ) : ( n49629 ) ;
assign n49631 =  ( n34820 ) ? ( VREG_6_9 ) : ( n49630 ) ;
assign n49632 =  ( n3051 ) ? ( n49631 ) : ( VREG_6_9 ) ;
assign n49633 =  ( n3040 ) ? ( n49625 ) : ( n49632 ) ;
assign n49634 =  ( n192 ) ? ( VREG_6_9 ) : ( VREG_6_9 ) ;
assign n49635 =  ( n157 ) ? ( n49633 ) : ( n49634 ) ;
assign n49636 =  ( n6 ) ? ( n49620 ) : ( n49635 ) ;
assign n49637 =  ( n791 ) ? ( n49636 ) : ( VREG_6_9 ) ;
assign n49638 =  ( n148 ) ? ( n1924 ) : ( VREG_7_0 ) ;
assign n49639 =  ( n146 ) ? ( n1923 ) : ( n49638 ) ;
assign n49640 =  ( n144 ) ? ( n1922 ) : ( n49639 ) ;
assign n49641 =  ( n142 ) ? ( n1921 ) : ( n49640 ) ;
assign n49642 =  ( n10 ) ? ( n1920 ) : ( n49641 ) ;
assign n49643 =  ( n148 ) ? ( n2959 ) : ( VREG_7_0 ) ;
assign n49644 =  ( n146 ) ? ( n2958 ) : ( n49643 ) ;
assign n49645 =  ( n144 ) ? ( n2957 ) : ( n49644 ) ;
assign n49646 =  ( n142 ) ? ( n2956 ) : ( n49645 ) ;
assign n49647 =  ( n10 ) ? ( n2955 ) : ( n49646 ) ;
assign n49648 =  ( n3032 ) ? ( VREG_7_0 ) : ( n49642 ) ;
assign n49649 =  ( n3032 ) ? ( VREG_7_0 ) : ( n49647 ) ;
assign n49650 =  ( n3034 ) ? ( n49649 ) : ( VREG_7_0 ) ;
assign n49651 =  ( n2965 ) ? ( n49648 ) : ( n49650 ) ;
assign n49652 =  ( n1930 ) ? ( n49647 ) : ( n49651 ) ;
assign n49653 =  ( n879 ) ? ( n49642 ) : ( n49652 ) ;
assign n49654 =  ( n172 ) ? ( n3045 ) : ( VREG_7_0 ) ;
assign n49655 =  ( n170 ) ? ( n3044 ) : ( n49654 ) ;
assign n49656 =  ( n168 ) ? ( n3043 ) : ( n49655 ) ;
assign n49657 =  ( n166 ) ? ( n3042 ) : ( n49656 ) ;
assign n49658 =  ( n162 ) ? ( n3041 ) : ( n49657 ) ;
assign n49659 =  ( n172 ) ? ( n3056 ) : ( VREG_7_0 ) ;
assign n49660 =  ( n170 ) ? ( n3055 ) : ( n49659 ) ;
assign n49661 =  ( n168 ) ? ( n3054 ) : ( n49660 ) ;
assign n49662 =  ( n166 ) ? ( n3053 ) : ( n49661 ) ;
assign n49663 =  ( n162 ) ? ( n3052 ) : ( n49662 ) ;
assign n49664 =  ( n3032 ) ? ( VREG_7_0 ) : ( n49663 ) ;
assign n49665 =  ( n3051 ) ? ( n49664 ) : ( VREG_7_0 ) ;
assign n49666 =  ( n3040 ) ? ( n49658 ) : ( n49665 ) ;
assign n49667 =  ( n192 ) ? ( VREG_7_0 ) : ( VREG_7_0 ) ;
assign n49668 =  ( n157 ) ? ( n49666 ) : ( n49667 ) ;
assign n49669 =  ( n6 ) ? ( n49653 ) : ( n49668 ) ;
assign n49670 =  ( n813 ) ? ( n49669 ) : ( VREG_7_0 ) ;
assign n49671 =  ( n148 ) ? ( n4113 ) : ( VREG_7_1 ) ;
assign n49672 =  ( n146 ) ? ( n4112 ) : ( n49671 ) ;
assign n49673 =  ( n144 ) ? ( n4111 ) : ( n49672 ) ;
assign n49674 =  ( n142 ) ? ( n4110 ) : ( n49673 ) ;
assign n49675 =  ( n10 ) ? ( n4109 ) : ( n49674 ) ;
assign n49676 =  ( n148 ) ? ( n5147 ) : ( VREG_7_1 ) ;
assign n49677 =  ( n146 ) ? ( n5146 ) : ( n49676 ) ;
assign n49678 =  ( n144 ) ? ( n5145 ) : ( n49677 ) ;
assign n49679 =  ( n142 ) ? ( n5144 ) : ( n49678 ) ;
assign n49680 =  ( n10 ) ? ( n5143 ) : ( n49679 ) ;
assign n49681 =  ( n5154 ) ? ( VREG_7_1 ) : ( n49675 ) ;
assign n49682 =  ( n5154 ) ? ( VREG_7_1 ) : ( n49680 ) ;
assign n49683 =  ( n3034 ) ? ( n49682 ) : ( VREG_7_1 ) ;
assign n49684 =  ( n2965 ) ? ( n49681 ) : ( n49683 ) ;
assign n49685 =  ( n1930 ) ? ( n49680 ) : ( n49684 ) ;
assign n49686 =  ( n879 ) ? ( n49675 ) : ( n49685 ) ;
assign n49687 =  ( n172 ) ? ( n5165 ) : ( VREG_7_1 ) ;
assign n49688 =  ( n170 ) ? ( n5164 ) : ( n49687 ) ;
assign n49689 =  ( n168 ) ? ( n5163 ) : ( n49688 ) ;
assign n49690 =  ( n166 ) ? ( n5162 ) : ( n49689 ) ;
assign n49691 =  ( n162 ) ? ( n5161 ) : ( n49690 ) ;
assign n49692 =  ( n172 ) ? ( n5175 ) : ( VREG_7_1 ) ;
assign n49693 =  ( n170 ) ? ( n5174 ) : ( n49692 ) ;
assign n49694 =  ( n168 ) ? ( n5173 ) : ( n49693 ) ;
assign n49695 =  ( n166 ) ? ( n5172 ) : ( n49694 ) ;
assign n49696 =  ( n162 ) ? ( n5171 ) : ( n49695 ) ;
assign n49697 =  ( n5154 ) ? ( VREG_7_1 ) : ( n49696 ) ;
assign n49698 =  ( n3051 ) ? ( n49697 ) : ( VREG_7_1 ) ;
assign n49699 =  ( n3040 ) ? ( n49691 ) : ( n49698 ) ;
assign n49700 =  ( n192 ) ? ( VREG_7_1 ) : ( VREG_7_1 ) ;
assign n49701 =  ( n157 ) ? ( n49699 ) : ( n49700 ) ;
assign n49702 =  ( n6 ) ? ( n49686 ) : ( n49701 ) ;
assign n49703 =  ( n813 ) ? ( n49702 ) : ( VREG_7_1 ) ;
assign n49704 =  ( n148 ) ? ( n6232 ) : ( VREG_7_10 ) ;
assign n49705 =  ( n146 ) ? ( n6231 ) : ( n49704 ) ;
assign n49706 =  ( n144 ) ? ( n6230 ) : ( n49705 ) ;
assign n49707 =  ( n142 ) ? ( n6229 ) : ( n49706 ) ;
assign n49708 =  ( n10 ) ? ( n6228 ) : ( n49707 ) ;
assign n49709 =  ( n148 ) ? ( n7266 ) : ( VREG_7_10 ) ;
assign n49710 =  ( n146 ) ? ( n7265 ) : ( n49709 ) ;
assign n49711 =  ( n144 ) ? ( n7264 ) : ( n49710 ) ;
assign n49712 =  ( n142 ) ? ( n7263 ) : ( n49711 ) ;
assign n49713 =  ( n10 ) ? ( n7262 ) : ( n49712 ) ;
assign n49714 =  ( n7273 ) ? ( VREG_7_10 ) : ( n49708 ) ;
assign n49715 =  ( n7273 ) ? ( VREG_7_10 ) : ( n49713 ) ;
assign n49716 =  ( n3034 ) ? ( n49715 ) : ( VREG_7_10 ) ;
assign n49717 =  ( n2965 ) ? ( n49714 ) : ( n49716 ) ;
assign n49718 =  ( n1930 ) ? ( n49713 ) : ( n49717 ) ;
assign n49719 =  ( n879 ) ? ( n49708 ) : ( n49718 ) ;
assign n49720 =  ( n172 ) ? ( n7284 ) : ( VREG_7_10 ) ;
assign n49721 =  ( n170 ) ? ( n7283 ) : ( n49720 ) ;
assign n49722 =  ( n168 ) ? ( n7282 ) : ( n49721 ) ;
assign n49723 =  ( n166 ) ? ( n7281 ) : ( n49722 ) ;
assign n49724 =  ( n162 ) ? ( n7280 ) : ( n49723 ) ;
assign n49725 =  ( n172 ) ? ( n7294 ) : ( VREG_7_10 ) ;
assign n49726 =  ( n170 ) ? ( n7293 ) : ( n49725 ) ;
assign n49727 =  ( n168 ) ? ( n7292 ) : ( n49726 ) ;
assign n49728 =  ( n166 ) ? ( n7291 ) : ( n49727 ) ;
assign n49729 =  ( n162 ) ? ( n7290 ) : ( n49728 ) ;
assign n49730 =  ( n7273 ) ? ( VREG_7_10 ) : ( n49729 ) ;
assign n49731 =  ( n3051 ) ? ( n49730 ) : ( VREG_7_10 ) ;
assign n49732 =  ( n3040 ) ? ( n49724 ) : ( n49731 ) ;
assign n49733 =  ( n192 ) ? ( VREG_7_10 ) : ( VREG_7_10 ) ;
assign n49734 =  ( n157 ) ? ( n49732 ) : ( n49733 ) ;
assign n49735 =  ( n6 ) ? ( n49719 ) : ( n49734 ) ;
assign n49736 =  ( n813 ) ? ( n49735 ) : ( VREG_7_10 ) ;
assign n49737 =  ( n148 ) ? ( n8351 ) : ( VREG_7_11 ) ;
assign n49738 =  ( n146 ) ? ( n8350 ) : ( n49737 ) ;
assign n49739 =  ( n144 ) ? ( n8349 ) : ( n49738 ) ;
assign n49740 =  ( n142 ) ? ( n8348 ) : ( n49739 ) ;
assign n49741 =  ( n10 ) ? ( n8347 ) : ( n49740 ) ;
assign n49742 =  ( n148 ) ? ( n9385 ) : ( VREG_7_11 ) ;
assign n49743 =  ( n146 ) ? ( n9384 ) : ( n49742 ) ;
assign n49744 =  ( n144 ) ? ( n9383 ) : ( n49743 ) ;
assign n49745 =  ( n142 ) ? ( n9382 ) : ( n49744 ) ;
assign n49746 =  ( n10 ) ? ( n9381 ) : ( n49745 ) ;
assign n49747 =  ( n9392 ) ? ( VREG_7_11 ) : ( n49741 ) ;
assign n49748 =  ( n9392 ) ? ( VREG_7_11 ) : ( n49746 ) ;
assign n49749 =  ( n3034 ) ? ( n49748 ) : ( VREG_7_11 ) ;
assign n49750 =  ( n2965 ) ? ( n49747 ) : ( n49749 ) ;
assign n49751 =  ( n1930 ) ? ( n49746 ) : ( n49750 ) ;
assign n49752 =  ( n879 ) ? ( n49741 ) : ( n49751 ) ;
assign n49753 =  ( n172 ) ? ( n9403 ) : ( VREG_7_11 ) ;
assign n49754 =  ( n170 ) ? ( n9402 ) : ( n49753 ) ;
assign n49755 =  ( n168 ) ? ( n9401 ) : ( n49754 ) ;
assign n49756 =  ( n166 ) ? ( n9400 ) : ( n49755 ) ;
assign n49757 =  ( n162 ) ? ( n9399 ) : ( n49756 ) ;
assign n49758 =  ( n172 ) ? ( n9413 ) : ( VREG_7_11 ) ;
assign n49759 =  ( n170 ) ? ( n9412 ) : ( n49758 ) ;
assign n49760 =  ( n168 ) ? ( n9411 ) : ( n49759 ) ;
assign n49761 =  ( n166 ) ? ( n9410 ) : ( n49760 ) ;
assign n49762 =  ( n162 ) ? ( n9409 ) : ( n49761 ) ;
assign n49763 =  ( n9392 ) ? ( VREG_7_11 ) : ( n49762 ) ;
assign n49764 =  ( n3051 ) ? ( n49763 ) : ( VREG_7_11 ) ;
assign n49765 =  ( n3040 ) ? ( n49757 ) : ( n49764 ) ;
assign n49766 =  ( n192 ) ? ( VREG_7_11 ) : ( VREG_7_11 ) ;
assign n49767 =  ( n157 ) ? ( n49765 ) : ( n49766 ) ;
assign n49768 =  ( n6 ) ? ( n49752 ) : ( n49767 ) ;
assign n49769 =  ( n813 ) ? ( n49768 ) : ( VREG_7_11 ) ;
assign n49770 =  ( n148 ) ? ( n10470 ) : ( VREG_7_12 ) ;
assign n49771 =  ( n146 ) ? ( n10469 ) : ( n49770 ) ;
assign n49772 =  ( n144 ) ? ( n10468 ) : ( n49771 ) ;
assign n49773 =  ( n142 ) ? ( n10467 ) : ( n49772 ) ;
assign n49774 =  ( n10 ) ? ( n10466 ) : ( n49773 ) ;
assign n49775 =  ( n148 ) ? ( n11504 ) : ( VREG_7_12 ) ;
assign n49776 =  ( n146 ) ? ( n11503 ) : ( n49775 ) ;
assign n49777 =  ( n144 ) ? ( n11502 ) : ( n49776 ) ;
assign n49778 =  ( n142 ) ? ( n11501 ) : ( n49777 ) ;
assign n49779 =  ( n10 ) ? ( n11500 ) : ( n49778 ) ;
assign n49780 =  ( n11511 ) ? ( VREG_7_12 ) : ( n49774 ) ;
assign n49781 =  ( n11511 ) ? ( VREG_7_12 ) : ( n49779 ) ;
assign n49782 =  ( n3034 ) ? ( n49781 ) : ( VREG_7_12 ) ;
assign n49783 =  ( n2965 ) ? ( n49780 ) : ( n49782 ) ;
assign n49784 =  ( n1930 ) ? ( n49779 ) : ( n49783 ) ;
assign n49785 =  ( n879 ) ? ( n49774 ) : ( n49784 ) ;
assign n49786 =  ( n172 ) ? ( n11522 ) : ( VREG_7_12 ) ;
assign n49787 =  ( n170 ) ? ( n11521 ) : ( n49786 ) ;
assign n49788 =  ( n168 ) ? ( n11520 ) : ( n49787 ) ;
assign n49789 =  ( n166 ) ? ( n11519 ) : ( n49788 ) ;
assign n49790 =  ( n162 ) ? ( n11518 ) : ( n49789 ) ;
assign n49791 =  ( n172 ) ? ( n11532 ) : ( VREG_7_12 ) ;
assign n49792 =  ( n170 ) ? ( n11531 ) : ( n49791 ) ;
assign n49793 =  ( n168 ) ? ( n11530 ) : ( n49792 ) ;
assign n49794 =  ( n166 ) ? ( n11529 ) : ( n49793 ) ;
assign n49795 =  ( n162 ) ? ( n11528 ) : ( n49794 ) ;
assign n49796 =  ( n11511 ) ? ( VREG_7_12 ) : ( n49795 ) ;
assign n49797 =  ( n3051 ) ? ( n49796 ) : ( VREG_7_12 ) ;
assign n49798 =  ( n3040 ) ? ( n49790 ) : ( n49797 ) ;
assign n49799 =  ( n192 ) ? ( VREG_7_12 ) : ( VREG_7_12 ) ;
assign n49800 =  ( n157 ) ? ( n49798 ) : ( n49799 ) ;
assign n49801 =  ( n6 ) ? ( n49785 ) : ( n49800 ) ;
assign n49802 =  ( n813 ) ? ( n49801 ) : ( VREG_7_12 ) ;
assign n49803 =  ( n148 ) ? ( n12589 ) : ( VREG_7_13 ) ;
assign n49804 =  ( n146 ) ? ( n12588 ) : ( n49803 ) ;
assign n49805 =  ( n144 ) ? ( n12587 ) : ( n49804 ) ;
assign n49806 =  ( n142 ) ? ( n12586 ) : ( n49805 ) ;
assign n49807 =  ( n10 ) ? ( n12585 ) : ( n49806 ) ;
assign n49808 =  ( n148 ) ? ( n13623 ) : ( VREG_7_13 ) ;
assign n49809 =  ( n146 ) ? ( n13622 ) : ( n49808 ) ;
assign n49810 =  ( n144 ) ? ( n13621 ) : ( n49809 ) ;
assign n49811 =  ( n142 ) ? ( n13620 ) : ( n49810 ) ;
assign n49812 =  ( n10 ) ? ( n13619 ) : ( n49811 ) ;
assign n49813 =  ( n13630 ) ? ( VREG_7_13 ) : ( n49807 ) ;
assign n49814 =  ( n13630 ) ? ( VREG_7_13 ) : ( n49812 ) ;
assign n49815 =  ( n3034 ) ? ( n49814 ) : ( VREG_7_13 ) ;
assign n49816 =  ( n2965 ) ? ( n49813 ) : ( n49815 ) ;
assign n49817 =  ( n1930 ) ? ( n49812 ) : ( n49816 ) ;
assign n49818 =  ( n879 ) ? ( n49807 ) : ( n49817 ) ;
assign n49819 =  ( n172 ) ? ( n13641 ) : ( VREG_7_13 ) ;
assign n49820 =  ( n170 ) ? ( n13640 ) : ( n49819 ) ;
assign n49821 =  ( n168 ) ? ( n13639 ) : ( n49820 ) ;
assign n49822 =  ( n166 ) ? ( n13638 ) : ( n49821 ) ;
assign n49823 =  ( n162 ) ? ( n13637 ) : ( n49822 ) ;
assign n49824 =  ( n172 ) ? ( n13651 ) : ( VREG_7_13 ) ;
assign n49825 =  ( n170 ) ? ( n13650 ) : ( n49824 ) ;
assign n49826 =  ( n168 ) ? ( n13649 ) : ( n49825 ) ;
assign n49827 =  ( n166 ) ? ( n13648 ) : ( n49826 ) ;
assign n49828 =  ( n162 ) ? ( n13647 ) : ( n49827 ) ;
assign n49829 =  ( n13630 ) ? ( VREG_7_13 ) : ( n49828 ) ;
assign n49830 =  ( n3051 ) ? ( n49829 ) : ( VREG_7_13 ) ;
assign n49831 =  ( n3040 ) ? ( n49823 ) : ( n49830 ) ;
assign n49832 =  ( n192 ) ? ( VREG_7_13 ) : ( VREG_7_13 ) ;
assign n49833 =  ( n157 ) ? ( n49831 ) : ( n49832 ) ;
assign n49834 =  ( n6 ) ? ( n49818 ) : ( n49833 ) ;
assign n49835 =  ( n813 ) ? ( n49834 ) : ( VREG_7_13 ) ;
assign n49836 =  ( n148 ) ? ( n14708 ) : ( VREG_7_14 ) ;
assign n49837 =  ( n146 ) ? ( n14707 ) : ( n49836 ) ;
assign n49838 =  ( n144 ) ? ( n14706 ) : ( n49837 ) ;
assign n49839 =  ( n142 ) ? ( n14705 ) : ( n49838 ) ;
assign n49840 =  ( n10 ) ? ( n14704 ) : ( n49839 ) ;
assign n49841 =  ( n148 ) ? ( n15742 ) : ( VREG_7_14 ) ;
assign n49842 =  ( n146 ) ? ( n15741 ) : ( n49841 ) ;
assign n49843 =  ( n144 ) ? ( n15740 ) : ( n49842 ) ;
assign n49844 =  ( n142 ) ? ( n15739 ) : ( n49843 ) ;
assign n49845 =  ( n10 ) ? ( n15738 ) : ( n49844 ) ;
assign n49846 =  ( n15749 ) ? ( VREG_7_14 ) : ( n49840 ) ;
assign n49847 =  ( n15749 ) ? ( VREG_7_14 ) : ( n49845 ) ;
assign n49848 =  ( n3034 ) ? ( n49847 ) : ( VREG_7_14 ) ;
assign n49849 =  ( n2965 ) ? ( n49846 ) : ( n49848 ) ;
assign n49850 =  ( n1930 ) ? ( n49845 ) : ( n49849 ) ;
assign n49851 =  ( n879 ) ? ( n49840 ) : ( n49850 ) ;
assign n49852 =  ( n172 ) ? ( n15760 ) : ( VREG_7_14 ) ;
assign n49853 =  ( n170 ) ? ( n15759 ) : ( n49852 ) ;
assign n49854 =  ( n168 ) ? ( n15758 ) : ( n49853 ) ;
assign n49855 =  ( n166 ) ? ( n15757 ) : ( n49854 ) ;
assign n49856 =  ( n162 ) ? ( n15756 ) : ( n49855 ) ;
assign n49857 =  ( n172 ) ? ( n15770 ) : ( VREG_7_14 ) ;
assign n49858 =  ( n170 ) ? ( n15769 ) : ( n49857 ) ;
assign n49859 =  ( n168 ) ? ( n15768 ) : ( n49858 ) ;
assign n49860 =  ( n166 ) ? ( n15767 ) : ( n49859 ) ;
assign n49861 =  ( n162 ) ? ( n15766 ) : ( n49860 ) ;
assign n49862 =  ( n15749 ) ? ( VREG_7_14 ) : ( n49861 ) ;
assign n49863 =  ( n3051 ) ? ( n49862 ) : ( VREG_7_14 ) ;
assign n49864 =  ( n3040 ) ? ( n49856 ) : ( n49863 ) ;
assign n49865 =  ( n192 ) ? ( VREG_7_14 ) : ( VREG_7_14 ) ;
assign n49866 =  ( n157 ) ? ( n49864 ) : ( n49865 ) ;
assign n49867 =  ( n6 ) ? ( n49851 ) : ( n49866 ) ;
assign n49868 =  ( n813 ) ? ( n49867 ) : ( VREG_7_14 ) ;
assign n49869 =  ( n148 ) ? ( n16827 ) : ( VREG_7_15 ) ;
assign n49870 =  ( n146 ) ? ( n16826 ) : ( n49869 ) ;
assign n49871 =  ( n144 ) ? ( n16825 ) : ( n49870 ) ;
assign n49872 =  ( n142 ) ? ( n16824 ) : ( n49871 ) ;
assign n49873 =  ( n10 ) ? ( n16823 ) : ( n49872 ) ;
assign n49874 =  ( n148 ) ? ( n17861 ) : ( VREG_7_15 ) ;
assign n49875 =  ( n146 ) ? ( n17860 ) : ( n49874 ) ;
assign n49876 =  ( n144 ) ? ( n17859 ) : ( n49875 ) ;
assign n49877 =  ( n142 ) ? ( n17858 ) : ( n49876 ) ;
assign n49878 =  ( n10 ) ? ( n17857 ) : ( n49877 ) ;
assign n49879 =  ( n17868 ) ? ( VREG_7_15 ) : ( n49873 ) ;
assign n49880 =  ( n17868 ) ? ( VREG_7_15 ) : ( n49878 ) ;
assign n49881 =  ( n3034 ) ? ( n49880 ) : ( VREG_7_15 ) ;
assign n49882 =  ( n2965 ) ? ( n49879 ) : ( n49881 ) ;
assign n49883 =  ( n1930 ) ? ( n49878 ) : ( n49882 ) ;
assign n49884 =  ( n879 ) ? ( n49873 ) : ( n49883 ) ;
assign n49885 =  ( n172 ) ? ( n17879 ) : ( VREG_7_15 ) ;
assign n49886 =  ( n170 ) ? ( n17878 ) : ( n49885 ) ;
assign n49887 =  ( n168 ) ? ( n17877 ) : ( n49886 ) ;
assign n49888 =  ( n166 ) ? ( n17876 ) : ( n49887 ) ;
assign n49889 =  ( n162 ) ? ( n17875 ) : ( n49888 ) ;
assign n49890 =  ( n172 ) ? ( n17889 ) : ( VREG_7_15 ) ;
assign n49891 =  ( n170 ) ? ( n17888 ) : ( n49890 ) ;
assign n49892 =  ( n168 ) ? ( n17887 ) : ( n49891 ) ;
assign n49893 =  ( n166 ) ? ( n17886 ) : ( n49892 ) ;
assign n49894 =  ( n162 ) ? ( n17885 ) : ( n49893 ) ;
assign n49895 =  ( n17868 ) ? ( VREG_7_15 ) : ( n49894 ) ;
assign n49896 =  ( n3051 ) ? ( n49895 ) : ( VREG_7_15 ) ;
assign n49897 =  ( n3040 ) ? ( n49889 ) : ( n49896 ) ;
assign n49898 =  ( n192 ) ? ( VREG_7_15 ) : ( VREG_7_15 ) ;
assign n49899 =  ( n157 ) ? ( n49897 ) : ( n49898 ) ;
assign n49900 =  ( n6 ) ? ( n49884 ) : ( n49899 ) ;
assign n49901 =  ( n813 ) ? ( n49900 ) : ( VREG_7_15 ) ;
assign n49902 =  ( n148 ) ? ( n18946 ) : ( VREG_7_2 ) ;
assign n49903 =  ( n146 ) ? ( n18945 ) : ( n49902 ) ;
assign n49904 =  ( n144 ) ? ( n18944 ) : ( n49903 ) ;
assign n49905 =  ( n142 ) ? ( n18943 ) : ( n49904 ) ;
assign n49906 =  ( n10 ) ? ( n18942 ) : ( n49905 ) ;
assign n49907 =  ( n148 ) ? ( n19980 ) : ( VREG_7_2 ) ;
assign n49908 =  ( n146 ) ? ( n19979 ) : ( n49907 ) ;
assign n49909 =  ( n144 ) ? ( n19978 ) : ( n49908 ) ;
assign n49910 =  ( n142 ) ? ( n19977 ) : ( n49909 ) ;
assign n49911 =  ( n10 ) ? ( n19976 ) : ( n49910 ) ;
assign n49912 =  ( n19987 ) ? ( VREG_7_2 ) : ( n49906 ) ;
assign n49913 =  ( n19987 ) ? ( VREG_7_2 ) : ( n49911 ) ;
assign n49914 =  ( n3034 ) ? ( n49913 ) : ( VREG_7_2 ) ;
assign n49915 =  ( n2965 ) ? ( n49912 ) : ( n49914 ) ;
assign n49916 =  ( n1930 ) ? ( n49911 ) : ( n49915 ) ;
assign n49917 =  ( n879 ) ? ( n49906 ) : ( n49916 ) ;
assign n49918 =  ( n172 ) ? ( n19998 ) : ( VREG_7_2 ) ;
assign n49919 =  ( n170 ) ? ( n19997 ) : ( n49918 ) ;
assign n49920 =  ( n168 ) ? ( n19996 ) : ( n49919 ) ;
assign n49921 =  ( n166 ) ? ( n19995 ) : ( n49920 ) ;
assign n49922 =  ( n162 ) ? ( n19994 ) : ( n49921 ) ;
assign n49923 =  ( n172 ) ? ( n20008 ) : ( VREG_7_2 ) ;
assign n49924 =  ( n170 ) ? ( n20007 ) : ( n49923 ) ;
assign n49925 =  ( n168 ) ? ( n20006 ) : ( n49924 ) ;
assign n49926 =  ( n166 ) ? ( n20005 ) : ( n49925 ) ;
assign n49927 =  ( n162 ) ? ( n20004 ) : ( n49926 ) ;
assign n49928 =  ( n19987 ) ? ( VREG_7_2 ) : ( n49927 ) ;
assign n49929 =  ( n3051 ) ? ( n49928 ) : ( VREG_7_2 ) ;
assign n49930 =  ( n3040 ) ? ( n49922 ) : ( n49929 ) ;
assign n49931 =  ( n192 ) ? ( VREG_7_2 ) : ( VREG_7_2 ) ;
assign n49932 =  ( n157 ) ? ( n49930 ) : ( n49931 ) ;
assign n49933 =  ( n6 ) ? ( n49917 ) : ( n49932 ) ;
assign n49934 =  ( n813 ) ? ( n49933 ) : ( VREG_7_2 ) ;
assign n49935 =  ( n148 ) ? ( n21065 ) : ( VREG_7_3 ) ;
assign n49936 =  ( n146 ) ? ( n21064 ) : ( n49935 ) ;
assign n49937 =  ( n144 ) ? ( n21063 ) : ( n49936 ) ;
assign n49938 =  ( n142 ) ? ( n21062 ) : ( n49937 ) ;
assign n49939 =  ( n10 ) ? ( n21061 ) : ( n49938 ) ;
assign n49940 =  ( n148 ) ? ( n22099 ) : ( VREG_7_3 ) ;
assign n49941 =  ( n146 ) ? ( n22098 ) : ( n49940 ) ;
assign n49942 =  ( n144 ) ? ( n22097 ) : ( n49941 ) ;
assign n49943 =  ( n142 ) ? ( n22096 ) : ( n49942 ) ;
assign n49944 =  ( n10 ) ? ( n22095 ) : ( n49943 ) ;
assign n49945 =  ( n22106 ) ? ( VREG_7_3 ) : ( n49939 ) ;
assign n49946 =  ( n22106 ) ? ( VREG_7_3 ) : ( n49944 ) ;
assign n49947 =  ( n3034 ) ? ( n49946 ) : ( VREG_7_3 ) ;
assign n49948 =  ( n2965 ) ? ( n49945 ) : ( n49947 ) ;
assign n49949 =  ( n1930 ) ? ( n49944 ) : ( n49948 ) ;
assign n49950 =  ( n879 ) ? ( n49939 ) : ( n49949 ) ;
assign n49951 =  ( n172 ) ? ( n22117 ) : ( VREG_7_3 ) ;
assign n49952 =  ( n170 ) ? ( n22116 ) : ( n49951 ) ;
assign n49953 =  ( n168 ) ? ( n22115 ) : ( n49952 ) ;
assign n49954 =  ( n166 ) ? ( n22114 ) : ( n49953 ) ;
assign n49955 =  ( n162 ) ? ( n22113 ) : ( n49954 ) ;
assign n49956 =  ( n172 ) ? ( n22127 ) : ( VREG_7_3 ) ;
assign n49957 =  ( n170 ) ? ( n22126 ) : ( n49956 ) ;
assign n49958 =  ( n168 ) ? ( n22125 ) : ( n49957 ) ;
assign n49959 =  ( n166 ) ? ( n22124 ) : ( n49958 ) ;
assign n49960 =  ( n162 ) ? ( n22123 ) : ( n49959 ) ;
assign n49961 =  ( n22106 ) ? ( VREG_7_3 ) : ( n49960 ) ;
assign n49962 =  ( n3051 ) ? ( n49961 ) : ( VREG_7_3 ) ;
assign n49963 =  ( n3040 ) ? ( n49955 ) : ( n49962 ) ;
assign n49964 =  ( n192 ) ? ( VREG_7_3 ) : ( VREG_7_3 ) ;
assign n49965 =  ( n157 ) ? ( n49963 ) : ( n49964 ) ;
assign n49966 =  ( n6 ) ? ( n49950 ) : ( n49965 ) ;
assign n49967 =  ( n813 ) ? ( n49966 ) : ( VREG_7_3 ) ;
assign n49968 =  ( n148 ) ? ( n23184 ) : ( VREG_7_4 ) ;
assign n49969 =  ( n146 ) ? ( n23183 ) : ( n49968 ) ;
assign n49970 =  ( n144 ) ? ( n23182 ) : ( n49969 ) ;
assign n49971 =  ( n142 ) ? ( n23181 ) : ( n49970 ) ;
assign n49972 =  ( n10 ) ? ( n23180 ) : ( n49971 ) ;
assign n49973 =  ( n148 ) ? ( n24218 ) : ( VREG_7_4 ) ;
assign n49974 =  ( n146 ) ? ( n24217 ) : ( n49973 ) ;
assign n49975 =  ( n144 ) ? ( n24216 ) : ( n49974 ) ;
assign n49976 =  ( n142 ) ? ( n24215 ) : ( n49975 ) ;
assign n49977 =  ( n10 ) ? ( n24214 ) : ( n49976 ) ;
assign n49978 =  ( n24225 ) ? ( VREG_7_4 ) : ( n49972 ) ;
assign n49979 =  ( n24225 ) ? ( VREG_7_4 ) : ( n49977 ) ;
assign n49980 =  ( n3034 ) ? ( n49979 ) : ( VREG_7_4 ) ;
assign n49981 =  ( n2965 ) ? ( n49978 ) : ( n49980 ) ;
assign n49982 =  ( n1930 ) ? ( n49977 ) : ( n49981 ) ;
assign n49983 =  ( n879 ) ? ( n49972 ) : ( n49982 ) ;
assign n49984 =  ( n172 ) ? ( n24236 ) : ( VREG_7_4 ) ;
assign n49985 =  ( n170 ) ? ( n24235 ) : ( n49984 ) ;
assign n49986 =  ( n168 ) ? ( n24234 ) : ( n49985 ) ;
assign n49987 =  ( n166 ) ? ( n24233 ) : ( n49986 ) ;
assign n49988 =  ( n162 ) ? ( n24232 ) : ( n49987 ) ;
assign n49989 =  ( n172 ) ? ( n24246 ) : ( VREG_7_4 ) ;
assign n49990 =  ( n170 ) ? ( n24245 ) : ( n49989 ) ;
assign n49991 =  ( n168 ) ? ( n24244 ) : ( n49990 ) ;
assign n49992 =  ( n166 ) ? ( n24243 ) : ( n49991 ) ;
assign n49993 =  ( n162 ) ? ( n24242 ) : ( n49992 ) ;
assign n49994 =  ( n24225 ) ? ( VREG_7_4 ) : ( n49993 ) ;
assign n49995 =  ( n3051 ) ? ( n49994 ) : ( VREG_7_4 ) ;
assign n49996 =  ( n3040 ) ? ( n49988 ) : ( n49995 ) ;
assign n49997 =  ( n192 ) ? ( VREG_7_4 ) : ( VREG_7_4 ) ;
assign n49998 =  ( n157 ) ? ( n49996 ) : ( n49997 ) ;
assign n49999 =  ( n6 ) ? ( n49983 ) : ( n49998 ) ;
assign n50000 =  ( n813 ) ? ( n49999 ) : ( VREG_7_4 ) ;
assign n50001 =  ( n148 ) ? ( n25303 ) : ( VREG_7_5 ) ;
assign n50002 =  ( n146 ) ? ( n25302 ) : ( n50001 ) ;
assign n50003 =  ( n144 ) ? ( n25301 ) : ( n50002 ) ;
assign n50004 =  ( n142 ) ? ( n25300 ) : ( n50003 ) ;
assign n50005 =  ( n10 ) ? ( n25299 ) : ( n50004 ) ;
assign n50006 =  ( n148 ) ? ( n26337 ) : ( VREG_7_5 ) ;
assign n50007 =  ( n146 ) ? ( n26336 ) : ( n50006 ) ;
assign n50008 =  ( n144 ) ? ( n26335 ) : ( n50007 ) ;
assign n50009 =  ( n142 ) ? ( n26334 ) : ( n50008 ) ;
assign n50010 =  ( n10 ) ? ( n26333 ) : ( n50009 ) ;
assign n50011 =  ( n26344 ) ? ( VREG_7_5 ) : ( n50005 ) ;
assign n50012 =  ( n26344 ) ? ( VREG_7_5 ) : ( n50010 ) ;
assign n50013 =  ( n3034 ) ? ( n50012 ) : ( VREG_7_5 ) ;
assign n50014 =  ( n2965 ) ? ( n50011 ) : ( n50013 ) ;
assign n50015 =  ( n1930 ) ? ( n50010 ) : ( n50014 ) ;
assign n50016 =  ( n879 ) ? ( n50005 ) : ( n50015 ) ;
assign n50017 =  ( n172 ) ? ( n26355 ) : ( VREG_7_5 ) ;
assign n50018 =  ( n170 ) ? ( n26354 ) : ( n50017 ) ;
assign n50019 =  ( n168 ) ? ( n26353 ) : ( n50018 ) ;
assign n50020 =  ( n166 ) ? ( n26352 ) : ( n50019 ) ;
assign n50021 =  ( n162 ) ? ( n26351 ) : ( n50020 ) ;
assign n50022 =  ( n172 ) ? ( n26365 ) : ( VREG_7_5 ) ;
assign n50023 =  ( n170 ) ? ( n26364 ) : ( n50022 ) ;
assign n50024 =  ( n168 ) ? ( n26363 ) : ( n50023 ) ;
assign n50025 =  ( n166 ) ? ( n26362 ) : ( n50024 ) ;
assign n50026 =  ( n162 ) ? ( n26361 ) : ( n50025 ) ;
assign n50027 =  ( n26344 ) ? ( VREG_7_5 ) : ( n50026 ) ;
assign n50028 =  ( n3051 ) ? ( n50027 ) : ( VREG_7_5 ) ;
assign n50029 =  ( n3040 ) ? ( n50021 ) : ( n50028 ) ;
assign n50030 =  ( n192 ) ? ( VREG_7_5 ) : ( VREG_7_5 ) ;
assign n50031 =  ( n157 ) ? ( n50029 ) : ( n50030 ) ;
assign n50032 =  ( n6 ) ? ( n50016 ) : ( n50031 ) ;
assign n50033 =  ( n813 ) ? ( n50032 ) : ( VREG_7_5 ) ;
assign n50034 =  ( n148 ) ? ( n27422 ) : ( VREG_7_6 ) ;
assign n50035 =  ( n146 ) ? ( n27421 ) : ( n50034 ) ;
assign n50036 =  ( n144 ) ? ( n27420 ) : ( n50035 ) ;
assign n50037 =  ( n142 ) ? ( n27419 ) : ( n50036 ) ;
assign n50038 =  ( n10 ) ? ( n27418 ) : ( n50037 ) ;
assign n50039 =  ( n148 ) ? ( n28456 ) : ( VREG_7_6 ) ;
assign n50040 =  ( n146 ) ? ( n28455 ) : ( n50039 ) ;
assign n50041 =  ( n144 ) ? ( n28454 ) : ( n50040 ) ;
assign n50042 =  ( n142 ) ? ( n28453 ) : ( n50041 ) ;
assign n50043 =  ( n10 ) ? ( n28452 ) : ( n50042 ) ;
assign n50044 =  ( n28463 ) ? ( VREG_7_6 ) : ( n50038 ) ;
assign n50045 =  ( n28463 ) ? ( VREG_7_6 ) : ( n50043 ) ;
assign n50046 =  ( n3034 ) ? ( n50045 ) : ( VREG_7_6 ) ;
assign n50047 =  ( n2965 ) ? ( n50044 ) : ( n50046 ) ;
assign n50048 =  ( n1930 ) ? ( n50043 ) : ( n50047 ) ;
assign n50049 =  ( n879 ) ? ( n50038 ) : ( n50048 ) ;
assign n50050 =  ( n172 ) ? ( n28474 ) : ( VREG_7_6 ) ;
assign n50051 =  ( n170 ) ? ( n28473 ) : ( n50050 ) ;
assign n50052 =  ( n168 ) ? ( n28472 ) : ( n50051 ) ;
assign n50053 =  ( n166 ) ? ( n28471 ) : ( n50052 ) ;
assign n50054 =  ( n162 ) ? ( n28470 ) : ( n50053 ) ;
assign n50055 =  ( n172 ) ? ( n28484 ) : ( VREG_7_6 ) ;
assign n50056 =  ( n170 ) ? ( n28483 ) : ( n50055 ) ;
assign n50057 =  ( n168 ) ? ( n28482 ) : ( n50056 ) ;
assign n50058 =  ( n166 ) ? ( n28481 ) : ( n50057 ) ;
assign n50059 =  ( n162 ) ? ( n28480 ) : ( n50058 ) ;
assign n50060 =  ( n28463 ) ? ( VREG_7_6 ) : ( n50059 ) ;
assign n50061 =  ( n3051 ) ? ( n50060 ) : ( VREG_7_6 ) ;
assign n50062 =  ( n3040 ) ? ( n50054 ) : ( n50061 ) ;
assign n50063 =  ( n192 ) ? ( VREG_7_6 ) : ( VREG_7_6 ) ;
assign n50064 =  ( n157 ) ? ( n50062 ) : ( n50063 ) ;
assign n50065 =  ( n6 ) ? ( n50049 ) : ( n50064 ) ;
assign n50066 =  ( n813 ) ? ( n50065 ) : ( VREG_7_6 ) ;
assign n50067 =  ( n148 ) ? ( n29541 ) : ( VREG_7_7 ) ;
assign n50068 =  ( n146 ) ? ( n29540 ) : ( n50067 ) ;
assign n50069 =  ( n144 ) ? ( n29539 ) : ( n50068 ) ;
assign n50070 =  ( n142 ) ? ( n29538 ) : ( n50069 ) ;
assign n50071 =  ( n10 ) ? ( n29537 ) : ( n50070 ) ;
assign n50072 =  ( n148 ) ? ( n30575 ) : ( VREG_7_7 ) ;
assign n50073 =  ( n146 ) ? ( n30574 ) : ( n50072 ) ;
assign n50074 =  ( n144 ) ? ( n30573 ) : ( n50073 ) ;
assign n50075 =  ( n142 ) ? ( n30572 ) : ( n50074 ) ;
assign n50076 =  ( n10 ) ? ( n30571 ) : ( n50075 ) ;
assign n50077 =  ( n30582 ) ? ( VREG_7_7 ) : ( n50071 ) ;
assign n50078 =  ( n30582 ) ? ( VREG_7_7 ) : ( n50076 ) ;
assign n50079 =  ( n3034 ) ? ( n50078 ) : ( VREG_7_7 ) ;
assign n50080 =  ( n2965 ) ? ( n50077 ) : ( n50079 ) ;
assign n50081 =  ( n1930 ) ? ( n50076 ) : ( n50080 ) ;
assign n50082 =  ( n879 ) ? ( n50071 ) : ( n50081 ) ;
assign n50083 =  ( n172 ) ? ( n30593 ) : ( VREG_7_7 ) ;
assign n50084 =  ( n170 ) ? ( n30592 ) : ( n50083 ) ;
assign n50085 =  ( n168 ) ? ( n30591 ) : ( n50084 ) ;
assign n50086 =  ( n166 ) ? ( n30590 ) : ( n50085 ) ;
assign n50087 =  ( n162 ) ? ( n30589 ) : ( n50086 ) ;
assign n50088 =  ( n172 ) ? ( n30603 ) : ( VREG_7_7 ) ;
assign n50089 =  ( n170 ) ? ( n30602 ) : ( n50088 ) ;
assign n50090 =  ( n168 ) ? ( n30601 ) : ( n50089 ) ;
assign n50091 =  ( n166 ) ? ( n30600 ) : ( n50090 ) ;
assign n50092 =  ( n162 ) ? ( n30599 ) : ( n50091 ) ;
assign n50093 =  ( n30582 ) ? ( VREG_7_7 ) : ( n50092 ) ;
assign n50094 =  ( n3051 ) ? ( n50093 ) : ( VREG_7_7 ) ;
assign n50095 =  ( n3040 ) ? ( n50087 ) : ( n50094 ) ;
assign n50096 =  ( n192 ) ? ( VREG_7_7 ) : ( VREG_7_7 ) ;
assign n50097 =  ( n157 ) ? ( n50095 ) : ( n50096 ) ;
assign n50098 =  ( n6 ) ? ( n50082 ) : ( n50097 ) ;
assign n50099 =  ( n813 ) ? ( n50098 ) : ( VREG_7_7 ) ;
assign n50100 =  ( n148 ) ? ( n31660 ) : ( VREG_7_8 ) ;
assign n50101 =  ( n146 ) ? ( n31659 ) : ( n50100 ) ;
assign n50102 =  ( n144 ) ? ( n31658 ) : ( n50101 ) ;
assign n50103 =  ( n142 ) ? ( n31657 ) : ( n50102 ) ;
assign n50104 =  ( n10 ) ? ( n31656 ) : ( n50103 ) ;
assign n50105 =  ( n148 ) ? ( n32694 ) : ( VREG_7_8 ) ;
assign n50106 =  ( n146 ) ? ( n32693 ) : ( n50105 ) ;
assign n50107 =  ( n144 ) ? ( n32692 ) : ( n50106 ) ;
assign n50108 =  ( n142 ) ? ( n32691 ) : ( n50107 ) ;
assign n50109 =  ( n10 ) ? ( n32690 ) : ( n50108 ) ;
assign n50110 =  ( n32701 ) ? ( VREG_7_8 ) : ( n50104 ) ;
assign n50111 =  ( n32701 ) ? ( VREG_7_8 ) : ( n50109 ) ;
assign n50112 =  ( n3034 ) ? ( n50111 ) : ( VREG_7_8 ) ;
assign n50113 =  ( n2965 ) ? ( n50110 ) : ( n50112 ) ;
assign n50114 =  ( n1930 ) ? ( n50109 ) : ( n50113 ) ;
assign n50115 =  ( n879 ) ? ( n50104 ) : ( n50114 ) ;
assign n50116 =  ( n172 ) ? ( n32712 ) : ( VREG_7_8 ) ;
assign n50117 =  ( n170 ) ? ( n32711 ) : ( n50116 ) ;
assign n50118 =  ( n168 ) ? ( n32710 ) : ( n50117 ) ;
assign n50119 =  ( n166 ) ? ( n32709 ) : ( n50118 ) ;
assign n50120 =  ( n162 ) ? ( n32708 ) : ( n50119 ) ;
assign n50121 =  ( n172 ) ? ( n32722 ) : ( VREG_7_8 ) ;
assign n50122 =  ( n170 ) ? ( n32721 ) : ( n50121 ) ;
assign n50123 =  ( n168 ) ? ( n32720 ) : ( n50122 ) ;
assign n50124 =  ( n166 ) ? ( n32719 ) : ( n50123 ) ;
assign n50125 =  ( n162 ) ? ( n32718 ) : ( n50124 ) ;
assign n50126 =  ( n32701 ) ? ( VREG_7_8 ) : ( n50125 ) ;
assign n50127 =  ( n3051 ) ? ( n50126 ) : ( VREG_7_8 ) ;
assign n50128 =  ( n3040 ) ? ( n50120 ) : ( n50127 ) ;
assign n50129 =  ( n192 ) ? ( VREG_7_8 ) : ( VREG_7_8 ) ;
assign n50130 =  ( n157 ) ? ( n50128 ) : ( n50129 ) ;
assign n50131 =  ( n6 ) ? ( n50115 ) : ( n50130 ) ;
assign n50132 =  ( n813 ) ? ( n50131 ) : ( VREG_7_8 ) ;
assign n50133 =  ( n148 ) ? ( n33779 ) : ( VREG_7_9 ) ;
assign n50134 =  ( n146 ) ? ( n33778 ) : ( n50133 ) ;
assign n50135 =  ( n144 ) ? ( n33777 ) : ( n50134 ) ;
assign n50136 =  ( n142 ) ? ( n33776 ) : ( n50135 ) ;
assign n50137 =  ( n10 ) ? ( n33775 ) : ( n50136 ) ;
assign n50138 =  ( n148 ) ? ( n34813 ) : ( VREG_7_9 ) ;
assign n50139 =  ( n146 ) ? ( n34812 ) : ( n50138 ) ;
assign n50140 =  ( n144 ) ? ( n34811 ) : ( n50139 ) ;
assign n50141 =  ( n142 ) ? ( n34810 ) : ( n50140 ) ;
assign n50142 =  ( n10 ) ? ( n34809 ) : ( n50141 ) ;
assign n50143 =  ( n34820 ) ? ( VREG_7_9 ) : ( n50137 ) ;
assign n50144 =  ( n34820 ) ? ( VREG_7_9 ) : ( n50142 ) ;
assign n50145 =  ( n3034 ) ? ( n50144 ) : ( VREG_7_9 ) ;
assign n50146 =  ( n2965 ) ? ( n50143 ) : ( n50145 ) ;
assign n50147 =  ( n1930 ) ? ( n50142 ) : ( n50146 ) ;
assign n50148 =  ( n879 ) ? ( n50137 ) : ( n50147 ) ;
assign n50149 =  ( n172 ) ? ( n34831 ) : ( VREG_7_9 ) ;
assign n50150 =  ( n170 ) ? ( n34830 ) : ( n50149 ) ;
assign n50151 =  ( n168 ) ? ( n34829 ) : ( n50150 ) ;
assign n50152 =  ( n166 ) ? ( n34828 ) : ( n50151 ) ;
assign n50153 =  ( n162 ) ? ( n34827 ) : ( n50152 ) ;
assign n50154 =  ( n172 ) ? ( n34841 ) : ( VREG_7_9 ) ;
assign n50155 =  ( n170 ) ? ( n34840 ) : ( n50154 ) ;
assign n50156 =  ( n168 ) ? ( n34839 ) : ( n50155 ) ;
assign n50157 =  ( n166 ) ? ( n34838 ) : ( n50156 ) ;
assign n50158 =  ( n162 ) ? ( n34837 ) : ( n50157 ) ;
assign n50159 =  ( n34820 ) ? ( VREG_7_9 ) : ( n50158 ) ;
assign n50160 =  ( n3051 ) ? ( n50159 ) : ( VREG_7_9 ) ;
assign n50161 =  ( n3040 ) ? ( n50153 ) : ( n50160 ) ;
assign n50162 =  ( n192 ) ? ( VREG_7_9 ) : ( VREG_7_9 ) ;
assign n50163 =  ( n157 ) ? ( n50161 ) : ( n50162 ) ;
assign n50164 =  ( n6 ) ? ( n50148 ) : ( n50163 ) ;
assign n50165 =  ( n813 ) ? ( n50164 ) : ( VREG_7_9 ) ;
assign n50166 =  ( n148 ) ? ( n1924 ) : ( VREG_8_0 ) ;
assign n50167 =  ( n146 ) ? ( n1923 ) : ( n50166 ) ;
assign n50168 =  ( n144 ) ? ( n1922 ) : ( n50167 ) ;
assign n50169 =  ( n142 ) ? ( n1921 ) : ( n50168 ) ;
assign n50170 =  ( n10 ) ? ( n1920 ) : ( n50169 ) ;
assign n50171 =  ( n148 ) ? ( n2959 ) : ( VREG_8_0 ) ;
assign n50172 =  ( n146 ) ? ( n2958 ) : ( n50171 ) ;
assign n50173 =  ( n144 ) ? ( n2957 ) : ( n50172 ) ;
assign n50174 =  ( n142 ) ? ( n2956 ) : ( n50173 ) ;
assign n50175 =  ( n10 ) ? ( n2955 ) : ( n50174 ) ;
assign n50176 =  ( n3032 ) ? ( VREG_8_0 ) : ( n50170 ) ;
assign n50177 =  ( n3032 ) ? ( VREG_8_0 ) : ( n50175 ) ;
assign n50178 =  ( n3034 ) ? ( n50177 ) : ( VREG_8_0 ) ;
assign n50179 =  ( n2965 ) ? ( n50176 ) : ( n50178 ) ;
assign n50180 =  ( n1930 ) ? ( n50175 ) : ( n50179 ) ;
assign n50181 =  ( n879 ) ? ( n50170 ) : ( n50180 ) ;
assign n50182 =  ( n172 ) ? ( n3045 ) : ( VREG_8_0 ) ;
assign n50183 =  ( n170 ) ? ( n3044 ) : ( n50182 ) ;
assign n50184 =  ( n168 ) ? ( n3043 ) : ( n50183 ) ;
assign n50185 =  ( n166 ) ? ( n3042 ) : ( n50184 ) ;
assign n50186 =  ( n162 ) ? ( n3041 ) : ( n50185 ) ;
assign n50187 =  ( n172 ) ? ( n3056 ) : ( VREG_8_0 ) ;
assign n50188 =  ( n170 ) ? ( n3055 ) : ( n50187 ) ;
assign n50189 =  ( n168 ) ? ( n3054 ) : ( n50188 ) ;
assign n50190 =  ( n166 ) ? ( n3053 ) : ( n50189 ) ;
assign n50191 =  ( n162 ) ? ( n3052 ) : ( n50190 ) ;
assign n50192 =  ( n3032 ) ? ( VREG_8_0 ) : ( n50191 ) ;
assign n50193 =  ( n3051 ) ? ( n50192 ) : ( VREG_8_0 ) ;
assign n50194 =  ( n3040 ) ? ( n50186 ) : ( n50193 ) ;
assign n50195 =  ( n192 ) ? ( VREG_8_0 ) : ( VREG_8_0 ) ;
assign n50196 =  ( n157 ) ? ( n50194 ) : ( n50195 ) ;
assign n50197 =  ( n6 ) ? ( n50181 ) : ( n50196 ) ;
assign n50198 =  ( n835 ) ? ( n50197 ) : ( VREG_8_0 ) ;
assign n50199 =  ( n148 ) ? ( n4113 ) : ( VREG_8_1 ) ;
assign n50200 =  ( n146 ) ? ( n4112 ) : ( n50199 ) ;
assign n50201 =  ( n144 ) ? ( n4111 ) : ( n50200 ) ;
assign n50202 =  ( n142 ) ? ( n4110 ) : ( n50201 ) ;
assign n50203 =  ( n10 ) ? ( n4109 ) : ( n50202 ) ;
assign n50204 =  ( n148 ) ? ( n5147 ) : ( VREG_8_1 ) ;
assign n50205 =  ( n146 ) ? ( n5146 ) : ( n50204 ) ;
assign n50206 =  ( n144 ) ? ( n5145 ) : ( n50205 ) ;
assign n50207 =  ( n142 ) ? ( n5144 ) : ( n50206 ) ;
assign n50208 =  ( n10 ) ? ( n5143 ) : ( n50207 ) ;
assign n50209 =  ( n5154 ) ? ( VREG_8_1 ) : ( n50203 ) ;
assign n50210 =  ( n5154 ) ? ( VREG_8_1 ) : ( n50208 ) ;
assign n50211 =  ( n3034 ) ? ( n50210 ) : ( VREG_8_1 ) ;
assign n50212 =  ( n2965 ) ? ( n50209 ) : ( n50211 ) ;
assign n50213 =  ( n1930 ) ? ( n50208 ) : ( n50212 ) ;
assign n50214 =  ( n879 ) ? ( n50203 ) : ( n50213 ) ;
assign n50215 =  ( n172 ) ? ( n5165 ) : ( VREG_8_1 ) ;
assign n50216 =  ( n170 ) ? ( n5164 ) : ( n50215 ) ;
assign n50217 =  ( n168 ) ? ( n5163 ) : ( n50216 ) ;
assign n50218 =  ( n166 ) ? ( n5162 ) : ( n50217 ) ;
assign n50219 =  ( n162 ) ? ( n5161 ) : ( n50218 ) ;
assign n50220 =  ( n172 ) ? ( n5175 ) : ( VREG_8_1 ) ;
assign n50221 =  ( n170 ) ? ( n5174 ) : ( n50220 ) ;
assign n50222 =  ( n168 ) ? ( n5173 ) : ( n50221 ) ;
assign n50223 =  ( n166 ) ? ( n5172 ) : ( n50222 ) ;
assign n50224 =  ( n162 ) ? ( n5171 ) : ( n50223 ) ;
assign n50225 =  ( n5154 ) ? ( VREG_8_1 ) : ( n50224 ) ;
assign n50226 =  ( n3051 ) ? ( n50225 ) : ( VREG_8_1 ) ;
assign n50227 =  ( n3040 ) ? ( n50219 ) : ( n50226 ) ;
assign n50228 =  ( n192 ) ? ( VREG_8_1 ) : ( VREG_8_1 ) ;
assign n50229 =  ( n157 ) ? ( n50227 ) : ( n50228 ) ;
assign n50230 =  ( n6 ) ? ( n50214 ) : ( n50229 ) ;
assign n50231 =  ( n835 ) ? ( n50230 ) : ( VREG_8_1 ) ;
assign n50232 =  ( n148 ) ? ( n6232 ) : ( VREG_8_10 ) ;
assign n50233 =  ( n146 ) ? ( n6231 ) : ( n50232 ) ;
assign n50234 =  ( n144 ) ? ( n6230 ) : ( n50233 ) ;
assign n50235 =  ( n142 ) ? ( n6229 ) : ( n50234 ) ;
assign n50236 =  ( n10 ) ? ( n6228 ) : ( n50235 ) ;
assign n50237 =  ( n148 ) ? ( n7266 ) : ( VREG_8_10 ) ;
assign n50238 =  ( n146 ) ? ( n7265 ) : ( n50237 ) ;
assign n50239 =  ( n144 ) ? ( n7264 ) : ( n50238 ) ;
assign n50240 =  ( n142 ) ? ( n7263 ) : ( n50239 ) ;
assign n50241 =  ( n10 ) ? ( n7262 ) : ( n50240 ) ;
assign n50242 =  ( n7273 ) ? ( VREG_8_10 ) : ( n50236 ) ;
assign n50243 =  ( n7273 ) ? ( VREG_8_10 ) : ( n50241 ) ;
assign n50244 =  ( n3034 ) ? ( n50243 ) : ( VREG_8_10 ) ;
assign n50245 =  ( n2965 ) ? ( n50242 ) : ( n50244 ) ;
assign n50246 =  ( n1930 ) ? ( n50241 ) : ( n50245 ) ;
assign n50247 =  ( n879 ) ? ( n50236 ) : ( n50246 ) ;
assign n50248 =  ( n172 ) ? ( n7284 ) : ( VREG_8_10 ) ;
assign n50249 =  ( n170 ) ? ( n7283 ) : ( n50248 ) ;
assign n50250 =  ( n168 ) ? ( n7282 ) : ( n50249 ) ;
assign n50251 =  ( n166 ) ? ( n7281 ) : ( n50250 ) ;
assign n50252 =  ( n162 ) ? ( n7280 ) : ( n50251 ) ;
assign n50253 =  ( n172 ) ? ( n7294 ) : ( VREG_8_10 ) ;
assign n50254 =  ( n170 ) ? ( n7293 ) : ( n50253 ) ;
assign n50255 =  ( n168 ) ? ( n7292 ) : ( n50254 ) ;
assign n50256 =  ( n166 ) ? ( n7291 ) : ( n50255 ) ;
assign n50257 =  ( n162 ) ? ( n7290 ) : ( n50256 ) ;
assign n50258 =  ( n7273 ) ? ( VREG_8_10 ) : ( n50257 ) ;
assign n50259 =  ( n3051 ) ? ( n50258 ) : ( VREG_8_10 ) ;
assign n50260 =  ( n3040 ) ? ( n50252 ) : ( n50259 ) ;
assign n50261 =  ( n192 ) ? ( VREG_8_10 ) : ( VREG_8_10 ) ;
assign n50262 =  ( n157 ) ? ( n50260 ) : ( n50261 ) ;
assign n50263 =  ( n6 ) ? ( n50247 ) : ( n50262 ) ;
assign n50264 =  ( n835 ) ? ( n50263 ) : ( VREG_8_10 ) ;
assign n50265 =  ( n148 ) ? ( n8351 ) : ( VREG_8_11 ) ;
assign n50266 =  ( n146 ) ? ( n8350 ) : ( n50265 ) ;
assign n50267 =  ( n144 ) ? ( n8349 ) : ( n50266 ) ;
assign n50268 =  ( n142 ) ? ( n8348 ) : ( n50267 ) ;
assign n50269 =  ( n10 ) ? ( n8347 ) : ( n50268 ) ;
assign n50270 =  ( n148 ) ? ( n9385 ) : ( VREG_8_11 ) ;
assign n50271 =  ( n146 ) ? ( n9384 ) : ( n50270 ) ;
assign n50272 =  ( n144 ) ? ( n9383 ) : ( n50271 ) ;
assign n50273 =  ( n142 ) ? ( n9382 ) : ( n50272 ) ;
assign n50274 =  ( n10 ) ? ( n9381 ) : ( n50273 ) ;
assign n50275 =  ( n9392 ) ? ( VREG_8_11 ) : ( n50269 ) ;
assign n50276 =  ( n9392 ) ? ( VREG_8_11 ) : ( n50274 ) ;
assign n50277 =  ( n3034 ) ? ( n50276 ) : ( VREG_8_11 ) ;
assign n50278 =  ( n2965 ) ? ( n50275 ) : ( n50277 ) ;
assign n50279 =  ( n1930 ) ? ( n50274 ) : ( n50278 ) ;
assign n50280 =  ( n879 ) ? ( n50269 ) : ( n50279 ) ;
assign n50281 =  ( n172 ) ? ( n9403 ) : ( VREG_8_11 ) ;
assign n50282 =  ( n170 ) ? ( n9402 ) : ( n50281 ) ;
assign n50283 =  ( n168 ) ? ( n9401 ) : ( n50282 ) ;
assign n50284 =  ( n166 ) ? ( n9400 ) : ( n50283 ) ;
assign n50285 =  ( n162 ) ? ( n9399 ) : ( n50284 ) ;
assign n50286 =  ( n172 ) ? ( n9413 ) : ( VREG_8_11 ) ;
assign n50287 =  ( n170 ) ? ( n9412 ) : ( n50286 ) ;
assign n50288 =  ( n168 ) ? ( n9411 ) : ( n50287 ) ;
assign n50289 =  ( n166 ) ? ( n9410 ) : ( n50288 ) ;
assign n50290 =  ( n162 ) ? ( n9409 ) : ( n50289 ) ;
assign n50291 =  ( n9392 ) ? ( VREG_8_11 ) : ( n50290 ) ;
assign n50292 =  ( n3051 ) ? ( n50291 ) : ( VREG_8_11 ) ;
assign n50293 =  ( n3040 ) ? ( n50285 ) : ( n50292 ) ;
assign n50294 =  ( n192 ) ? ( VREG_8_11 ) : ( VREG_8_11 ) ;
assign n50295 =  ( n157 ) ? ( n50293 ) : ( n50294 ) ;
assign n50296 =  ( n6 ) ? ( n50280 ) : ( n50295 ) ;
assign n50297 =  ( n835 ) ? ( n50296 ) : ( VREG_8_11 ) ;
assign n50298 =  ( n148 ) ? ( n10470 ) : ( VREG_8_12 ) ;
assign n50299 =  ( n146 ) ? ( n10469 ) : ( n50298 ) ;
assign n50300 =  ( n144 ) ? ( n10468 ) : ( n50299 ) ;
assign n50301 =  ( n142 ) ? ( n10467 ) : ( n50300 ) ;
assign n50302 =  ( n10 ) ? ( n10466 ) : ( n50301 ) ;
assign n50303 =  ( n148 ) ? ( n11504 ) : ( VREG_8_12 ) ;
assign n50304 =  ( n146 ) ? ( n11503 ) : ( n50303 ) ;
assign n50305 =  ( n144 ) ? ( n11502 ) : ( n50304 ) ;
assign n50306 =  ( n142 ) ? ( n11501 ) : ( n50305 ) ;
assign n50307 =  ( n10 ) ? ( n11500 ) : ( n50306 ) ;
assign n50308 =  ( n11511 ) ? ( VREG_8_12 ) : ( n50302 ) ;
assign n50309 =  ( n11511 ) ? ( VREG_8_12 ) : ( n50307 ) ;
assign n50310 =  ( n3034 ) ? ( n50309 ) : ( VREG_8_12 ) ;
assign n50311 =  ( n2965 ) ? ( n50308 ) : ( n50310 ) ;
assign n50312 =  ( n1930 ) ? ( n50307 ) : ( n50311 ) ;
assign n50313 =  ( n879 ) ? ( n50302 ) : ( n50312 ) ;
assign n50314 =  ( n172 ) ? ( n11522 ) : ( VREG_8_12 ) ;
assign n50315 =  ( n170 ) ? ( n11521 ) : ( n50314 ) ;
assign n50316 =  ( n168 ) ? ( n11520 ) : ( n50315 ) ;
assign n50317 =  ( n166 ) ? ( n11519 ) : ( n50316 ) ;
assign n50318 =  ( n162 ) ? ( n11518 ) : ( n50317 ) ;
assign n50319 =  ( n172 ) ? ( n11532 ) : ( VREG_8_12 ) ;
assign n50320 =  ( n170 ) ? ( n11531 ) : ( n50319 ) ;
assign n50321 =  ( n168 ) ? ( n11530 ) : ( n50320 ) ;
assign n50322 =  ( n166 ) ? ( n11529 ) : ( n50321 ) ;
assign n50323 =  ( n162 ) ? ( n11528 ) : ( n50322 ) ;
assign n50324 =  ( n11511 ) ? ( VREG_8_12 ) : ( n50323 ) ;
assign n50325 =  ( n3051 ) ? ( n50324 ) : ( VREG_8_12 ) ;
assign n50326 =  ( n3040 ) ? ( n50318 ) : ( n50325 ) ;
assign n50327 =  ( n192 ) ? ( VREG_8_12 ) : ( VREG_8_12 ) ;
assign n50328 =  ( n157 ) ? ( n50326 ) : ( n50327 ) ;
assign n50329 =  ( n6 ) ? ( n50313 ) : ( n50328 ) ;
assign n50330 =  ( n835 ) ? ( n50329 ) : ( VREG_8_12 ) ;
assign n50331 =  ( n148 ) ? ( n12589 ) : ( VREG_8_13 ) ;
assign n50332 =  ( n146 ) ? ( n12588 ) : ( n50331 ) ;
assign n50333 =  ( n144 ) ? ( n12587 ) : ( n50332 ) ;
assign n50334 =  ( n142 ) ? ( n12586 ) : ( n50333 ) ;
assign n50335 =  ( n10 ) ? ( n12585 ) : ( n50334 ) ;
assign n50336 =  ( n148 ) ? ( n13623 ) : ( VREG_8_13 ) ;
assign n50337 =  ( n146 ) ? ( n13622 ) : ( n50336 ) ;
assign n50338 =  ( n144 ) ? ( n13621 ) : ( n50337 ) ;
assign n50339 =  ( n142 ) ? ( n13620 ) : ( n50338 ) ;
assign n50340 =  ( n10 ) ? ( n13619 ) : ( n50339 ) ;
assign n50341 =  ( n13630 ) ? ( VREG_8_13 ) : ( n50335 ) ;
assign n50342 =  ( n13630 ) ? ( VREG_8_13 ) : ( n50340 ) ;
assign n50343 =  ( n3034 ) ? ( n50342 ) : ( VREG_8_13 ) ;
assign n50344 =  ( n2965 ) ? ( n50341 ) : ( n50343 ) ;
assign n50345 =  ( n1930 ) ? ( n50340 ) : ( n50344 ) ;
assign n50346 =  ( n879 ) ? ( n50335 ) : ( n50345 ) ;
assign n50347 =  ( n172 ) ? ( n13641 ) : ( VREG_8_13 ) ;
assign n50348 =  ( n170 ) ? ( n13640 ) : ( n50347 ) ;
assign n50349 =  ( n168 ) ? ( n13639 ) : ( n50348 ) ;
assign n50350 =  ( n166 ) ? ( n13638 ) : ( n50349 ) ;
assign n50351 =  ( n162 ) ? ( n13637 ) : ( n50350 ) ;
assign n50352 =  ( n172 ) ? ( n13651 ) : ( VREG_8_13 ) ;
assign n50353 =  ( n170 ) ? ( n13650 ) : ( n50352 ) ;
assign n50354 =  ( n168 ) ? ( n13649 ) : ( n50353 ) ;
assign n50355 =  ( n166 ) ? ( n13648 ) : ( n50354 ) ;
assign n50356 =  ( n162 ) ? ( n13647 ) : ( n50355 ) ;
assign n50357 =  ( n13630 ) ? ( VREG_8_13 ) : ( n50356 ) ;
assign n50358 =  ( n3051 ) ? ( n50357 ) : ( VREG_8_13 ) ;
assign n50359 =  ( n3040 ) ? ( n50351 ) : ( n50358 ) ;
assign n50360 =  ( n192 ) ? ( VREG_8_13 ) : ( VREG_8_13 ) ;
assign n50361 =  ( n157 ) ? ( n50359 ) : ( n50360 ) ;
assign n50362 =  ( n6 ) ? ( n50346 ) : ( n50361 ) ;
assign n50363 =  ( n835 ) ? ( n50362 ) : ( VREG_8_13 ) ;
assign n50364 =  ( n148 ) ? ( n14708 ) : ( VREG_8_14 ) ;
assign n50365 =  ( n146 ) ? ( n14707 ) : ( n50364 ) ;
assign n50366 =  ( n144 ) ? ( n14706 ) : ( n50365 ) ;
assign n50367 =  ( n142 ) ? ( n14705 ) : ( n50366 ) ;
assign n50368 =  ( n10 ) ? ( n14704 ) : ( n50367 ) ;
assign n50369 =  ( n148 ) ? ( n15742 ) : ( VREG_8_14 ) ;
assign n50370 =  ( n146 ) ? ( n15741 ) : ( n50369 ) ;
assign n50371 =  ( n144 ) ? ( n15740 ) : ( n50370 ) ;
assign n50372 =  ( n142 ) ? ( n15739 ) : ( n50371 ) ;
assign n50373 =  ( n10 ) ? ( n15738 ) : ( n50372 ) ;
assign n50374 =  ( n15749 ) ? ( VREG_8_14 ) : ( n50368 ) ;
assign n50375 =  ( n15749 ) ? ( VREG_8_14 ) : ( n50373 ) ;
assign n50376 =  ( n3034 ) ? ( n50375 ) : ( VREG_8_14 ) ;
assign n50377 =  ( n2965 ) ? ( n50374 ) : ( n50376 ) ;
assign n50378 =  ( n1930 ) ? ( n50373 ) : ( n50377 ) ;
assign n50379 =  ( n879 ) ? ( n50368 ) : ( n50378 ) ;
assign n50380 =  ( n172 ) ? ( n15760 ) : ( VREG_8_14 ) ;
assign n50381 =  ( n170 ) ? ( n15759 ) : ( n50380 ) ;
assign n50382 =  ( n168 ) ? ( n15758 ) : ( n50381 ) ;
assign n50383 =  ( n166 ) ? ( n15757 ) : ( n50382 ) ;
assign n50384 =  ( n162 ) ? ( n15756 ) : ( n50383 ) ;
assign n50385 =  ( n172 ) ? ( n15770 ) : ( VREG_8_14 ) ;
assign n50386 =  ( n170 ) ? ( n15769 ) : ( n50385 ) ;
assign n50387 =  ( n168 ) ? ( n15768 ) : ( n50386 ) ;
assign n50388 =  ( n166 ) ? ( n15767 ) : ( n50387 ) ;
assign n50389 =  ( n162 ) ? ( n15766 ) : ( n50388 ) ;
assign n50390 =  ( n15749 ) ? ( VREG_8_14 ) : ( n50389 ) ;
assign n50391 =  ( n3051 ) ? ( n50390 ) : ( VREG_8_14 ) ;
assign n50392 =  ( n3040 ) ? ( n50384 ) : ( n50391 ) ;
assign n50393 =  ( n192 ) ? ( VREG_8_14 ) : ( VREG_8_14 ) ;
assign n50394 =  ( n157 ) ? ( n50392 ) : ( n50393 ) ;
assign n50395 =  ( n6 ) ? ( n50379 ) : ( n50394 ) ;
assign n50396 =  ( n835 ) ? ( n50395 ) : ( VREG_8_14 ) ;
assign n50397 =  ( n148 ) ? ( n16827 ) : ( VREG_8_15 ) ;
assign n50398 =  ( n146 ) ? ( n16826 ) : ( n50397 ) ;
assign n50399 =  ( n144 ) ? ( n16825 ) : ( n50398 ) ;
assign n50400 =  ( n142 ) ? ( n16824 ) : ( n50399 ) ;
assign n50401 =  ( n10 ) ? ( n16823 ) : ( n50400 ) ;
assign n50402 =  ( n148 ) ? ( n17861 ) : ( VREG_8_15 ) ;
assign n50403 =  ( n146 ) ? ( n17860 ) : ( n50402 ) ;
assign n50404 =  ( n144 ) ? ( n17859 ) : ( n50403 ) ;
assign n50405 =  ( n142 ) ? ( n17858 ) : ( n50404 ) ;
assign n50406 =  ( n10 ) ? ( n17857 ) : ( n50405 ) ;
assign n50407 =  ( n17868 ) ? ( VREG_8_15 ) : ( n50401 ) ;
assign n50408 =  ( n17868 ) ? ( VREG_8_15 ) : ( n50406 ) ;
assign n50409 =  ( n3034 ) ? ( n50408 ) : ( VREG_8_15 ) ;
assign n50410 =  ( n2965 ) ? ( n50407 ) : ( n50409 ) ;
assign n50411 =  ( n1930 ) ? ( n50406 ) : ( n50410 ) ;
assign n50412 =  ( n879 ) ? ( n50401 ) : ( n50411 ) ;
assign n50413 =  ( n172 ) ? ( n17879 ) : ( VREG_8_15 ) ;
assign n50414 =  ( n170 ) ? ( n17878 ) : ( n50413 ) ;
assign n50415 =  ( n168 ) ? ( n17877 ) : ( n50414 ) ;
assign n50416 =  ( n166 ) ? ( n17876 ) : ( n50415 ) ;
assign n50417 =  ( n162 ) ? ( n17875 ) : ( n50416 ) ;
assign n50418 =  ( n172 ) ? ( n17889 ) : ( VREG_8_15 ) ;
assign n50419 =  ( n170 ) ? ( n17888 ) : ( n50418 ) ;
assign n50420 =  ( n168 ) ? ( n17887 ) : ( n50419 ) ;
assign n50421 =  ( n166 ) ? ( n17886 ) : ( n50420 ) ;
assign n50422 =  ( n162 ) ? ( n17885 ) : ( n50421 ) ;
assign n50423 =  ( n17868 ) ? ( VREG_8_15 ) : ( n50422 ) ;
assign n50424 =  ( n3051 ) ? ( n50423 ) : ( VREG_8_15 ) ;
assign n50425 =  ( n3040 ) ? ( n50417 ) : ( n50424 ) ;
assign n50426 =  ( n192 ) ? ( VREG_8_15 ) : ( VREG_8_15 ) ;
assign n50427 =  ( n157 ) ? ( n50425 ) : ( n50426 ) ;
assign n50428 =  ( n6 ) ? ( n50412 ) : ( n50427 ) ;
assign n50429 =  ( n835 ) ? ( n50428 ) : ( VREG_8_15 ) ;
assign n50430 =  ( n148 ) ? ( n18946 ) : ( VREG_8_2 ) ;
assign n50431 =  ( n146 ) ? ( n18945 ) : ( n50430 ) ;
assign n50432 =  ( n144 ) ? ( n18944 ) : ( n50431 ) ;
assign n50433 =  ( n142 ) ? ( n18943 ) : ( n50432 ) ;
assign n50434 =  ( n10 ) ? ( n18942 ) : ( n50433 ) ;
assign n50435 =  ( n148 ) ? ( n19980 ) : ( VREG_8_2 ) ;
assign n50436 =  ( n146 ) ? ( n19979 ) : ( n50435 ) ;
assign n50437 =  ( n144 ) ? ( n19978 ) : ( n50436 ) ;
assign n50438 =  ( n142 ) ? ( n19977 ) : ( n50437 ) ;
assign n50439 =  ( n10 ) ? ( n19976 ) : ( n50438 ) ;
assign n50440 =  ( n19987 ) ? ( VREG_8_2 ) : ( n50434 ) ;
assign n50441 =  ( n19987 ) ? ( VREG_8_2 ) : ( n50439 ) ;
assign n50442 =  ( n3034 ) ? ( n50441 ) : ( VREG_8_2 ) ;
assign n50443 =  ( n2965 ) ? ( n50440 ) : ( n50442 ) ;
assign n50444 =  ( n1930 ) ? ( n50439 ) : ( n50443 ) ;
assign n50445 =  ( n879 ) ? ( n50434 ) : ( n50444 ) ;
assign n50446 =  ( n172 ) ? ( n19998 ) : ( VREG_8_2 ) ;
assign n50447 =  ( n170 ) ? ( n19997 ) : ( n50446 ) ;
assign n50448 =  ( n168 ) ? ( n19996 ) : ( n50447 ) ;
assign n50449 =  ( n166 ) ? ( n19995 ) : ( n50448 ) ;
assign n50450 =  ( n162 ) ? ( n19994 ) : ( n50449 ) ;
assign n50451 =  ( n172 ) ? ( n20008 ) : ( VREG_8_2 ) ;
assign n50452 =  ( n170 ) ? ( n20007 ) : ( n50451 ) ;
assign n50453 =  ( n168 ) ? ( n20006 ) : ( n50452 ) ;
assign n50454 =  ( n166 ) ? ( n20005 ) : ( n50453 ) ;
assign n50455 =  ( n162 ) ? ( n20004 ) : ( n50454 ) ;
assign n50456 =  ( n19987 ) ? ( VREG_8_2 ) : ( n50455 ) ;
assign n50457 =  ( n3051 ) ? ( n50456 ) : ( VREG_8_2 ) ;
assign n50458 =  ( n3040 ) ? ( n50450 ) : ( n50457 ) ;
assign n50459 =  ( n192 ) ? ( VREG_8_2 ) : ( VREG_8_2 ) ;
assign n50460 =  ( n157 ) ? ( n50458 ) : ( n50459 ) ;
assign n50461 =  ( n6 ) ? ( n50445 ) : ( n50460 ) ;
assign n50462 =  ( n835 ) ? ( n50461 ) : ( VREG_8_2 ) ;
assign n50463 =  ( n148 ) ? ( n21065 ) : ( VREG_8_3 ) ;
assign n50464 =  ( n146 ) ? ( n21064 ) : ( n50463 ) ;
assign n50465 =  ( n144 ) ? ( n21063 ) : ( n50464 ) ;
assign n50466 =  ( n142 ) ? ( n21062 ) : ( n50465 ) ;
assign n50467 =  ( n10 ) ? ( n21061 ) : ( n50466 ) ;
assign n50468 =  ( n148 ) ? ( n22099 ) : ( VREG_8_3 ) ;
assign n50469 =  ( n146 ) ? ( n22098 ) : ( n50468 ) ;
assign n50470 =  ( n144 ) ? ( n22097 ) : ( n50469 ) ;
assign n50471 =  ( n142 ) ? ( n22096 ) : ( n50470 ) ;
assign n50472 =  ( n10 ) ? ( n22095 ) : ( n50471 ) ;
assign n50473 =  ( n22106 ) ? ( VREG_8_3 ) : ( n50467 ) ;
assign n50474 =  ( n22106 ) ? ( VREG_8_3 ) : ( n50472 ) ;
assign n50475 =  ( n3034 ) ? ( n50474 ) : ( VREG_8_3 ) ;
assign n50476 =  ( n2965 ) ? ( n50473 ) : ( n50475 ) ;
assign n50477 =  ( n1930 ) ? ( n50472 ) : ( n50476 ) ;
assign n50478 =  ( n879 ) ? ( n50467 ) : ( n50477 ) ;
assign n50479 =  ( n172 ) ? ( n22117 ) : ( VREG_8_3 ) ;
assign n50480 =  ( n170 ) ? ( n22116 ) : ( n50479 ) ;
assign n50481 =  ( n168 ) ? ( n22115 ) : ( n50480 ) ;
assign n50482 =  ( n166 ) ? ( n22114 ) : ( n50481 ) ;
assign n50483 =  ( n162 ) ? ( n22113 ) : ( n50482 ) ;
assign n50484 =  ( n172 ) ? ( n22127 ) : ( VREG_8_3 ) ;
assign n50485 =  ( n170 ) ? ( n22126 ) : ( n50484 ) ;
assign n50486 =  ( n168 ) ? ( n22125 ) : ( n50485 ) ;
assign n50487 =  ( n166 ) ? ( n22124 ) : ( n50486 ) ;
assign n50488 =  ( n162 ) ? ( n22123 ) : ( n50487 ) ;
assign n50489 =  ( n22106 ) ? ( VREG_8_3 ) : ( n50488 ) ;
assign n50490 =  ( n3051 ) ? ( n50489 ) : ( VREG_8_3 ) ;
assign n50491 =  ( n3040 ) ? ( n50483 ) : ( n50490 ) ;
assign n50492 =  ( n192 ) ? ( VREG_8_3 ) : ( VREG_8_3 ) ;
assign n50493 =  ( n157 ) ? ( n50491 ) : ( n50492 ) ;
assign n50494 =  ( n6 ) ? ( n50478 ) : ( n50493 ) ;
assign n50495 =  ( n835 ) ? ( n50494 ) : ( VREG_8_3 ) ;
assign n50496 =  ( n148 ) ? ( n23184 ) : ( VREG_8_4 ) ;
assign n50497 =  ( n146 ) ? ( n23183 ) : ( n50496 ) ;
assign n50498 =  ( n144 ) ? ( n23182 ) : ( n50497 ) ;
assign n50499 =  ( n142 ) ? ( n23181 ) : ( n50498 ) ;
assign n50500 =  ( n10 ) ? ( n23180 ) : ( n50499 ) ;
assign n50501 =  ( n148 ) ? ( n24218 ) : ( VREG_8_4 ) ;
assign n50502 =  ( n146 ) ? ( n24217 ) : ( n50501 ) ;
assign n50503 =  ( n144 ) ? ( n24216 ) : ( n50502 ) ;
assign n50504 =  ( n142 ) ? ( n24215 ) : ( n50503 ) ;
assign n50505 =  ( n10 ) ? ( n24214 ) : ( n50504 ) ;
assign n50506 =  ( n24225 ) ? ( VREG_8_4 ) : ( n50500 ) ;
assign n50507 =  ( n24225 ) ? ( VREG_8_4 ) : ( n50505 ) ;
assign n50508 =  ( n3034 ) ? ( n50507 ) : ( VREG_8_4 ) ;
assign n50509 =  ( n2965 ) ? ( n50506 ) : ( n50508 ) ;
assign n50510 =  ( n1930 ) ? ( n50505 ) : ( n50509 ) ;
assign n50511 =  ( n879 ) ? ( n50500 ) : ( n50510 ) ;
assign n50512 =  ( n172 ) ? ( n24236 ) : ( VREG_8_4 ) ;
assign n50513 =  ( n170 ) ? ( n24235 ) : ( n50512 ) ;
assign n50514 =  ( n168 ) ? ( n24234 ) : ( n50513 ) ;
assign n50515 =  ( n166 ) ? ( n24233 ) : ( n50514 ) ;
assign n50516 =  ( n162 ) ? ( n24232 ) : ( n50515 ) ;
assign n50517 =  ( n172 ) ? ( n24246 ) : ( VREG_8_4 ) ;
assign n50518 =  ( n170 ) ? ( n24245 ) : ( n50517 ) ;
assign n50519 =  ( n168 ) ? ( n24244 ) : ( n50518 ) ;
assign n50520 =  ( n166 ) ? ( n24243 ) : ( n50519 ) ;
assign n50521 =  ( n162 ) ? ( n24242 ) : ( n50520 ) ;
assign n50522 =  ( n24225 ) ? ( VREG_8_4 ) : ( n50521 ) ;
assign n50523 =  ( n3051 ) ? ( n50522 ) : ( VREG_8_4 ) ;
assign n50524 =  ( n3040 ) ? ( n50516 ) : ( n50523 ) ;
assign n50525 =  ( n192 ) ? ( VREG_8_4 ) : ( VREG_8_4 ) ;
assign n50526 =  ( n157 ) ? ( n50524 ) : ( n50525 ) ;
assign n50527 =  ( n6 ) ? ( n50511 ) : ( n50526 ) ;
assign n50528 =  ( n835 ) ? ( n50527 ) : ( VREG_8_4 ) ;
assign n50529 =  ( n148 ) ? ( n25303 ) : ( VREG_8_5 ) ;
assign n50530 =  ( n146 ) ? ( n25302 ) : ( n50529 ) ;
assign n50531 =  ( n144 ) ? ( n25301 ) : ( n50530 ) ;
assign n50532 =  ( n142 ) ? ( n25300 ) : ( n50531 ) ;
assign n50533 =  ( n10 ) ? ( n25299 ) : ( n50532 ) ;
assign n50534 =  ( n148 ) ? ( n26337 ) : ( VREG_8_5 ) ;
assign n50535 =  ( n146 ) ? ( n26336 ) : ( n50534 ) ;
assign n50536 =  ( n144 ) ? ( n26335 ) : ( n50535 ) ;
assign n50537 =  ( n142 ) ? ( n26334 ) : ( n50536 ) ;
assign n50538 =  ( n10 ) ? ( n26333 ) : ( n50537 ) ;
assign n50539 =  ( n26344 ) ? ( VREG_8_5 ) : ( n50533 ) ;
assign n50540 =  ( n26344 ) ? ( VREG_8_5 ) : ( n50538 ) ;
assign n50541 =  ( n3034 ) ? ( n50540 ) : ( VREG_8_5 ) ;
assign n50542 =  ( n2965 ) ? ( n50539 ) : ( n50541 ) ;
assign n50543 =  ( n1930 ) ? ( n50538 ) : ( n50542 ) ;
assign n50544 =  ( n879 ) ? ( n50533 ) : ( n50543 ) ;
assign n50545 =  ( n172 ) ? ( n26355 ) : ( VREG_8_5 ) ;
assign n50546 =  ( n170 ) ? ( n26354 ) : ( n50545 ) ;
assign n50547 =  ( n168 ) ? ( n26353 ) : ( n50546 ) ;
assign n50548 =  ( n166 ) ? ( n26352 ) : ( n50547 ) ;
assign n50549 =  ( n162 ) ? ( n26351 ) : ( n50548 ) ;
assign n50550 =  ( n172 ) ? ( n26365 ) : ( VREG_8_5 ) ;
assign n50551 =  ( n170 ) ? ( n26364 ) : ( n50550 ) ;
assign n50552 =  ( n168 ) ? ( n26363 ) : ( n50551 ) ;
assign n50553 =  ( n166 ) ? ( n26362 ) : ( n50552 ) ;
assign n50554 =  ( n162 ) ? ( n26361 ) : ( n50553 ) ;
assign n50555 =  ( n26344 ) ? ( VREG_8_5 ) : ( n50554 ) ;
assign n50556 =  ( n3051 ) ? ( n50555 ) : ( VREG_8_5 ) ;
assign n50557 =  ( n3040 ) ? ( n50549 ) : ( n50556 ) ;
assign n50558 =  ( n192 ) ? ( VREG_8_5 ) : ( VREG_8_5 ) ;
assign n50559 =  ( n157 ) ? ( n50557 ) : ( n50558 ) ;
assign n50560 =  ( n6 ) ? ( n50544 ) : ( n50559 ) ;
assign n50561 =  ( n835 ) ? ( n50560 ) : ( VREG_8_5 ) ;
assign n50562 =  ( n148 ) ? ( n27422 ) : ( VREG_8_6 ) ;
assign n50563 =  ( n146 ) ? ( n27421 ) : ( n50562 ) ;
assign n50564 =  ( n144 ) ? ( n27420 ) : ( n50563 ) ;
assign n50565 =  ( n142 ) ? ( n27419 ) : ( n50564 ) ;
assign n50566 =  ( n10 ) ? ( n27418 ) : ( n50565 ) ;
assign n50567 =  ( n148 ) ? ( n28456 ) : ( VREG_8_6 ) ;
assign n50568 =  ( n146 ) ? ( n28455 ) : ( n50567 ) ;
assign n50569 =  ( n144 ) ? ( n28454 ) : ( n50568 ) ;
assign n50570 =  ( n142 ) ? ( n28453 ) : ( n50569 ) ;
assign n50571 =  ( n10 ) ? ( n28452 ) : ( n50570 ) ;
assign n50572 =  ( n28463 ) ? ( VREG_8_6 ) : ( n50566 ) ;
assign n50573 =  ( n28463 ) ? ( VREG_8_6 ) : ( n50571 ) ;
assign n50574 =  ( n3034 ) ? ( n50573 ) : ( VREG_8_6 ) ;
assign n50575 =  ( n2965 ) ? ( n50572 ) : ( n50574 ) ;
assign n50576 =  ( n1930 ) ? ( n50571 ) : ( n50575 ) ;
assign n50577 =  ( n879 ) ? ( n50566 ) : ( n50576 ) ;
assign n50578 =  ( n172 ) ? ( n28474 ) : ( VREG_8_6 ) ;
assign n50579 =  ( n170 ) ? ( n28473 ) : ( n50578 ) ;
assign n50580 =  ( n168 ) ? ( n28472 ) : ( n50579 ) ;
assign n50581 =  ( n166 ) ? ( n28471 ) : ( n50580 ) ;
assign n50582 =  ( n162 ) ? ( n28470 ) : ( n50581 ) ;
assign n50583 =  ( n172 ) ? ( n28484 ) : ( VREG_8_6 ) ;
assign n50584 =  ( n170 ) ? ( n28483 ) : ( n50583 ) ;
assign n50585 =  ( n168 ) ? ( n28482 ) : ( n50584 ) ;
assign n50586 =  ( n166 ) ? ( n28481 ) : ( n50585 ) ;
assign n50587 =  ( n162 ) ? ( n28480 ) : ( n50586 ) ;
assign n50588 =  ( n28463 ) ? ( VREG_8_6 ) : ( n50587 ) ;
assign n50589 =  ( n3051 ) ? ( n50588 ) : ( VREG_8_6 ) ;
assign n50590 =  ( n3040 ) ? ( n50582 ) : ( n50589 ) ;
assign n50591 =  ( n192 ) ? ( VREG_8_6 ) : ( VREG_8_6 ) ;
assign n50592 =  ( n157 ) ? ( n50590 ) : ( n50591 ) ;
assign n50593 =  ( n6 ) ? ( n50577 ) : ( n50592 ) ;
assign n50594 =  ( n835 ) ? ( n50593 ) : ( VREG_8_6 ) ;
assign n50595 =  ( n148 ) ? ( n29541 ) : ( VREG_8_7 ) ;
assign n50596 =  ( n146 ) ? ( n29540 ) : ( n50595 ) ;
assign n50597 =  ( n144 ) ? ( n29539 ) : ( n50596 ) ;
assign n50598 =  ( n142 ) ? ( n29538 ) : ( n50597 ) ;
assign n50599 =  ( n10 ) ? ( n29537 ) : ( n50598 ) ;
assign n50600 =  ( n148 ) ? ( n30575 ) : ( VREG_8_7 ) ;
assign n50601 =  ( n146 ) ? ( n30574 ) : ( n50600 ) ;
assign n50602 =  ( n144 ) ? ( n30573 ) : ( n50601 ) ;
assign n50603 =  ( n142 ) ? ( n30572 ) : ( n50602 ) ;
assign n50604 =  ( n10 ) ? ( n30571 ) : ( n50603 ) ;
assign n50605 =  ( n30582 ) ? ( VREG_8_7 ) : ( n50599 ) ;
assign n50606 =  ( n30582 ) ? ( VREG_8_7 ) : ( n50604 ) ;
assign n50607 =  ( n3034 ) ? ( n50606 ) : ( VREG_8_7 ) ;
assign n50608 =  ( n2965 ) ? ( n50605 ) : ( n50607 ) ;
assign n50609 =  ( n1930 ) ? ( n50604 ) : ( n50608 ) ;
assign n50610 =  ( n879 ) ? ( n50599 ) : ( n50609 ) ;
assign n50611 =  ( n172 ) ? ( n30593 ) : ( VREG_8_7 ) ;
assign n50612 =  ( n170 ) ? ( n30592 ) : ( n50611 ) ;
assign n50613 =  ( n168 ) ? ( n30591 ) : ( n50612 ) ;
assign n50614 =  ( n166 ) ? ( n30590 ) : ( n50613 ) ;
assign n50615 =  ( n162 ) ? ( n30589 ) : ( n50614 ) ;
assign n50616 =  ( n172 ) ? ( n30603 ) : ( VREG_8_7 ) ;
assign n50617 =  ( n170 ) ? ( n30602 ) : ( n50616 ) ;
assign n50618 =  ( n168 ) ? ( n30601 ) : ( n50617 ) ;
assign n50619 =  ( n166 ) ? ( n30600 ) : ( n50618 ) ;
assign n50620 =  ( n162 ) ? ( n30599 ) : ( n50619 ) ;
assign n50621 =  ( n30582 ) ? ( VREG_8_7 ) : ( n50620 ) ;
assign n50622 =  ( n3051 ) ? ( n50621 ) : ( VREG_8_7 ) ;
assign n50623 =  ( n3040 ) ? ( n50615 ) : ( n50622 ) ;
assign n50624 =  ( n192 ) ? ( VREG_8_7 ) : ( VREG_8_7 ) ;
assign n50625 =  ( n157 ) ? ( n50623 ) : ( n50624 ) ;
assign n50626 =  ( n6 ) ? ( n50610 ) : ( n50625 ) ;
assign n50627 =  ( n835 ) ? ( n50626 ) : ( VREG_8_7 ) ;
assign n50628 =  ( n148 ) ? ( n31660 ) : ( VREG_8_8 ) ;
assign n50629 =  ( n146 ) ? ( n31659 ) : ( n50628 ) ;
assign n50630 =  ( n144 ) ? ( n31658 ) : ( n50629 ) ;
assign n50631 =  ( n142 ) ? ( n31657 ) : ( n50630 ) ;
assign n50632 =  ( n10 ) ? ( n31656 ) : ( n50631 ) ;
assign n50633 =  ( n148 ) ? ( n32694 ) : ( VREG_8_8 ) ;
assign n50634 =  ( n146 ) ? ( n32693 ) : ( n50633 ) ;
assign n50635 =  ( n144 ) ? ( n32692 ) : ( n50634 ) ;
assign n50636 =  ( n142 ) ? ( n32691 ) : ( n50635 ) ;
assign n50637 =  ( n10 ) ? ( n32690 ) : ( n50636 ) ;
assign n50638 =  ( n32701 ) ? ( VREG_8_8 ) : ( n50632 ) ;
assign n50639 =  ( n32701 ) ? ( VREG_8_8 ) : ( n50637 ) ;
assign n50640 =  ( n3034 ) ? ( n50639 ) : ( VREG_8_8 ) ;
assign n50641 =  ( n2965 ) ? ( n50638 ) : ( n50640 ) ;
assign n50642 =  ( n1930 ) ? ( n50637 ) : ( n50641 ) ;
assign n50643 =  ( n879 ) ? ( n50632 ) : ( n50642 ) ;
assign n50644 =  ( n172 ) ? ( n32712 ) : ( VREG_8_8 ) ;
assign n50645 =  ( n170 ) ? ( n32711 ) : ( n50644 ) ;
assign n50646 =  ( n168 ) ? ( n32710 ) : ( n50645 ) ;
assign n50647 =  ( n166 ) ? ( n32709 ) : ( n50646 ) ;
assign n50648 =  ( n162 ) ? ( n32708 ) : ( n50647 ) ;
assign n50649 =  ( n172 ) ? ( n32722 ) : ( VREG_8_8 ) ;
assign n50650 =  ( n170 ) ? ( n32721 ) : ( n50649 ) ;
assign n50651 =  ( n168 ) ? ( n32720 ) : ( n50650 ) ;
assign n50652 =  ( n166 ) ? ( n32719 ) : ( n50651 ) ;
assign n50653 =  ( n162 ) ? ( n32718 ) : ( n50652 ) ;
assign n50654 =  ( n32701 ) ? ( VREG_8_8 ) : ( n50653 ) ;
assign n50655 =  ( n3051 ) ? ( n50654 ) : ( VREG_8_8 ) ;
assign n50656 =  ( n3040 ) ? ( n50648 ) : ( n50655 ) ;
assign n50657 =  ( n192 ) ? ( VREG_8_8 ) : ( VREG_8_8 ) ;
assign n50658 =  ( n157 ) ? ( n50656 ) : ( n50657 ) ;
assign n50659 =  ( n6 ) ? ( n50643 ) : ( n50658 ) ;
assign n50660 =  ( n835 ) ? ( n50659 ) : ( VREG_8_8 ) ;
assign n50661 =  ( n148 ) ? ( n33779 ) : ( VREG_8_9 ) ;
assign n50662 =  ( n146 ) ? ( n33778 ) : ( n50661 ) ;
assign n50663 =  ( n144 ) ? ( n33777 ) : ( n50662 ) ;
assign n50664 =  ( n142 ) ? ( n33776 ) : ( n50663 ) ;
assign n50665 =  ( n10 ) ? ( n33775 ) : ( n50664 ) ;
assign n50666 =  ( n148 ) ? ( n34813 ) : ( VREG_8_9 ) ;
assign n50667 =  ( n146 ) ? ( n34812 ) : ( n50666 ) ;
assign n50668 =  ( n144 ) ? ( n34811 ) : ( n50667 ) ;
assign n50669 =  ( n142 ) ? ( n34810 ) : ( n50668 ) ;
assign n50670 =  ( n10 ) ? ( n34809 ) : ( n50669 ) ;
assign n50671 =  ( n34820 ) ? ( VREG_8_9 ) : ( n50665 ) ;
assign n50672 =  ( n34820 ) ? ( VREG_8_9 ) : ( n50670 ) ;
assign n50673 =  ( n3034 ) ? ( n50672 ) : ( VREG_8_9 ) ;
assign n50674 =  ( n2965 ) ? ( n50671 ) : ( n50673 ) ;
assign n50675 =  ( n1930 ) ? ( n50670 ) : ( n50674 ) ;
assign n50676 =  ( n879 ) ? ( n50665 ) : ( n50675 ) ;
assign n50677 =  ( n172 ) ? ( n34831 ) : ( VREG_8_9 ) ;
assign n50678 =  ( n170 ) ? ( n34830 ) : ( n50677 ) ;
assign n50679 =  ( n168 ) ? ( n34829 ) : ( n50678 ) ;
assign n50680 =  ( n166 ) ? ( n34828 ) : ( n50679 ) ;
assign n50681 =  ( n162 ) ? ( n34827 ) : ( n50680 ) ;
assign n50682 =  ( n172 ) ? ( n34841 ) : ( VREG_8_9 ) ;
assign n50683 =  ( n170 ) ? ( n34840 ) : ( n50682 ) ;
assign n50684 =  ( n168 ) ? ( n34839 ) : ( n50683 ) ;
assign n50685 =  ( n166 ) ? ( n34838 ) : ( n50684 ) ;
assign n50686 =  ( n162 ) ? ( n34837 ) : ( n50685 ) ;
assign n50687 =  ( n34820 ) ? ( VREG_8_9 ) : ( n50686 ) ;
assign n50688 =  ( n3051 ) ? ( n50687 ) : ( VREG_8_9 ) ;
assign n50689 =  ( n3040 ) ? ( n50681 ) : ( n50688 ) ;
assign n50690 =  ( n192 ) ? ( VREG_8_9 ) : ( VREG_8_9 ) ;
assign n50691 =  ( n157 ) ? ( n50689 ) : ( n50690 ) ;
assign n50692 =  ( n6 ) ? ( n50676 ) : ( n50691 ) ;
assign n50693 =  ( n835 ) ? ( n50692 ) : ( VREG_8_9 ) ;
assign n50694 =  ( n148 ) ? ( n1924 ) : ( VREG_9_0 ) ;
assign n50695 =  ( n146 ) ? ( n1923 ) : ( n50694 ) ;
assign n50696 =  ( n144 ) ? ( n1922 ) : ( n50695 ) ;
assign n50697 =  ( n142 ) ? ( n1921 ) : ( n50696 ) ;
assign n50698 =  ( n10 ) ? ( n1920 ) : ( n50697 ) ;
assign n50699 =  ( n148 ) ? ( n2959 ) : ( VREG_9_0 ) ;
assign n50700 =  ( n146 ) ? ( n2958 ) : ( n50699 ) ;
assign n50701 =  ( n144 ) ? ( n2957 ) : ( n50700 ) ;
assign n50702 =  ( n142 ) ? ( n2956 ) : ( n50701 ) ;
assign n50703 =  ( n10 ) ? ( n2955 ) : ( n50702 ) ;
assign n50704 =  ( n3032 ) ? ( VREG_9_0 ) : ( n50698 ) ;
assign n50705 =  ( n3032 ) ? ( VREG_9_0 ) : ( n50703 ) ;
assign n50706 =  ( n3034 ) ? ( n50705 ) : ( VREG_9_0 ) ;
assign n50707 =  ( n2965 ) ? ( n50704 ) : ( n50706 ) ;
assign n50708 =  ( n1930 ) ? ( n50703 ) : ( n50707 ) ;
assign n50709 =  ( n879 ) ? ( n50698 ) : ( n50708 ) ;
assign n50710 =  ( n172 ) ? ( n3045 ) : ( VREG_9_0 ) ;
assign n50711 =  ( n170 ) ? ( n3044 ) : ( n50710 ) ;
assign n50712 =  ( n168 ) ? ( n3043 ) : ( n50711 ) ;
assign n50713 =  ( n166 ) ? ( n3042 ) : ( n50712 ) ;
assign n50714 =  ( n162 ) ? ( n3041 ) : ( n50713 ) ;
assign n50715 =  ( n172 ) ? ( n3056 ) : ( VREG_9_0 ) ;
assign n50716 =  ( n170 ) ? ( n3055 ) : ( n50715 ) ;
assign n50717 =  ( n168 ) ? ( n3054 ) : ( n50716 ) ;
assign n50718 =  ( n166 ) ? ( n3053 ) : ( n50717 ) ;
assign n50719 =  ( n162 ) ? ( n3052 ) : ( n50718 ) ;
assign n50720 =  ( n3032 ) ? ( VREG_9_0 ) : ( n50719 ) ;
assign n50721 =  ( n3051 ) ? ( n50720 ) : ( VREG_9_0 ) ;
assign n50722 =  ( n3040 ) ? ( n50714 ) : ( n50721 ) ;
assign n50723 =  ( n192 ) ? ( VREG_9_0 ) : ( VREG_9_0 ) ;
assign n50724 =  ( n157 ) ? ( n50722 ) : ( n50723 ) ;
assign n50725 =  ( n6 ) ? ( n50709 ) : ( n50724 ) ;
assign n50726 =  ( n857 ) ? ( n50725 ) : ( VREG_9_0 ) ;
assign n50727 =  ( n148 ) ? ( n4113 ) : ( VREG_9_1 ) ;
assign n50728 =  ( n146 ) ? ( n4112 ) : ( n50727 ) ;
assign n50729 =  ( n144 ) ? ( n4111 ) : ( n50728 ) ;
assign n50730 =  ( n142 ) ? ( n4110 ) : ( n50729 ) ;
assign n50731 =  ( n10 ) ? ( n4109 ) : ( n50730 ) ;
assign n50732 =  ( n148 ) ? ( n5147 ) : ( VREG_9_1 ) ;
assign n50733 =  ( n146 ) ? ( n5146 ) : ( n50732 ) ;
assign n50734 =  ( n144 ) ? ( n5145 ) : ( n50733 ) ;
assign n50735 =  ( n142 ) ? ( n5144 ) : ( n50734 ) ;
assign n50736 =  ( n10 ) ? ( n5143 ) : ( n50735 ) ;
assign n50737 =  ( n5154 ) ? ( VREG_9_1 ) : ( n50731 ) ;
assign n50738 =  ( n5154 ) ? ( VREG_9_1 ) : ( n50736 ) ;
assign n50739 =  ( n3034 ) ? ( n50738 ) : ( VREG_9_1 ) ;
assign n50740 =  ( n2965 ) ? ( n50737 ) : ( n50739 ) ;
assign n50741 =  ( n1930 ) ? ( n50736 ) : ( n50740 ) ;
assign n50742 =  ( n879 ) ? ( n50731 ) : ( n50741 ) ;
assign n50743 =  ( n172 ) ? ( n5165 ) : ( VREG_9_1 ) ;
assign n50744 =  ( n170 ) ? ( n5164 ) : ( n50743 ) ;
assign n50745 =  ( n168 ) ? ( n5163 ) : ( n50744 ) ;
assign n50746 =  ( n166 ) ? ( n5162 ) : ( n50745 ) ;
assign n50747 =  ( n162 ) ? ( n5161 ) : ( n50746 ) ;
assign n50748 =  ( n172 ) ? ( n5175 ) : ( VREG_9_1 ) ;
assign n50749 =  ( n170 ) ? ( n5174 ) : ( n50748 ) ;
assign n50750 =  ( n168 ) ? ( n5173 ) : ( n50749 ) ;
assign n50751 =  ( n166 ) ? ( n5172 ) : ( n50750 ) ;
assign n50752 =  ( n162 ) ? ( n5171 ) : ( n50751 ) ;
assign n50753 =  ( n5154 ) ? ( VREG_9_1 ) : ( n50752 ) ;
assign n50754 =  ( n3051 ) ? ( n50753 ) : ( VREG_9_1 ) ;
assign n50755 =  ( n3040 ) ? ( n50747 ) : ( n50754 ) ;
assign n50756 =  ( n192 ) ? ( VREG_9_1 ) : ( VREG_9_1 ) ;
assign n50757 =  ( n157 ) ? ( n50755 ) : ( n50756 ) ;
assign n50758 =  ( n6 ) ? ( n50742 ) : ( n50757 ) ;
assign n50759 =  ( n857 ) ? ( n50758 ) : ( VREG_9_1 ) ;
assign n50760 =  ( n148 ) ? ( n6232 ) : ( VREG_9_10 ) ;
assign n50761 =  ( n146 ) ? ( n6231 ) : ( n50760 ) ;
assign n50762 =  ( n144 ) ? ( n6230 ) : ( n50761 ) ;
assign n50763 =  ( n142 ) ? ( n6229 ) : ( n50762 ) ;
assign n50764 =  ( n10 ) ? ( n6228 ) : ( n50763 ) ;
assign n50765 =  ( n148 ) ? ( n7266 ) : ( VREG_9_10 ) ;
assign n50766 =  ( n146 ) ? ( n7265 ) : ( n50765 ) ;
assign n50767 =  ( n144 ) ? ( n7264 ) : ( n50766 ) ;
assign n50768 =  ( n142 ) ? ( n7263 ) : ( n50767 ) ;
assign n50769 =  ( n10 ) ? ( n7262 ) : ( n50768 ) ;
assign n50770 =  ( n7273 ) ? ( VREG_9_10 ) : ( n50764 ) ;
assign n50771 =  ( n7273 ) ? ( VREG_9_10 ) : ( n50769 ) ;
assign n50772 =  ( n3034 ) ? ( n50771 ) : ( VREG_9_10 ) ;
assign n50773 =  ( n2965 ) ? ( n50770 ) : ( n50772 ) ;
assign n50774 =  ( n1930 ) ? ( n50769 ) : ( n50773 ) ;
assign n50775 =  ( n879 ) ? ( n50764 ) : ( n50774 ) ;
assign n50776 =  ( n172 ) ? ( n7284 ) : ( VREG_9_10 ) ;
assign n50777 =  ( n170 ) ? ( n7283 ) : ( n50776 ) ;
assign n50778 =  ( n168 ) ? ( n7282 ) : ( n50777 ) ;
assign n50779 =  ( n166 ) ? ( n7281 ) : ( n50778 ) ;
assign n50780 =  ( n162 ) ? ( n7280 ) : ( n50779 ) ;
assign n50781 =  ( n172 ) ? ( n7294 ) : ( VREG_9_10 ) ;
assign n50782 =  ( n170 ) ? ( n7293 ) : ( n50781 ) ;
assign n50783 =  ( n168 ) ? ( n7292 ) : ( n50782 ) ;
assign n50784 =  ( n166 ) ? ( n7291 ) : ( n50783 ) ;
assign n50785 =  ( n162 ) ? ( n7290 ) : ( n50784 ) ;
assign n50786 =  ( n7273 ) ? ( VREG_9_10 ) : ( n50785 ) ;
assign n50787 =  ( n3051 ) ? ( n50786 ) : ( VREG_9_10 ) ;
assign n50788 =  ( n3040 ) ? ( n50780 ) : ( n50787 ) ;
assign n50789 =  ( n192 ) ? ( VREG_9_10 ) : ( VREG_9_10 ) ;
assign n50790 =  ( n157 ) ? ( n50788 ) : ( n50789 ) ;
assign n50791 =  ( n6 ) ? ( n50775 ) : ( n50790 ) ;
assign n50792 =  ( n857 ) ? ( n50791 ) : ( VREG_9_10 ) ;
assign n50793 =  ( n148 ) ? ( n8351 ) : ( VREG_9_11 ) ;
assign n50794 =  ( n146 ) ? ( n8350 ) : ( n50793 ) ;
assign n50795 =  ( n144 ) ? ( n8349 ) : ( n50794 ) ;
assign n50796 =  ( n142 ) ? ( n8348 ) : ( n50795 ) ;
assign n50797 =  ( n10 ) ? ( n8347 ) : ( n50796 ) ;
assign n50798 =  ( n148 ) ? ( n9385 ) : ( VREG_9_11 ) ;
assign n50799 =  ( n146 ) ? ( n9384 ) : ( n50798 ) ;
assign n50800 =  ( n144 ) ? ( n9383 ) : ( n50799 ) ;
assign n50801 =  ( n142 ) ? ( n9382 ) : ( n50800 ) ;
assign n50802 =  ( n10 ) ? ( n9381 ) : ( n50801 ) ;
assign n50803 =  ( n9392 ) ? ( VREG_9_11 ) : ( n50797 ) ;
assign n50804 =  ( n9392 ) ? ( VREG_9_11 ) : ( n50802 ) ;
assign n50805 =  ( n3034 ) ? ( n50804 ) : ( VREG_9_11 ) ;
assign n50806 =  ( n2965 ) ? ( n50803 ) : ( n50805 ) ;
assign n50807 =  ( n1930 ) ? ( n50802 ) : ( n50806 ) ;
assign n50808 =  ( n879 ) ? ( n50797 ) : ( n50807 ) ;
assign n50809 =  ( n172 ) ? ( n9403 ) : ( VREG_9_11 ) ;
assign n50810 =  ( n170 ) ? ( n9402 ) : ( n50809 ) ;
assign n50811 =  ( n168 ) ? ( n9401 ) : ( n50810 ) ;
assign n50812 =  ( n166 ) ? ( n9400 ) : ( n50811 ) ;
assign n50813 =  ( n162 ) ? ( n9399 ) : ( n50812 ) ;
assign n50814 =  ( n172 ) ? ( n9413 ) : ( VREG_9_11 ) ;
assign n50815 =  ( n170 ) ? ( n9412 ) : ( n50814 ) ;
assign n50816 =  ( n168 ) ? ( n9411 ) : ( n50815 ) ;
assign n50817 =  ( n166 ) ? ( n9410 ) : ( n50816 ) ;
assign n50818 =  ( n162 ) ? ( n9409 ) : ( n50817 ) ;
assign n50819 =  ( n9392 ) ? ( VREG_9_11 ) : ( n50818 ) ;
assign n50820 =  ( n3051 ) ? ( n50819 ) : ( VREG_9_11 ) ;
assign n50821 =  ( n3040 ) ? ( n50813 ) : ( n50820 ) ;
assign n50822 =  ( n192 ) ? ( VREG_9_11 ) : ( VREG_9_11 ) ;
assign n50823 =  ( n157 ) ? ( n50821 ) : ( n50822 ) ;
assign n50824 =  ( n6 ) ? ( n50808 ) : ( n50823 ) ;
assign n50825 =  ( n857 ) ? ( n50824 ) : ( VREG_9_11 ) ;
assign n50826 =  ( n148 ) ? ( n10470 ) : ( VREG_9_12 ) ;
assign n50827 =  ( n146 ) ? ( n10469 ) : ( n50826 ) ;
assign n50828 =  ( n144 ) ? ( n10468 ) : ( n50827 ) ;
assign n50829 =  ( n142 ) ? ( n10467 ) : ( n50828 ) ;
assign n50830 =  ( n10 ) ? ( n10466 ) : ( n50829 ) ;
assign n50831 =  ( n148 ) ? ( n11504 ) : ( VREG_9_12 ) ;
assign n50832 =  ( n146 ) ? ( n11503 ) : ( n50831 ) ;
assign n50833 =  ( n144 ) ? ( n11502 ) : ( n50832 ) ;
assign n50834 =  ( n142 ) ? ( n11501 ) : ( n50833 ) ;
assign n50835 =  ( n10 ) ? ( n11500 ) : ( n50834 ) ;
assign n50836 =  ( n11511 ) ? ( VREG_9_12 ) : ( n50830 ) ;
assign n50837 =  ( n11511 ) ? ( VREG_9_12 ) : ( n50835 ) ;
assign n50838 =  ( n3034 ) ? ( n50837 ) : ( VREG_9_12 ) ;
assign n50839 =  ( n2965 ) ? ( n50836 ) : ( n50838 ) ;
assign n50840 =  ( n1930 ) ? ( n50835 ) : ( n50839 ) ;
assign n50841 =  ( n879 ) ? ( n50830 ) : ( n50840 ) ;
assign n50842 =  ( n172 ) ? ( n11522 ) : ( VREG_9_12 ) ;
assign n50843 =  ( n170 ) ? ( n11521 ) : ( n50842 ) ;
assign n50844 =  ( n168 ) ? ( n11520 ) : ( n50843 ) ;
assign n50845 =  ( n166 ) ? ( n11519 ) : ( n50844 ) ;
assign n50846 =  ( n162 ) ? ( n11518 ) : ( n50845 ) ;
assign n50847 =  ( n172 ) ? ( n11532 ) : ( VREG_9_12 ) ;
assign n50848 =  ( n170 ) ? ( n11531 ) : ( n50847 ) ;
assign n50849 =  ( n168 ) ? ( n11530 ) : ( n50848 ) ;
assign n50850 =  ( n166 ) ? ( n11529 ) : ( n50849 ) ;
assign n50851 =  ( n162 ) ? ( n11528 ) : ( n50850 ) ;
assign n50852 =  ( n11511 ) ? ( VREG_9_12 ) : ( n50851 ) ;
assign n50853 =  ( n3051 ) ? ( n50852 ) : ( VREG_9_12 ) ;
assign n50854 =  ( n3040 ) ? ( n50846 ) : ( n50853 ) ;
assign n50855 =  ( n192 ) ? ( VREG_9_12 ) : ( VREG_9_12 ) ;
assign n50856 =  ( n157 ) ? ( n50854 ) : ( n50855 ) ;
assign n50857 =  ( n6 ) ? ( n50841 ) : ( n50856 ) ;
assign n50858 =  ( n857 ) ? ( n50857 ) : ( VREG_9_12 ) ;
assign n50859 =  ( n148 ) ? ( n12589 ) : ( VREG_9_13 ) ;
assign n50860 =  ( n146 ) ? ( n12588 ) : ( n50859 ) ;
assign n50861 =  ( n144 ) ? ( n12587 ) : ( n50860 ) ;
assign n50862 =  ( n142 ) ? ( n12586 ) : ( n50861 ) ;
assign n50863 =  ( n10 ) ? ( n12585 ) : ( n50862 ) ;
assign n50864 =  ( n148 ) ? ( n13623 ) : ( VREG_9_13 ) ;
assign n50865 =  ( n146 ) ? ( n13622 ) : ( n50864 ) ;
assign n50866 =  ( n144 ) ? ( n13621 ) : ( n50865 ) ;
assign n50867 =  ( n142 ) ? ( n13620 ) : ( n50866 ) ;
assign n50868 =  ( n10 ) ? ( n13619 ) : ( n50867 ) ;
assign n50869 =  ( n13630 ) ? ( VREG_9_13 ) : ( n50863 ) ;
assign n50870 =  ( n13630 ) ? ( VREG_9_13 ) : ( n50868 ) ;
assign n50871 =  ( n3034 ) ? ( n50870 ) : ( VREG_9_13 ) ;
assign n50872 =  ( n2965 ) ? ( n50869 ) : ( n50871 ) ;
assign n50873 =  ( n1930 ) ? ( n50868 ) : ( n50872 ) ;
assign n50874 =  ( n879 ) ? ( n50863 ) : ( n50873 ) ;
assign n50875 =  ( n172 ) ? ( n13641 ) : ( VREG_9_13 ) ;
assign n50876 =  ( n170 ) ? ( n13640 ) : ( n50875 ) ;
assign n50877 =  ( n168 ) ? ( n13639 ) : ( n50876 ) ;
assign n50878 =  ( n166 ) ? ( n13638 ) : ( n50877 ) ;
assign n50879 =  ( n162 ) ? ( n13637 ) : ( n50878 ) ;
assign n50880 =  ( n172 ) ? ( n13651 ) : ( VREG_9_13 ) ;
assign n50881 =  ( n170 ) ? ( n13650 ) : ( n50880 ) ;
assign n50882 =  ( n168 ) ? ( n13649 ) : ( n50881 ) ;
assign n50883 =  ( n166 ) ? ( n13648 ) : ( n50882 ) ;
assign n50884 =  ( n162 ) ? ( n13647 ) : ( n50883 ) ;
assign n50885 =  ( n13630 ) ? ( VREG_9_13 ) : ( n50884 ) ;
assign n50886 =  ( n3051 ) ? ( n50885 ) : ( VREG_9_13 ) ;
assign n50887 =  ( n3040 ) ? ( n50879 ) : ( n50886 ) ;
assign n50888 =  ( n192 ) ? ( VREG_9_13 ) : ( VREG_9_13 ) ;
assign n50889 =  ( n157 ) ? ( n50887 ) : ( n50888 ) ;
assign n50890 =  ( n6 ) ? ( n50874 ) : ( n50889 ) ;
assign n50891 =  ( n857 ) ? ( n50890 ) : ( VREG_9_13 ) ;
assign n50892 =  ( n148 ) ? ( n14708 ) : ( VREG_9_14 ) ;
assign n50893 =  ( n146 ) ? ( n14707 ) : ( n50892 ) ;
assign n50894 =  ( n144 ) ? ( n14706 ) : ( n50893 ) ;
assign n50895 =  ( n142 ) ? ( n14705 ) : ( n50894 ) ;
assign n50896 =  ( n10 ) ? ( n14704 ) : ( n50895 ) ;
assign n50897 =  ( n148 ) ? ( n15742 ) : ( VREG_9_14 ) ;
assign n50898 =  ( n146 ) ? ( n15741 ) : ( n50897 ) ;
assign n50899 =  ( n144 ) ? ( n15740 ) : ( n50898 ) ;
assign n50900 =  ( n142 ) ? ( n15739 ) : ( n50899 ) ;
assign n50901 =  ( n10 ) ? ( n15738 ) : ( n50900 ) ;
assign n50902 =  ( n15749 ) ? ( VREG_9_14 ) : ( n50896 ) ;
assign n50903 =  ( n15749 ) ? ( VREG_9_14 ) : ( n50901 ) ;
assign n50904 =  ( n3034 ) ? ( n50903 ) : ( VREG_9_14 ) ;
assign n50905 =  ( n2965 ) ? ( n50902 ) : ( n50904 ) ;
assign n50906 =  ( n1930 ) ? ( n50901 ) : ( n50905 ) ;
assign n50907 =  ( n879 ) ? ( n50896 ) : ( n50906 ) ;
assign n50908 =  ( n172 ) ? ( n15760 ) : ( VREG_9_14 ) ;
assign n50909 =  ( n170 ) ? ( n15759 ) : ( n50908 ) ;
assign n50910 =  ( n168 ) ? ( n15758 ) : ( n50909 ) ;
assign n50911 =  ( n166 ) ? ( n15757 ) : ( n50910 ) ;
assign n50912 =  ( n162 ) ? ( n15756 ) : ( n50911 ) ;
assign n50913 =  ( n172 ) ? ( n15770 ) : ( VREG_9_14 ) ;
assign n50914 =  ( n170 ) ? ( n15769 ) : ( n50913 ) ;
assign n50915 =  ( n168 ) ? ( n15768 ) : ( n50914 ) ;
assign n50916 =  ( n166 ) ? ( n15767 ) : ( n50915 ) ;
assign n50917 =  ( n162 ) ? ( n15766 ) : ( n50916 ) ;
assign n50918 =  ( n15749 ) ? ( VREG_9_14 ) : ( n50917 ) ;
assign n50919 =  ( n3051 ) ? ( n50918 ) : ( VREG_9_14 ) ;
assign n50920 =  ( n3040 ) ? ( n50912 ) : ( n50919 ) ;
assign n50921 =  ( n192 ) ? ( VREG_9_14 ) : ( VREG_9_14 ) ;
assign n50922 =  ( n157 ) ? ( n50920 ) : ( n50921 ) ;
assign n50923 =  ( n6 ) ? ( n50907 ) : ( n50922 ) ;
assign n50924 =  ( n857 ) ? ( n50923 ) : ( VREG_9_14 ) ;
assign n50925 =  ( n148 ) ? ( n16827 ) : ( VREG_9_15 ) ;
assign n50926 =  ( n146 ) ? ( n16826 ) : ( n50925 ) ;
assign n50927 =  ( n144 ) ? ( n16825 ) : ( n50926 ) ;
assign n50928 =  ( n142 ) ? ( n16824 ) : ( n50927 ) ;
assign n50929 =  ( n10 ) ? ( n16823 ) : ( n50928 ) ;
assign n50930 =  ( n148 ) ? ( n17861 ) : ( VREG_9_15 ) ;
assign n50931 =  ( n146 ) ? ( n17860 ) : ( n50930 ) ;
assign n50932 =  ( n144 ) ? ( n17859 ) : ( n50931 ) ;
assign n50933 =  ( n142 ) ? ( n17858 ) : ( n50932 ) ;
assign n50934 =  ( n10 ) ? ( n17857 ) : ( n50933 ) ;
assign n50935 =  ( n17868 ) ? ( VREG_9_15 ) : ( n50929 ) ;
assign n50936 =  ( n17868 ) ? ( VREG_9_15 ) : ( n50934 ) ;
assign n50937 =  ( n3034 ) ? ( n50936 ) : ( VREG_9_15 ) ;
assign n50938 =  ( n2965 ) ? ( n50935 ) : ( n50937 ) ;
assign n50939 =  ( n1930 ) ? ( n50934 ) : ( n50938 ) ;
assign n50940 =  ( n879 ) ? ( n50929 ) : ( n50939 ) ;
assign n50941 =  ( n172 ) ? ( n17879 ) : ( VREG_9_15 ) ;
assign n50942 =  ( n170 ) ? ( n17878 ) : ( n50941 ) ;
assign n50943 =  ( n168 ) ? ( n17877 ) : ( n50942 ) ;
assign n50944 =  ( n166 ) ? ( n17876 ) : ( n50943 ) ;
assign n50945 =  ( n162 ) ? ( n17875 ) : ( n50944 ) ;
assign n50946 =  ( n172 ) ? ( n17889 ) : ( VREG_9_15 ) ;
assign n50947 =  ( n170 ) ? ( n17888 ) : ( n50946 ) ;
assign n50948 =  ( n168 ) ? ( n17887 ) : ( n50947 ) ;
assign n50949 =  ( n166 ) ? ( n17886 ) : ( n50948 ) ;
assign n50950 =  ( n162 ) ? ( n17885 ) : ( n50949 ) ;
assign n50951 =  ( n17868 ) ? ( VREG_9_15 ) : ( n50950 ) ;
assign n50952 =  ( n3051 ) ? ( n50951 ) : ( VREG_9_15 ) ;
assign n50953 =  ( n3040 ) ? ( n50945 ) : ( n50952 ) ;
assign n50954 =  ( n192 ) ? ( VREG_9_15 ) : ( VREG_9_15 ) ;
assign n50955 =  ( n157 ) ? ( n50953 ) : ( n50954 ) ;
assign n50956 =  ( n6 ) ? ( n50940 ) : ( n50955 ) ;
assign n50957 =  ( n857 ) ? ( n50956 ) : ( VREG_9_15 ) ;
assign n50958 =  ( n148 ) ? ( n18946 ) : ( VREG_9_2 ) ;
assign n50959 =  ( n146 ) ? ( n18945 ) : ( n50958 ) ;
assign n50960 =  ( n144 ) ? ( n18944 ) : ( n50959 ) ;
assign n50961 =  ( n142 ) ? ( n18943 ) : ( n50960 ) ;
assign n50962 =  ( n10 ) ? ( n18942 ) : ( n50961 ) ;
assign n50963 =  ( n148 ) ? ( n19980 ) : ( VREG_9_2 ) ;
assign n50964 =  ( n146 ) ? ( n19979 ) : ( n50963 ) ;
assign n50965 =  ( n144 ) ? ( n19978 ) : ( n50964 ) ;
assign n50966 =  ( n142 ) ? ( n19977 ) : ( n50965 ) ;
assign n50967 =  ( n10 ) ? ( n19976 ) : ( n50966 ) ;
assign n50968 =  ( n19987 ) ? ( VREG_9_2 ) : ( n50962 ) ;
assign n50969 =  ( n19987 ) ? ( VREG_9_2 ) : ( n50967 ) ;
assign n50970 =  ( n3034 ) ? ( n50969 ) : ( VREG_9_2 ) ;
assign n50971 =  ( n2965 ) ? ( n50968 ) : ( n50970 ) ;
assign n50972 =  ( n1930 ) ? ( n50967 ) : ( n50971 ) ;
assign n50973 =  ( n879 ) ? ( n50962 ) : ( n50972 ) ;
assign n50974 =  ( n172 ) ? ( n19998 ) : ( VREG_9_2 ) ;
assign n50975 =  ( n170 ) ? ( n19997 ) : ( n50974 ) ;
assign n50976 =  ( n168 ) ? ( n19996 ) : ( n50975 ) ;
assign n50977 =  ( n166 ) ? ( n19995 ) : ( n50976 ) ;
assign n50978 =  ( n162 ) ? ( n19994 ) : ( n50977 ) ;
assign n50979 =  ( n172 ) ? ( n20008 ) : ( VREG_9_2 ) ;
assign n50980 =  ( n170 ) ? ( n20007 ) : ( n50979 ) ;
assign n50981 =  ( n168 ) ? ( n20006 ) : ( n50980 ) ;
assign n50982 =  ( n166 ) ? ( n20005 ) : ( n50981 ) ;
assign n50983 =  ( n162 ) ? ( n20004 ) : ( n50982 ) ;
assign n50984 =  ( n19987 ) ? ( VREG_9_2 ) : ( n50983 ) ;
assign n50985 =  ( n3051 ) ? ( n50984 ) : ( VREG_9_2 ) ;
assign n50986 =  ( n3040 ) ? ( n50978 ) : ( n50985 ) ;
assign n50987 =  ( n192 ) ? ( VREG_9_2 ) : ( VREG_9_2 ) ;
assign n50988 =  ( n157 ) ? ( n50986 ) : ( n50987 ) ;
assign n50989 =  ( n6 ) ? ( n50973 ) : ( n50988 ) ;
assign n50990 =  ( n857 ) ? ( n50989 ) : ( VREG_9_2 ) ;
assign n50991 =  ( n148 ) ? ( n21065 ) : ( VREG_9_3 ) ;
assign n50992 =  ( n146 ) ? ( n21064 ) : ( n50991 ) ;
assign n50993 =  ( n144 ) ? ( n21063 ) : ( n50992 ) ;
assign n50994 =  ( n142 ) ? ( n21062 ) : ( n50993 ) ;
assign n50995 =  ( n10 ) ? ( n21061 ) : ( n50994 ) ;
assign n50996 =  ( n148 ) ? ( n22099 ) : ( VREG_9_3 ) ;
assign n50997 =  ( n146 ) ? ( n22098 ) : ( n50996 ) ;
assign n50998 =  ( n144 ) ? ( n22097 ) : ( n50997 ) ;
assign n50999 =  ( n142 ) ? ( n22096 ) : ( n50998 ) ;
assign n51000 =  ( n10 ) ? ( n22095 ) : ( n50999 ) ;
assign n51001 =  ( n22106 ) ? ( VREG_9_3 ) : ( n50995 ) ;
assign n51002 =  ( n22106 ) ? ( VREG_9_3 ) : ( n51000 ) ;
assign n51003 =  ( n3034 ) ? ( n51002 ) : ( VREG_9_3 ) ;
assign n51004 =  ( n2965 ) ? ( n51001 ) : ( n51003 ) ;
assign n51005 =  ( n1930 ) ? ( n51000 ) : ( n51004 ) ;
assign n51006 =  ( n879 ) ? ( n50995 ) : ( n51005 ) ;
assign n51007 =  ( n172 ) ? ( n22117 ) : ( VREG_9_3 ) ;
assign n51008 =  ( n170 ) ? ( n22116 ) : ( n51007 ) ;
assign n51009 =  ( n168 ) ? ( n22115 ) : ( n51008 ) ;
assign n51010 =  ( n166 ) ? ( n22114 ) : ( n51009 ) ;
assign n51011 =  ( n162 ) ? ( n22113 ) : ( n51010 ) ;
assign n51012 =  ( n172 ) ? ( n22127 ) : ( VREG_9_3 ) ;
assign n51013 =  ( n170 ) ? ( n22126 ) : ( n51012 ) ;
assign n51014 =  ( n168 ) ? ( n22125 ) : ( n51013 ) ;
assign n51015 =  ( n166 ) ? ( n22124 ) : ( n51014 ) ;
assign n51016 =  ( n162 ) ? ( n22123 ) : ( n51015 ) ;
assign n51017 =  ( n22106 ) ? ( VREG_9_3 ) : ( n51016 ) ;
assign n51018 =  ( n3051 ) ? ( n51017 ) : ( VREG_9_3 ) ;
assign n51019 =  ( n3040 ) ? ( n51011 ) : ( n51018 ) ;
assign n51020 =  ( n192 ) ? ( VREG_9_3 ) : ( VREG_9_3 ) ;
assign n51021 =  ( n157 ) ? ( n51019 ) : ( n51020 ) ;
assign n51022 =  ( n6 ) ? ( n51006 ) : ( n51021 ) ;
assign n51023 =  ( n857 ) ? ( n51022 ) : ( VREG_9_3 ) ;
assign n51024 =  ( n148 ) ? ( n23184 ) : ( VREG_9_4 ) ;
assign n51025 =  ( n146 ) ? ( n23183 ) : ( n51024 ) ;
assign n51026 =  ( n144 ) ? ( n23182 ) : ( n51025 ) ;
assign n51027 =  ( n142 ) ? ( n23181 ) : ( n51026 ) ;
assign n51028 =  ( n10 ) ? ( n23180 ) : ( n51027 ) ;
assign n51029 =  ( n148 ) ? ( n24218 ) : ( VREG_9_4 ) ;
assign n51030 =  ( n146 ) ? ( n24217 ) : ( n51029 ) ;
assign n51031 =  ( n144 ) ? ( n24216 ) : ( n51030 ) ;
assign n51032 =  ( n142 ) ? ( n24215 ) : ( n51031 ) ;
assign n51033 =  ( n10 ) ? ( n24214 ) : ( n51032 ) ;
assign n51034 =  ( n24225 ) ? ( VREG_9_4 ) : ( n51028 ) ;
assign n51035 =  ( n24225 ) ? ( VREG_9_4 ) : ( n51033 ) ;
assign n51036 =  ( n3034 ) ? ( n51035 ) : ( VREG_9_4 ) ;
assign n51037 =  ( n2965 ) ? ( n51034 ) : ( n51036 ) ;
assign n51038 =  ( n1930 ) ? ( n51033 ) : ( n51037 ) ;
assign n51039 =  ( n879 ) ? ( n51028 ) : ( n51038 ) ;
assign n51040 =  ( n172 ) ? ( n24236 ) : ( VREG_9_4 ) ;
assign n51041 =  ( n170 ) ? ( n24235 ) : ( n51040 ) ;
assign n51042 =  ( n168 ) ? ( n24234 ) : ( n51041 ) ;
assign n51043 =  ( n166 ) ? ( n24233 ) : ( n51042 ) ;
assign n51044 =  ( n162 ) ? ( n24232 ) : ( n51043 ) ;
assign n51045 =  ( n172 ) ? ( n24246 ) : ( VREG_9_4 ) ;
assign n51046 =  ( n170 ) ? ( n24245 ) : ( n51045 ) ;
assign n51047 =  ( n168 ) ? ( n24244 ) : ( n51046 ) ;
assign n51048 =  ( n166 ) ? ( n24243 ) : ( n51047 ) ;
assign n51049 =  ( n162 ) ? ( n24242 ) : ( n51048 ) ;
assign n51050 =  ( n24225 ) ? ( VREG_9_4 ) : ( n51049 ) ;
assign n51051 =  ( n3051 ) ? ( n51050 ) : ( VREG_9_4 ) ;
assign n51052 =  ( n3040 ) ? ( n51044 ) : ( n51051 ) ;
assign n51053 =  ( n192 ) ? ( VREG_9_4 ) : ( VREG_9_4 ) ;
assign n51054 =  ( n157 ) ? ( n51052 ) : ( n51053 ) ;
assign n51055 =  ( n6 ) ? ( n51039 ) : ( n51054 ) ;
assign n51056 =  ( n857 ) ? ( n51055 ) : ( VREG_9_4 ) ;
assign n51057 =  ( n148 ) ? ( n25303 ) : ( VREG_9_5 ) ;
assign n51058 =  ( n146 ) ? ( n25302 ) : ( n51057 ) ;
assign n51059 =  ( n144 ) ? ( n25301 ) : ( n51058 ) ;
assign n51060 =  ( n142 ) ? ( n25300 ) : ( n51059 ) ;
assign n51061 =  ( n10 ) ? ( n25299 ) : ( n51060 ) ;
assign n51062 =  ( n148 ) ? ( n26337 ) : ( VREG_9_5 ) ;
assign n51063 =  ( n146 ) ? ( n26336 ) : ( n51062 ) ;
assign n51064 =  ( n144 ) ? ( n26335 ) : ( n51063 ) ;
assign n51065 =  ( n142 ) ? ( n26334 ) : ( n51064 ) ;
assign n51066 =  ( n10 ) ? ( n26333 ) : ( n51065 ) ;
assign n51067 =  ( n26344 ) ? ( VREG_9_5 ) : ( n51061 ) ;
assign n51068 =  ( n26344 ) ? ( VREG_9_5 ) : ( n51066 ) ;
assign n51069 =  ( n3034 ) ? ( n51068 ) : ( VREG_9_5 ) ;
assign n51070 =  ( n2965 ) ? ( n51067 ) : ( n51069 ) ;
assign n51071 =  ( n1930 ) ? ( n51066 ) : ( n51070 ) ;
assign n51072 =  ( n879 ) ? ( n51061 ) : ( n51071 ) ;
assign n51073 =  ( n172 ) ? ( n26355 ) : ( VREG_9_5 ) ;
assign n51074 =  ( n170 ) ? ( n26354 ) : ( n51073 ) ;
assign n51075 =  ( n168 ) ? ( n26353 ) : ( n51074 ) ;
assign n51076 =  ( n166 ) ? ( n26352 ) : ( n51075 ) ;
assign n51077 =  ( n162 ) ? ( n26351 ) : ( n51076 ) ;
assign n51078 =  ( n172 ) ? ( n26365 ) : ( VREG_9_5 ) ;
assign n51079 =  ( n170 ) ? ( n26364 ) : ( n51078 ) ;
assign n51080 =  ( n168 ) ? ( n26363 ) : ( n51079 ) ;
assign n51081 =  ( n166 ) ? ( n26362 ) : ( n51080 ) ;
assign n51082 =  ( n162 ) ? ( n26361 ) : ( n51081 ) ;
assign n51083 =  ( n26344 ) ? ( VREG_9_5 ) : ( n51082 ) ;
assign n51084 =  ( n3051 ) ? ( n51083 ) : ( VREG_9_5 ) ;
assign n51085 =  ( n3040 ) ? ( n51077 ) : ( n51084 ) ;
assign n51086 =  ( n192 ) ? ( VREG_9_5 ) : ( VREG_9_5 ) ;
assign n51087 =  ( n157 ) ? ( n51085 ) : ( n51086 ) ;
assign n51088 =  ( n6 ) ? ( n51072 ) : ( n51087 ) ;
assign n51089 =  ( n857 ) ? ( n51088 ) : ( VREG_9_5 ) ;
assign n51090 =  ( n148 ) ? ( n27422 ) : ( VREG_9_6 ) ;
assign n51091 =  ( n146 ) ? ( n27421 ) : ( n51090 ) ;
assign n51092 =  ( n144 ) ? ( n27420 ) : ( n51091 ) ;
assign n51093 =  ( n142 ) ? ( n27419 ) : ( n51092 ) ;
assign n51094 =  ( n10 ) ? ( n27418 ) : ( n51093 ) ;
assign n51095 =  ( n148 ) ? ( n28456 ) : ( VREG_9_6 ) ;
assign n51096 =  ( n146 ) ? ( n28455 ) : ( n51095 ) ;
assign n51097 =  ( n144 ) ? ( n28454 ) : ( n51096 ) ;
assign n51098 =  ( n142 ) ? ( n28453 ) : ( n51097 ) ;
assign n51099 =  ( n10 ) ? ( n28452 ) : ( n51098 ) ;
assign n51100 =  ( n28463 ) ? ( VREG_9_6 ) : ( n51094 ) ;
assign n51101 =  ( n28463 ) ? ( VREG_9_6 ) : ( n51099 ) ;
assign n51102 =  ( n3034 ) ? ( n51101 ) : ( VREG_9_6 ) ;
assign n51103 =  ( n2965 ) ? ( n51100 ) : ( n51102 ) ;
assign n51104 =  ( n1930 ) ? ( n51099 ) : ( n51103 ) ;
assign n51105 =  ( n879 ) ? ( n51094 ) : ( n51104 ) ;
assign n51106 =  ( n172 ) ? ( n28474 ) : ( VREG_9_6 ) ;
assign n51107 =  ( n170 ) ? ( n28473 ) : ( n51106 ) ;
assign n51108 =  ( n168 ) ? ( n28472 ) : ( n51107 ) ;
assign n51109 =  ( n166 ) ? ( n28471 ) : ( n51108 ) ;
assign n51110 =  ( n162 ) ? ( n28470 ) : ( n51109 ) ;
assign n51111 =  ( n172 ) ? ( n28484 ) : ( VREG_9_6 ) ;
assign n51112 =  ( n170 ) ? ( n28483 ) : ( n51111 ) ;
assign n51113 =  ( n168 ) ? ( n28482 ) : ( n51112 ) ;
assign n51114 =  ( n166 ) ? ( n28481 ) : ( n51113 ) ;
assign n51115 =  ( n162 ) ? ( n28480 ) : ( n51114 ) ;
assign n51116 =  ( n28463 ) ? ( VREG_9_6 ) : ( n51115 ) ;
assign n51117 =  ( n3051 ) ? ( n51116 ) : ( VREG_9_6 ) ;
assign n51118 =  ( n3040 ) ? ( n51110 ) : ( n51117 ) ;
assign n51119 =  ( n192 ) ? ( VREG_9_6 ) : ( VREG_9_6 ) ;
assign n51120 =  ( n157 ) ? ( n51118 ) : ( n51119 ) ;
assign n51121 =  ( n6 ) ? ( n51105 ) : ( n51120 ) ;
assign n51122 =  ( n857 ) ? ( n51121 ) : ( VREG_9_6 ) ;
assign n51123 =  ( n148 ) ? ( n29541 ) : ( VREG_9_7 ) ;
assign n51124 =  ( n146 ) ? ( n29540 ) : ( n51123 ) ;
assign n51125 =  ( n144 ) ? ( n29539 ) : ( n51124 ) ;
assign n51126 =  ( n142 ) ? ( n29538 ) : ( n51125 ) ;
assign n51127 =  ( n10 ) ? ( n29537 ) : ( n51126 ) ;
assign n51128 =  ( n148 ) ? ( n30575 ) : ( VREG_9_7 ) ;
assign n51129 =  ( n146 ) ? ( n30574 ) : ( n51128 ) ;
assign n51130 =  ( n144 ) ? ( n30573 ) : ( n51129 ) ;
assign n51131 =  ( n142 ) ? ( n30572 ) : ( n51130 ) ;
assign n51132 =  ( n10 ) ? ( n30571 ) : ( n51131 ) ;
assign n51133 =  ( n30582 ) ? ( VREG_9_7 ) : ( n51127 ) ;
assign n51134 =  ( n30582 ) ? ( VREG_9_7 ) : ( n51132 ) ;
assign n51135 =  ( n3034 ) ? ( n51134 ) : ( VREG_9_7 ) ;
assign n51136 =  ( n2965 ) ? ( n51133 ) : ( n51135 ) ;
assign n51137 =  ( n1930 ) ? ( n51132 ) : ( n51136 ) ;
assign n51138 =  ( n879 ) ? ( n51127 ) : ( n51137 ) ;
assign n51139 =  ( n172 ) ? ( n30593 ) : ( VREG_9_7 ) ;
assign n51140 =  ( n170 ) ? ( n30592 ) : ( n51139 ) ;
assign n51141 =  ( n168 ) ? ( n30591 ) : ( n51140 ) ;
assign n51142 =  ( n166 ) ? ( n30590 ) : ( n51141 ) ;
assign n51143 =  ( n162 ) ? ( n30589 ) : ( n51142 ) ;
assign n51144 =  ( n172 ) ? ( n30603 ) : ( VREG_9_7 ) ;
assign n51145 =  ( n170 ) ? ( n30602 ) : ( n51144 ) ;
assign n51146 =  ( n168 ) ? ( n30601 ) : ( n51145 ) ;
assign n51147 =  ( n166 ) ? ( n30600 ) : ( n51146 ) ;
assign n51148 =  ( n162 ) ? ( n30599 ) : ( n51147 ) ;
assign n51149 =  ( n30582 ) ? ( VREG_9_7 ) : ( n51148 ) ;
assign n51150 =  ( n3051 ) ? ( n51149 ) : ( VREG_9_7 ) ;
assign n51151 =  ( n3040 ) ? ( n51143 ) : ( n51150 ) ;
assign n51152 =  ( n192 ) ? ( VREG_9_7 ) : ( VREG_9_7 ) ;
assign n51153 =  ( n157 ) ? ( n51151 ) : ( n51152 ) ;
assign n51154 =  ( n6 ) ? ( n51138 ) : ( n51153 ) ;
assign n51155 =  ( n857 ) ? ( n51154 ) : ( VREG_9_7 ) ;
assign n51156 =  ( n148 ) ? ( n31660 ) : ( VREG_9_8 ) ;
assign n51157 =  ( n146 ) ? ( n31659 ) : ( n51156 ) ;
assign n51158 =  ( n144 ) ? ( n31658 ) : ( n51157 ) ;
assign n51159 =  ( n142 ) ? ( n31657 ) : ( n51158 ) ;
assign n51160 =  ( n10 ) ? ( n31656 ) : ( n51159 ) ;
assign n51161 =  ( n148 ) ? ( n32694 ) : ( VREG_9_8 ) ;
assign n51162 =  ( n146 ) ? ( n32693 ) : ( n51161 ) ;
assign n51163 =  ( n144 ) ? ( n32692 ) : ( n51162 ) ;
assign n51164 =  ( n142 ) ? ( n32691 ) : ( n51163 ) ;
assign n51165 =  ( n10 ) ? ( n32690 ) : ( n51164 ) ;
assign n51166 =  ( n32701 ) ? ( VREG_9_8 ) : ( n51160 ) ;
assign n51167 =  ( n32701 ) ? ( VREG_9_8 ) : ( n51165 ) ;
assign n51168 =  ( n3034 ) ? ( n51167 ) : ( VREG_9_8 ) ;
assign n51169 =  ( n2965 ) ? ( n51166 ) : ( n51168 ) ;
assign n51170 =  ( n1930 ) ? ( n51165 ) : ( n51169 ) ;
assign n51171 =  ( n879 ) ? ( n51160 ) : ( n51170 ) ;
assign n51172 =  ( n172 ) ? ( n32712 ) : ( VREG_9_8 ) ;
assign n51173 =  ( n170 ) ? ( n32711 ) : ( n51172 ) ;
assign n51174 =  ( n168 ) ? ( n32710 ) : ( n51173 ) ;
assign n51175 =  ( n166 ) ? ( n32709 ) : ( n51174 ) ;
assign n51176 =  ( n162 ) ? ( n32708 ) : ( n51175 ) ;
assign n51177 =  ( n172 ) ? ( n32722 ) : ( VREG_9_8 ) ;
assign n51178 =  ( n170 ) ? ( n32721 ) : ( n51177 ) ;
assign n51179 =  ( n168 ) ? ( n32720 ) : ( n51178 ) ;
assign n51180 =  ( n166 ) ? ( n32719 ) : ( n51179 ) ;
assign n51181 =  ( n162 ) ? ( n32718 ) : ( n51180 ) ;
assign n51182 =  ( n32701 ) ? ( VREG_9_8 ) : ( n51181 ) ;
assign n51183 =  ( n3051 ) ? ( n51182 ) : ( VREG_9_8 ) ;
assign n51184 =  ( n3040 ) ? ( n51176 ) : ( n51183 ) ;
assign n51185 =  ( n192 ) ? ( VREG_9_8 ) : ( VREG_9_8 ) ;
assign n51186 =  ( n157 ) ? ( n51184 ) : ( n51185 ) ;
assign n51187 =  ( n6 ) ? ( n51171 ) : ( n51186 ) ;
assign n51188 =  ( n857 ) ? ( n51187 ) : ( VREG_9_8 ) ;
assign n51189 =  ( n148 ) ? ( n33779 ) : ( VREG_9_9 ) ;
assign n51190 =  ( n146 ) ? ( n33778 ) : ( n51189 ) ;
assign n51191 =  ( n144 ) ? ( n33777 ) : ( n51190 ) ;
assign n51192 =  ( n142 ) ? ( n33776 ) : ( n51191 ) ;
assign n51193 =  ( n10 ) ? ( n33775 ) : ( n51192 ) ;
assign n51194 =  ( n148 ) ? ( n34813 ) : ( VREG_9_9 ) ;
assign n51195 =  ( n146 ) ? ( n34812 ) : ( n51194 ) ;
assign n51196 =  ( n144 ) ? ( n34811 ) : ( n51195 ) ;
assign n51197 =  ( n142 ) ? ( n34810 ) : ( n51196 ) ;
assign n51198 =  ( n10 ) ? ( n34809 ) : ( n51197 ) ;
assign n51199 =  ( n34820 ) ? ( VREG_9_9 ) : ( n51193 ) ;
assign n51200 =  ( n34820 ) ? ( VREG_9_9 ) : ( n51198 ) ;
assign n51201 =  ( n3034 ) ? ( n51200 ) : ( VREG_9_9 ) ;
assign n51202 =  ( n2965 ) ? ( n51199 ) : ( n51201 ) ;
assign n51203 =  ( n1930 ) ? ( n51198 ) : ( n51202 ) ;
assign n51204 =  ( n879 ) ? ( n51193 ) : ( n51203 ) ;
assign n51205 =  ( n172 ) ? ( n34831 ) : ( VREG_9_9 ) ;
assign n51206 =  ( n170 ) ? ( n34830 ) : ( n51205 ) ;
assign n51207 =  ( n168 ) ? ( n34829 ) : ( n51206 ) ;
assign n51208 =  ( n166 ) ? ( n34828 ) : ( n51207 ) ;
assign n51209 =  ( n162 ) ? ( n34827 ) : ( n51208 ) ;
assign n51210 =  ( n172 ) ? ( n34841 ) : ( VREG_9_9 ) ;
assign n51211 =  ( n170 ) ? ( n34840 ) : ( n51210 ) ;
assign n51212 =  ( n168 ) ? ( n34839 ) : ( n51211 ) ;
assign n51213 =  ( n166 ) ? ( n34838 ) : ( n51212 ) ;
assign n51214 =  ( n162 ) ? ( n34837 ) : ( n51213 ) ;
assign n51215 =  ( n34820 ) ? ( VREG_9_9 ) : ( n51214 ) ;
assign n51216 =  ( n3051 ) ? ( n51215 ) : ( VREG_9_9 ) ;
assign n51217 =  ( n3040 ) ? ( n51209 ) : ( n51216 ) ;
assign n51218 =  ( n192 ) ? ( VREG_9_9 ) : ( VREG_9_9 ) ;
assign n51219 =  ( n157 ) ? ( n51217 ) : ( n51218 ) ;
assign n51220 =  ( n6 ) ? ( n51204 ) : ( n51219 ) ;
assign n51221 =  ( n857 ) ? ( n51220 ) : ( VREG_9_9 ) ;
assign n51222 =  ( pc ) + ( 32'd4 )  ;
always @(posedge clk, posedge rst) begin
   if(rst) begin
       SREG_0 <= SREG_0;
       SREG_1 <= SREG_1;
       SREG_10 <= SREG_10;
       SREG_11 <= SREG_11;
       SREG_12 <= SREG_12;
       SREG_13 <= SREG_13;
       SREG_14 <= SREG_14;
       SREG_15 <= SREG_15;
       SREG_16 <= SREG_16;
       SREG_17 <= SREG_17;
       SREG_18 <= SREG_18;
       SREG_19 <= SREG_19;
       SREG_2 <= SREG_2;
       SREG_20 <= SREG_20;
       SREG_21 <= SREG_21;
       SREG_22 <= SREG_22;
       SREG_23 <= SREG_23;
       SREG_24 <= SREG_24;
       SREG_25 <= SREG_25;
       SREG_26 <= SREG_26;
       SREG_27 <= SREG_27;
       SREG_28 <= SREG_28;
       SREG_29 <= SREG_29;
       SREG_3 <= SREG_3;
       SREG_30 <= SREG_30;
       SREG_31 <= SREG_31;
       SREG_4 <= SREG_4;
       SREG_5 <= SREG_5;
       SREG_6 <= SREG_6;
       SREG_7 <= SREG_7;
       SREG_8 <= SREG_8;
       SREG_9 <= SREG_9;
       VREG_0_0 <= VREG_0_0;
       VREG_0_1 <= VREG_0_1;
       VREG_0_10 <= VREG_0_10;
       VREG_0_11 <= VREG_0_11;
       VREG_0_12 <= VREG_0_12;
       VREG_0_13 <= VREG_0_13;
       VREG_0_14 <= VREG_0_14;
       VREG_0_15 <= VREG_0_15;
       VREG_0_2 <= VREG_0_2;
       VREG_0_3 <= VREG_0_3;
       VREG_0_4 <= VREG_0_4;
       VREG_0_5 <= VREG_0_5;
       VREG_0_6 <= VREG_0_6;
       VREG_0_7 <= VREG_0_7;
       VREG_0_8 <= VREG_0_8;
       VREG_0_9 <= VREG_0_9;
       VREG_10_0 <= VREG_10_0;
       VREG_10_1 <= VREG_10_1;
       VREG_10_10 <= VREG_10_10;
       VREG_10_11 <= VREG_10_11;
       VREG_10_12 <= VREG_10_12;
       VREG_10_13 <= VREG_10_13;
       VREG_10_14 <= VREG_10_14;
       VREG_10_15 <= VREG_10_15;
       VREG_10_2 <= VREG_10_2;
       VREG_10_3 <= VREG_10_3;
       VREG_10_4 <= VREG_10_4;
       VREG_10_5 <= VREG_10_5;
       VREG_10_6 <= VREG_10_6;
       VREG_10_7 <= VREG_10_7;
       VREG_10_8 <= VREG_10_8;
       VREG_10_9 <= VREG_10_9;
       VREG_11_0 <= VREG_11_0;
       VREG_11_1 <= VREG_11_1;
       VREG_11_10 <= VREG_11_10;
       VREG_11_11 <= VREG_11_11;
       VREG_11_12 <= VREG_11_12;
       VREG_11_13 <= VREG_11_13;
       VREG_11_14 <= VREG_11_14;
       VREG_11_15 <= VREG_11_15;
       VREG_11_2 <= VREG_11_2;
       VREG_11_3 <= VREG_11_3;
       VREG_11_4 <= VREG_11_4;
       VREG_11_5 <= VREG_11_5;
       VREG_11_6 <= VREG_11_6;
       VREG_11_7 <= VREG_11_7;
       VREG_11_8 <= VREG_11_8;
       VREG_11_9 <= VREG_11_9;
       VREG_12_0 <= VREG_12_0;
       VREG_12_1 <= VREG_12_1;
       VREG_12_10 <= VREG_12_10;
       VREG_12_11 <= VREG_12_11;
       VREG_12_12 <= VREG_12_12;
       VREG_12_13 <= VREG_12_13;
       VREG_12_14 <= VREG_12_14;
       VREG_12_15 <= VREG_12_15;
       VREG_12_2 <= VREG_12_2;
       VREG_12_3 <= VREG_12_3;
       VREG_12_4 <= VREG_12_4;
       VREG_12_5 <= VREG_12_5;
       VREG_12_6 <= VREG_12_6;
       VREG_12_7 <= VREG_12_7;
       VREG_12_8 <= VREG_12_8;
       VREG_12_9 <= VREG_12_9;
       VREG_13_0 <= VREG_13_0;
       VREG_13_1 <= VREG_13_1;
       VREG_13_10 <= VREG_13_10;
       VREG_13_11 <= VREG_13_11;
       VREG_13_12 <= VREG_13_12;
       VREG_13_13 <= VREG_13_13;
       VREG_13_14 <= VREG_13_14;
       VREG_13_15 <= VREG_13_15;
       VREG_13_2 <= VREG_13_2;
       VREG_13_3 <= VREG_13_3;
       VREG_13_4 <= VREG_13_4;
       VREG_13_5 <= VREG_13_5;
       VREG_13_6 <= VREG_13_6;
       VREG_13_7 <= VREG_13_7;
       VREG_13_8 <= VREG_13_8;
       VREG_13_9 <= VREG_13_9;
       VREG_14_0 <= VREG_14_0;
       VREG_14_1 <= VREG_14_1;
       VREG_14_10 <= VREG_14_10;
       VREG_14_11 <= VREG_14_11;
       VREG_14_12 <= VREG_14_12;
       VREG_14_13 <= VREG_14_13;
       VREG_14_14 <= VREG_14_14;
       VREG_14_15 <= VREG_14_15;
       VREG_14_2 <= VREG_14_2;
       VREG_14_3 <= VREG_14_3;
       VREG_14_4 <= VREG_14_4;
       VREG_14_5 <= VREG_14_5;
       VREG_14_6 <= VREG_14_6;
       VREG_14_7 <= VREG_14_7;
       VREG_14_8 <= VREG_14_8;
       VREG_14_9 <= VREG_14_9;
       VREG_15_0 <= VREG_15_0;
       VREG_15_1 <= VREG_15_1;
       VREG_15_10 <= VREG_15_10;
       VREG_15_11 <= VREG_15_11;
       VREG_15_12 <= VREG_15_12;
       VREG_15_13 <= VREG_15_13;
       VREG_15_14 <= VREG_15_14;
       VREG_15_15 <= VREG_15_15;
       VREG_15_2 <= VREG_15_2;
       VREG_15_3 <= VREG_15_3;
       VREG_15_4 <= VREG_15_4;
       VREG_15_5 <= VREG_15_5;
       VREG_15_6 <= VREG_15_6;
       VREG_15_7 <= VREG_15_7;
       VREG_15_8 <= VREG_15_8;
       VREG_15_9 <= VREG_15_9;
       VREG_16_0 <= VREG_16_0;
       VREG_16_1 <= VREG_16_1;
       VREG_16_10 <= VREG_16_10;
       VREG_16_11 <= VREG_16_11;
       VREG_16_12 <= VREG_16_12;
       VREG_16_13 <= VREG_16_13;
       VREG_16_14 <= VREG_16_14;
       VREG_16_15 <= VREG_16_15;
       VREG_16_2 <= VREG_16_2;
       VREG_16_3 <= VREG_16_3;
       VREG_16_4 <= VREG_16_4;
       VREG_16_5 <= VREG_16_5;
       VREG_16_6 <= VREG_16_6;
       VREG_16_7 <= VREG_16_7;
       VREG_16_8 <= VREG_16_8;
       VREG_16_9 <= VREG_16_9;
       VREG_17_0 <= VREG_17_0;
       VREG_17_1 <= VREG_17_1;
       VREG_17_10 <= VREG_17_10;
       VREG_17_11 <= VREG_17_11;
       VREG_17_12 <= VREG_17_12;
       VREG_17_13 <= VREG_17_13;
       VREG_17_14 <= VREG_17_14;
       VREG_17_15 <= VREG_17_15;
       VREG_17_2 <= VREG_17_2;
       VREG_17_3 <= VREG_17_3;
       VREG_17_4 <= VREG_17_4;
       VREG_17_5 <= VREG_17_5;
       VREG_17_6 <= VREG_17_6;
       VREG_17_7 <= VREG_17_7;
       VREG_17_8 <= VREG_17_8;
       VREG_17_9 <= VREG_17_9;
       VREG_18_0 <= VREG_18_0;
       VREG_18_1 <= VREG_18_1;
       VREG_18_10 <= VREG_18_10;
       VREG_18_11 <= VREG_18_11;
       VREG_18_12 <= VREG_18_12;
       VREG_18_13 <= VREG_18_13;
       VREG_18_14 <= VREG_18_14;
       VREG_18_15 <= VREG_18_15;
       VREG_18_2 <= VREG_18_2;
       VREG_18_3 <= VREG_18_3;
       VREG_18_4 <= VREG_18_4;
       VREG_18_5 <= VREG_18_5;
       VREG_18_6 <= VREG_18_6;
       VREG_18_7 <= VREG_18_7;
       VREG_18_8 <= VREG_18_8;
       VREG_18_9 <= VREG_18_9;
       VREG_19_0 <= VREG_19_0;
       VREG_19_1 <= VREG_19_1;
       VREG_19_10 <= VREG_19_10;
       VREG_19_11 <= VREG_19_11;
       VREG_19_12 <= VREG_19_12;
       VREG_19_13 <= VREG_19_13;
       VREG_19_14 <= VREG_19_14;
       VREG_19_15 <= VREG_19_15;
       VREG_19_2 <= VREG_19_2;
       VREG_19_3 <= VREG_19_3;
       VREG_19_4 <= VREG_19_4;
       VREG_19_5 <= VREG_19_5;
       VREG_19_6 <= VREG_19_6;
       VREG_19_7 <= VREG_19_7;
       VREG_19_8 <= VREG_19_8;
       VREG_19_9 <= VREG_19_9;
       VREG_1_0 <= VREG_1_0;
       VREG_1_1 <= VREG_1_1;
       VREG_1_10 <= VREG_1_10;
       VREG_1_11 <= VREG_1_11;
       VREG_1_12 <= VREG_1_12;
       VREG_1_13 <= VREG_1_13;
       VREG_1_14 <= VREG_1_14;
       VREG_1_15 <= VREG_1_15;
       VREG_1_2 <= VREG_1_2;
       VREG_1_3 <= VREG_1_3;
       VREG_1_4 <= VREG_1_4;
       VREG_1_5 <= VREG_1_5;
       VREG_1_6 <= VREG_1_6;
       VREG_1_7 <= VREG_1_7;
       VREG_1_8 <= VREG_1_8;
       VREG_1_9 <= VREG_1_9;
       VREG_20_0 <= VREG_20_0;
       VREG_20_1 <= VREG_20_1;
       VREG_20_10 <= VREG_20_10;
       VREG_20_11 <= VREG_20_11;
       VREG_20_12 <= VREG_20_12;
       VREG_20_13 <= VREG_20_13;
       VREG_20_14 <= VREG_20_14;
       VREG_20_15 <= VREG_20_15;
       VREG_20_2 <= VREG_20_2;
       VREG_20_3 <= VREG_20_3;
       VREG_20_4 <= VREG_20_4;
       VREG_20_5 <= VREG_20_5;
       VREG_20_6 <= VREG_20_6;
       VREG_20_7 <= VREG_20_7;
       VREG_20_8 <= VREG_20_8;
       VREG_20_9 <= VREG_20_9;
       VREG_21_0 <= VREG_21_0;
       VREG_21_1 <= VREG_21_1;
       VREG_21_10 <= VREG_21_10;
       VREG_21_11 <= VREG_21_11;
       VREG_21_12 <= VREG_21_12;
       VREG_21_13 <= VREG_21_13;
       VREG_21_14 <= VREG_21_14;
       VREG_21_15 <= VREG_21_15;
       VREG_21_2 <= VREG_21_2;
       VREG_21_3 <= VREG_21_3;
       VREG_21_4 <= VREG_21_4;
       VREG_21_5 <= VREG_21_5;
       VREG_21_6 <= VREG_21_6;
       VREG_21_7 <= VREG_21_7;
       VREG_21_8 <= VREG_21_8;
       VREG_21_9 <= VREG_21_9;
       VREG_22_0 <= VREG_22_0;
       VREG_22_1 <= VREG_22_1;
       VREG_22_10 <= VREG_22_10;
       VREG_22_11 <= VREG_22_11;
       VREG_22_12 <= VREG_22_12;
       VREG_22_13 <= VREG_22_13;
       VREG_22_14 <= VREG_22_14;
       VREG_22_15 <= VREG_22_15;
       VREG_22_2 <= VREG_22_2;
       VREG_22_3 <= VREG_22_3;
       VREG_22_4 <= VREG_22_4;
       VREG_22_5 <= VREG_22_5;
       VREG_22_6 <= VREG_22_6;
       VREG_22_7 <= VREG_22_7;
       VREG_22_8 <= VREG_22_8;
       VREG_22_9 <= VREG_22_9;
       VREG_23_0 <= VREG_23_0;
       VREG_23_1 <= VREG_23_1;
       VREG_23_10 <= VREG_23_10;
       VREG_23_11 <= VREG_23_11;
       VREG_23_12 <= VREG_23_12;
       VREG_23_13 <= VREG_23_13;
       VREG_23_14 <= VREG_23_14;
       VREG_23_15 <= VREG_23_15;
       VREG_23_2 <= VREG_23_2;
       VREG_23_3 <= VREG_23_3;
       VREG_23_4 <= VREG_23_4;
       VREG_23_5 <= VREG_23_5;
       VREG_23_6 <= VREG_23_6;
       VREG_23_7 <= VREG_23_7;
       VREG_23_8 <= VREG_23_8;
       VREG_23_9 <= VREG_23_9;
       VREG_24_0 <= VREG_24_0;
       VREG_24_1 <= VREG_24_1;
       VREG_24_10 <= VREG_24_10;
       VREG_24_11 <= VREG_24_11;
       VREG_24_12 <= VREG_24_12;
       VREG_24_13 <= VREG_24_13;
       VREG_24_14 <= VREG_24_14;
       VREG_24_15 <= VREG_24_15;
       VREG_24_2 <= VREG_24_2;
       VREG_24_3 <= VREG_24_3;
       VREG_24_4 <= VREG_24_4;
       VREG_24_5 <= VREG_24_5;
       VREG_24_6 <= VREG_24_6;
       VREG_24_7 <= VREG_24_7;
       VREG_24_8 <= VREG_24_8;
       VREG_24_9 <= VREG_24_9;
       VREG_25_0 <= VREG_25_0;
       VREG_25_1 <= VREG_25_1;
       VREG_25_10 <= VREG_25_10;
       VREG_25_11 <= VREG_25_11;
       VREG_25_12 <= VREG_25_12;
       VREG_25_13 <= VREG_25_13;
       VREG_25_14 <= VREG_25_14;
       VREG_25_15 <= VREG_25_15;
       VREG_25_2 <= VREG_25_2;
       VREG_25_3 <= VREG_25_3;
       VREG_25_4 <= VREG_25_4;
       VREG_25_5 <= VREG_25_5;
       VREG_25_6 <= VREG_25_6;
       VREG_25_7 <= VREG_25_7;
       VREG_25_8 <= VREG_25_8;
       VREG_25_9 <= VREG_25_9;
       VREG_26_0 <= VREG_26_0;
       VREG_26_1 <= VREG_26_1;
       VREG_26_10 <= VREG_26_10;
       VREG_26_11 <= VREG_26_11;
       VREG_26_12 <= VREG_26_12;
       VREG_26_13 <= VREG_26_13;
       VREG_26_14 <= VREG_26_14;
       VREG_26_15 <= VREG_26_15;
       VREG_26_2 <= VREG_26_2;
       VREG_26_3 <= VREG_26_3;
       VREG_26_4 <= VREG_26_4;
       VREG_26_5 <= VREG_26_5;
       VREG_26_6 <= VREG_26_6;
       VREG_26_7 <= VREG_26_7;
       VREG_26_8 <= VREG_26_8;
       VREG_26_9 <= VREG_26_9;
       VREG_27_0 <= VREG_27_0;
       VREG_27_1 <= VREG_27_1;
       VREG_27_10 <= VREG_27_10;
       VREG_27_11 <= VREG_27_11;
       VREG_27_12 <= VREG_27_12;
       VREG_27_13 <= VREG_27_13;
       VREG_27_14 <= VREG_27_14;
       VREG_27_15 <= VREG_27_15;
       VREG_27_2 <= VREG_27_2;
       VREG_27_3 <= VREG_27_3;
       VREG_27_4 <= VREG_27_4;
       VREG_27_5 <= VREG_27_5;
       VREG_27_6 <= VREG_27_6;
       VREG_27_7 <= VREG_27_7;
       VREG_27_8 <= VREG_27_8;
       VREG_27_9 <= VREG_27_9;
       VREG_28_0 <= VREG_28_0;
       VREG_28_1 <= VREG_28_1;
       VREG_28_10 <= VREG_28_10;
       VREG_28_11 <= VREG_28_11;
       VREG_28_12 <= VREG_28_12;
       VREG_28_13 <= VREG_28_13;
       VREG_28_14 <= VREG_28_14;
       VREG_28_15 <= VREG_28_15;
       VREG_28_2 <= VREG_28_2;
       VREG_28_3 <= VREG_28_3;
       VREG_28_4 <= VREG_28_4;
       VREG_28_5 <= VREG_28_5;
       VREG_28_6 <= VREG_28_6;
       VREG_28_7 <= VREG_28_7;
       VREG_28_8 <= VREG_28_8;
       VREG_28_9 <= VREG_28_9;
       VREG_29_0 <= VREG_29_0;
       VREG_29_1 <= VREG_29_1;
       VREG_29_10 <= VREG_29_10;
       VREG_29_11 <= VREG_29_11;
       VREG_29_12 <= VREG_29_12;
       VREG_29_13 <= VREG_29_13;
       VREG_29_14 <= VREG_29_14;
       VREG_29_15 <= VREG_29_15;
       VREG_29_2 <= VREG_29_2;
       VREG_29_3 <= VREG_29_3;
       VREG_29_4 <= VREG_29_4;
       VREG_29_5 <= VREG_29_5;
       VREG_29_6 <= VREG_29_6;
       VREG_29_7 <= VREG_29_7;
       VREG_29_8 <= VREG_29_8;
       VREG_29_9 <= VREG_29_9;
       VREG_2_0 <= VREG_2_0;
       VREG_2_1 <= VREG_2_1;
       VREG_2_10 <= VREG_2_10;
       VREG_2_11 <= VREG_2_11;
       VREG_2_12 <= VREG_2_12;
       VREG_2_13 <= VREG_2_13;
       VREG_2_14 <= VREG_2_14;
       VREG_2_15 <= VREG_2_15;
       VREG_2_2 <= VREG_2_2;
       VREG_2_3 <= VREG_2_3;
       VREG_2_4 <= VREG_2_4;
       VREG_2_5 <= VREG_2_5;
       VREG_2_6 <= VREG_2_6;
       VREG_2_7 <= VREG_2_7;
       VREG_2_8 <= VREG_2_8;
       VREG_2_9 <= VREG_2_9;
       VREG_30_0 <= VREG_30_0;
       VREG_30_1 <= VREG_30_1;
       VREG_30_10 <= VREG_30_10;
       VREG_30_11 <= VREG_30_11;
       VREG_30_12 <= VREG_30_12;
       VREG_30_13 <= VREG_30_13;
       VREG_30_14 <= VREG_30_14;
       VREG_30_15 <= VREG_30_15;
       VREG_30_2 <= VREG_30_2;
       VREG_30_3 <= VREG_30_3;
       VREG_30_4 <= VREG_30_4;
       VREG_30_5 <= VREG_30_5;
       VREG_30_6 <= VREG_30_6;
       VREG_30_7 <= VREG_30_7;
       VREG_30_8 <= VREG_30_8;
       VREG_30_9 <= VREG_30_9;
       VREG_31_0 <= VREG_31_0;
       VREG_31_1 <= VREG_31_1;
       VREG_31_10 <= VREG_31_10;
       VREG_31_11 <= VREG_31_11;
       VREG_31_12 <= VREG_31_12;
       VREG_31_13 <= VREG_31_13;
       VREG_31_14 <= VREG_31_14;
       VREG_31_15 <= VREG_31_15;
       VREG_31_2 <= VREG_31_2;
       VREG_31_3 <= VREG_31_3;
       VREG_31_4 <= VREG_31_4;
       VREG_31_5 <= VREG_31_5;
       VREG_31_6 <= VREG_31_6;
       VREG_31_7 <= VREG_31_7;
       VREG_31_8 <= VREG_31_8;
       VREG_31_9 <= VREG_31_9;
       VREG_3_0 <= VREG_3_0;
       VREG_3_1 <= VREG_3_1;
       VREG_3_10 <= VREG_3_10;
       VREG_3_11 <= VREG_3_11;
       VREG_3_12 <= VREG_3_12;
       VREG_3_13 <= VREG_3_13;
       VREG_3_14 <= VREG_3_14;
       VREG_3_15 <= VREG_3_15;
       VREG_3_2 <= VREG_3_2;
       VREG_3_3 <= VREG_3_3;
       VREG_3_4 <= VREG_3_4;
       VREG_3_5 <= VREG_3_5;
       VREG_3_6 <= VREG_3_6;
       VREG_3_7 <= VREG_3_7;
       VREG_3_8 <= VREG_3_8;
       VREG_3_9 <= VREG_3_9;
       VREG_4_0 <= VREG_4_0;
       VREG_4_1 <= VREG_4_1;
       VREG_4_10 <= VREG_4_10;
       VREG_4_11 <= VREG_4_11;
       VREG_4_12 <= VREG_4_12;
       VREG_4_13 <= VREG_4_13;
       VREG_4_14 <= VREG_4_14;
       VREG_4_15 <= VREG_4_15;
       VREG_4_2 <= VREG_4_2;
       VREG_4_3 <= VREG_4_3;
       VREG_4_4 <= VREG_4_4;
       VREG_4_5 <= VREG_4_5;
       VREG_4_6 <= VREG_4_6;
       VREG_4_7 <= VREG_4_7;
       VREG_4_8 <= VREG_4_8;
       VREG_4_9 <= VREG_4_9;
       VREG_5_0 <= VREG_5_0;
       VREG_5_1 <= VREG_5_1;
       VREG_5_10 <= VREG_5_10;
       VREG_5_11 <= VREG_5_11;
       VREG_5_12 <= VREG_5_12;
       VREG_5_13 <= VREG_5_13;
       VREG_5_14 <= VREG_5_14;
       VREG_5_15 <= VREG_5_15;
       VREG_5_2 <= VREG_5_2;
       VREG_5_3 <= VREG_5_3;
       VREG_5_4 <= VREG_5_4;
       VREG_5_5 <= VREG_5_5;
       VREG_5_6 <= VREG_5_6;
       VREG_5_7 <= VREG_5_7;
       VREG_5_8 <= VREG_5_8;
       VREG_5_9 <= VREG_5_9;
       VREG_6_0 <= VREG_6_0;
       VREG_6_1 <= VREG_6_1;
       VREG_6_10 <= VREG_6_10;
       VREG_6_11 <= VREG_6_11;
       VREG_6_12 <= VREG_6_12;
       VREG_6_13 <= VREG_6_13;
       VREG_6_14 <= VREG_6_14;
       VREG_6_15 <= VREG_6_15;
       VREG_6_2 <= VREG_6_2;
       VREG_6_3 <= VREG_6_3;
       VREG_6_4 <= VREG_6_4;
       VREG_6_5 <= VREG_6_5;
       VREG_6_6 <= VREG_6_6;
       VREG_6_7 <= VREG_6_7;
       VREG_6_8 <= VREG_6_8;
       VREG_6_9 <= VREG_6_9;
       VREG_7_0 <= VREG_7_0;
       VREG_7_1 <= VREG_7_1;
       VREG_7_10 <= VREG_7_10;
       VREG_7_11 <= VREG_7_11;
       VREG_7_12 <= VREG_7_12;
       VREG_7_13 <= VREG_7_13;
       VREG_7_14 <= VREG_7_14;
       VREG_7_15 <= VREG_7_15;
       VREG_7_2 <= VREG_7_2;
       VREG_7_3 <= VREG_7_3;
       VREG_7_4 <= VREG_7_4;
       VREG_7_5 <= VREG_7_5;
       VREG_7_6 <= VREG_7_6;
       VREG_7_7 <= VREG_7_7;
       VREG_7_8 <= VREG_7_8;
       VREG_7_9 <= VREG_7_9;
       VREG_8_0 <= VREG_8_0;
       VREG_8_1 <= VREG_8_1;
       VREG_8_10 <= VREG_8_10;
       VREG_8_11 <= VREG_8_11;
       VREG_8_12 <= VREG_8_12;
       VREG_8_13 <= VREG_8_13;
       VREG_8_14 <= VREG_8_14;
       VREG_8_15 <= VREG_8_15;
       VREG_8_2 <= VREG_8_2;
       VREG_8_3 <= VREG_8_3;
       VREG_8_4 <= VREG_8_4;
       VREG_8_5 <= VREG_8_5;
       VREG_8_6 <= VREG_8_6;
       VREG_8_7 <= VREG_8_7;
       VREG_8_8 <= VREG_8_8;
       VREG_8_9 <= VREG_8_9;
       VREG_9_0 <= VREG_9_0;
       VREG_9_1 <= VREG_9_1;
       VREG_9_10 <= VREG_9_10;
       VREG_9_11 <= VREG_9_11;
       VREG_9_12 <= VREG_9_12;
       VREG_9_13 <= VREG_9_13;
       VREG_9_14 <= VREG_9_14;
       VREG_9_15 <= VREG_9_15;
       VREG_9_2 <= VREG_9_2;
       VREG_9_3 <= VREG_9_3;
       VREG_9_4 <= VREG_9_4;
       VREG_9_5 <= VREG_9_5;
       VREG_9_6 <= VREG_9_6;
       VREG_9_7 <= VREG_9_7;
       VREG_9_8 <= VREG_9_8;
       VREG_9_9 <= VREG_9_9;
       pc <= pc;
       vector_mask_register <= vector_mask_register;
   end
   else if(step) begin
       SREG_0 <= n196;
       SREG_1 <= n218;
       SREG_10 <= n240;
       SREG_11 <= n262;
       SREG_12 <= n284;
       SREG_13 <= n306;
       SREG_14 <= n328;
       SREG_15 <= n350;
       SREG_16 <= n372;
       SREG_17 <= n394;
       SREG_18 <= n416;
       SREG_19 <= n438;
       SREG_2 <= n460;
       SREG_20 <= n482;
       SREG_21 <= n504;
       SREG_22 <= n526;
       SREG_23 <= n548;
       SREG_24 <= n570;
       SREG_25 <= n592;
       SREG_26 <= n614;
       SREG_27 <= n636;
       SREG_28 <= n658;
       SREG_29 <= n680;
       SREG_3 <= n702;
       SREG_30 <= n724;
       SREG_31 <= n746;
       SREG_4 <= n768;
       SREG_5 <= n790;
       SREG_6 <= n812;
       SREG_7 <= n834;
       SREG_8 <= n856;
       SREG_9 <= n878;
       VREG_0_0 <= n3068;
       VREG_0_1 <= n5187;
       VREG_0_10 <= n7306;
       VREG_0_11 <= n9425;
       VREG_0_12 <= n11544;
       VREG_0_13 <= n13663;
       VREG_0_14 <= n15782;
       VREG_0_15 <= n17901;
       VREG_0_2 <= n20020;
       VREG_0_3 <= n22139;
       VREG_0_4 <= n24258;
       VREG_0_5 <= n26377;
       VREG_0_6 <= n28496;
       VREG_0_7 <= n30615;
       VREG_0_8 <= n32734;
       VREG_0_9 <= n34853;
       VREG_10_0 <= n34886;
       VREG_10_1 <= n34919;
       VREG_10_10 <= n34952;
       VREG_10_11 <= n34985;
       VREG_10_12 <= n35018;
       VREG_10_13 <= n35051;
       VREG_10_14 <= n35084;
       VREG_10_15 <= n35117;
       VREG_10_2 <= n35150;
       VREG_10_3 <= n35183;
       VREG_10_4 <= n35216;
       VREG_10_5 <= n35249;
       VREG_10_6 <= n35282;
       VREG_10_7 <= n35315;
       VREG_10_8 <= n35348;
       VREG_10_9 <= n35381;
       VREG_11_0 <= n35414;
       VREG_11_1 <= n35447;
       VREG_11_10 <= n35480;
       VREG_11_11 <= n35513;
       VREG_11_12 <= n35546;
       VREG_11_13 <= n35579;
       VREG_11_14 <= n35612;
       VREG_11_15 <= n35645;
       VREG_11_2 <= n35678;
       VREG_11_3 <= n35711;
       VREG_11_4 <= n35744;
       VREG_11_5 <= n35777;
       VREG_11_6 <= n35810;
       VREG_11_7 <= n35843;
       VREG_11_8 <= n35876;
       VREG_11_9 <= n35909;
       VREG_12_0 <= n35942;
       VREG_12_1 <= n35975;
       VREG_12_10 <= n36008;
       VREG_12_11 <= n36041;
       VREG_12_12 <= n36074;
       VREG_12_13 <= n36107;
       VREG_12_14 <= n36140;
       VREG_12_15 <= n36173;
       VREG_12_2 <= n36206;
       VREG_12_3 <= n36239;
       VREG_12_4 <= n36272;
       VREG_12_5 <= n36305;
       VREG_12_6 <= n36338;
       VREG_12_7 <= n36371;
       VREG_12_8 <= n36404;
       VREG_12_9 <= n36437;
       VREG_13_0 <= n36470;
       VREG_13_1 <= n36503;
       VREG_13_10 <= n36536;
       VREG_13_11 <= n36569;
       VREG_13_12 <= n36602;
       VREG_13_13 <= n36635;
       VREG_13_14 <= n36668;
       VREG_13_15 <= n36701;
       VREG_13_2 <= n36734;
       VREG_13_3 <= n36767;
       VREG_13_4 <= n36800;
       VREG_13_5 <= n36833;
       VREG_13_6 <= n36866;
       VREG_13_7 <= n36899;
       VREG_13_8 <= n36932;
       VREG_13_9 <= n36965;
       VREG_14_0 <= n36998;
       VREG_14_1 <= n37031;
       VREG_14_10 <= n37064;
       VREG_14_11 <= n37097;
       VREG_14_12 <= n37130;
       VREG_14_13 <= n37163;
       VREG_14_14 <= n37196;
       VREG_14_15 <= n37229;
       VREG_14_2 <= n37262;
       VREG_14_3 <= n37295;
       VREG_14_4 <= n37328;
       VREG_14_5 <= n37361;
       VREG_14_6 <= n37394;
       VREG_14_7 <= n37427;
       VREG_14_8 <= n37460;
       VREG_14_9 <= n37493;
       VREG_15_0 <= n37526;
       VREG_15_1 <= n37559;
       VREG_15_10 <= n37592;
       VREG_15_11 <= n37625;
       VREG_15_12 <= n37658;
       VREG_15_13 <= n37691;
       VREG_15_14 <= n37724;
       VREG_15_15 <= n37757;
       VREG_15_2 <= n37790;
       VREG_15_3 <= n37823;
       VREG_15_4 <= n37856;
       VREG_15_5 <= n37889;
       VREG_15_6 <= n37922;
       VREG_15_7 <= n37955;
       VREG_15_8 <= n37988;
       VREG_15_9 <= n38021;
       VREG_16_0 <= n38054;
       VREG_16_1 <= n38087;
       VREG_16_10 <= n38120;
       VREG_16_11 <= n38153;
       VREG_16_12 <= n38186;
       VREG_16_13 <= n38219;
       VREG_16_14 <= n38252;
       VREG_16_15 <= n38285;
       VREG_16_2 <= n38318;
       VREG_16_3 <= n38351;
       VREG_16_4 <= n38384;
       VREG_16_5 <= n38417;
       VREG_16_6 <= n38450;
       VREG_16_7 <= n38483;
       VREG_16_8 <= n38516;
       VREG_16_9 <= n38549;
       VREG_17_0 <= n38582;
       VREG_17_1 <= n38615;
       VREG_17_10 <= n38648;
       VREG_17_11 <= n38681;
       VREG_17_12 <= n38714;
       VREG_17_13 <= n38747;
       VREG_17_14 <= n38780;
       VREG_17_15 <= n38813;
       VREG_17_2 <= n38846;
       VREG_17_3 <= n38879;
       VREG_17_4 <= n38912;
       VREG_17_5 <= n38945;
       VREG_17_6 <= n38978;
       VREG_17_7 <= n39011;
       VREG_17_8 <= n39044;
       VREG_17_9 <= n39077;
       VREG_18_0 <= n39110;
       VREG_18_1 <= n39143;
       VREG_18_10 <= n39176;
       VREG_18_11 <= n39209;
       VREG_18_12 <= n39242;
       VREG_18_13 <= n39275;
       VREG_18_14 <= n39308;
       VREG_18_15 <= n39341;
       VREG_18_2 <= n39374;
       VREG_18_3 <= n39407;
       VREG_18_4 <= n39440;
       VREG_18_5 <= n39473;
       VREG_18_6 <= n39506;
       VREG_18_7 <= n39539;
       VREG_18_8 <= n39572;
       VREG_18_9 <= n39605;
       VREG_19_0 <= n39638;
       VREG_19_1 <= n39671;
       VREG_19_10 <= n39704;
       VREG_19_11 <= n39737;
       VREG_19_12 <= n39770;
       VREG_19_13 <= n39803;
       VREG_19_14 <= n39836;
       VREG_19_15 <= n39869;
       VREG_19_2 <= n39902;
       VREG_19_3 <= n39935;
       VREG_19_4 <= n39968;
       VREG_19_5 <= n40001;
       VREG_19_6 <= n40034;
       VREG_19_7 <= n40067;
       VREG_19_8 <= n40100;
       VREG_19_9 <= n40133;
       VREG_1_0 <= n40166;
       VREG_1_1 <= n40199;
       VREG_1_10 <= n40232;
       VREG_1_11 <= n40265;
       VREG_1_12 <= n40298;
       VREG_1_13 <= n40331;
       VREG_1_14 <= n40364;
       VREG_1_15 <= n40397;
       VREG_1_2 <= n40430;
       VREG_1_3 <= n40463;
       VREG_1_4 <= n40496;
       VREG_1_5 <= n40529;
       VREG_1_6 <= n40562;
       VREG_1_7 <= n40595;
       VREG_1_8 <= n40628;
       VREG_1_9 <= n40661;
       VREG_20_0 <= n40694;
       VREG_20_1 <= n40727;
       VREG_20_10 <= n40760;
       VREG_20_11 <= n40793;
       VREG_20_12 <= n40826;
       VREG_20_13 <= n40859;
       VREG_20_14 <= n40892;
       VREG_20_15 <= n40925;
       VREG_20_2 <= n40958;
       VREG_20_3 <= n40991;
       VREG_20_4 <= n41024;
       VREG_20_5 <= n41057;
       VREG_20_6 <= n41090;
       VREG_20_7 <= n41123;
       VREG_20_8 <= n41156;
       VREG_20_9 <= n41189;
       VREG_21_0 <= n41222;
       VREG_21_1 <= n41255;
       VREG_21_10 <= n41288;
       VREG_21_11 <= n41321;
       VREG_21_12 <= n41354;
       VREG_21_13 <= n41387;
       VREG_21_14 <= n41420;
       VREG_21_15 <= n41453;
       VREG_21_2 <= n41486;
       VREG_21_3 <= n41519;
       VREG_21_4 <= n41552;
       VREG_21_5 <= n41585;
       VREG_21_6 <= n41618;
       VREG_21_7 <= n41651;
       VREG_21_8 <= n41684;
       VREG_21_9 <= n41717;
       VREG_22_0 <= n41750;
       VREG_22_1 <= n41783;
       VREG_22_10 <= n41816;
       VREG_22_11 <= n41849;
       VREG_22_12 <= n41882;
       VREG_22_13 <= n41915;
       VREG_22_14 <= n41948;
       VREG_22_15 <= n41981;
       VREG_22_2 <= n42014;
       VREG_22_3 <= n42047;
       VREG_22_4 <= n42080;
       VREG_22_5 <= n42113;
       VREG_22_6 <= n42146;
       VREG_22_7 <= n42179;
       VREG_22_8 <= n42212;
       VREG_22_9 <= n42245;
       VREG_23_0 <= n42278;
       VREG_23_1 <= n42311;
       VREG_23_10 <= n42344;
       VREG_23_11 <= n42377;
       VREG_23_12 <= n42410;
       VREG_23_13 <= n42443;
       VREG_23_14 <= n42476;
       VREG_23_15 <= n42509;
       VREG_23_2 <= n42542;
       VREG_23_3 <= n42575;
       VREG_23_4 <= n42608;
       VREG_23_5 <= n42641;
       VREG_23_6 <= n42674;
       VREG_23_7 <= n42707;
       VREG_23_8 <= n42740;
       VREG_23_9 <= n42773;
       VREG_24_0 <= n42806;
       VREG_24_1 <= n42839;
       VREG_24_10 <= n42872;
       VREG_24_11 <= n42905;
       VREG_24_12 <= n42938;
       VREG_24_13 <= n42971;
       VREG_24_14 <= n43004;
       VREG_24_15 <= n43037;
       VREG_24_2 <= n43070;
       VREG_24_3 <= n43103;
       VREG_24_4 <= n43136;
       VREG_24_5 <= n43169;
       VREG_24_6 <= n43202;
       VREG_24_7 <= n43235;
       VREG_24_8 <= n43268;
       VREG_24_9 <= n43301;
       VREG_25_0 <= n43334;
       VREG_25_1 <= n43367;
       VREG_25_10 <= n43400;
       VREG_25_11 <= n43433;
       VREG_25_12 <= n43466;
       VREG_25_13 <= n43499;
       VREG_25_14 <= n43532;
       VREG_25_15 <= n43565;
       VREG_25_2 <= n43598;
       VREG_25_3 <= n43631;
       VREG_25_4 <= n43664;
       VREG_25_5 <= n43697;
       VREG_25_6 <= n43730;
       VREG_25_7 <= n43763;
       VREG_25_8 <= n43796;
       VREG_25_9 <= n43829;
       VREG_26_0 <= n43862;
       VREG_26_1 <= n43895;
       VREG_26_10 <= n43928;
       VREG_26_11 <= n43961;
       VREG_26_12 <= n43994;
       VREG_26_13 <= n44027;
       VREG_26_14 <= n44060;
       VREG_26_15 <= n44093;
       VREG_26_2 <= n44126;
       VREG_26_3 <= n44159;
       VREG_26_4 <= n44192;
       VREG_26_5 <= n44225;
       VREG_26_6 <= n44258;
       VREG_26_7 <= n44291;
       VREG_26_8 <= n44324;
       VREG_26_9 <= n44357;
       VREG_27_0 <= n44390;
       VREG_27_1 <= n44423;
       VREG_27_10 <= n44456;
       VREG_27_11 <= n44489;
       VREG_27_12 <= n44522;
       VREG_27_13 <= n44555;
       VREG_27_14 <= n44588;
       VREG_27_15 <= n44621;
       VREG_27_2 <= n44654;
       VREG_27_3 <= n44687;
       VREG_27_4 <= n44720;
       VREG_27_5 <= n44753;
       VREG_27_6 <= n44786;
       VREG_27_7 <= n44819;
       VREG_27_8 <= n44852;
       VREG_27_9 <= n44885;
       VREG_28_0 <= n44918;
       VREG_28_1 <= n44951;
       VREG_28_10 <= n44984;
       VREG_28_11 <= n45017;
       VREG_28_12 <= n45050;
       VREG_28_13 <= n45083;
       VREG_28_14 <= n45116;
       VREG_28_15 <= n45149;
       VREG_28_2 <= n45182;
       VREG_28_3 <= n45215;
       VREG_28_4 <= n45248;
       VREG_28_5 <= n45281;
       VREG_28_6 <= n45314;
       VREG_28_7 <= n45347;
       VREG_28_8 <= n45380;
       VREG_28_9 <= n45413;
       VREG_29_0 <= n45446;
       VREG_29_1 <= n45479;
       VREG_29_10 <= n45512;
       VREG_29_11 <= n45545;
       VREG_29_12 <= n45578;
       VREG_29_13 <= n45611;
       VREG_29_14 <= n45644;
       VREG_29_15 <= n45677;
       VREG_29_2 <= n45710;
       VREG_29_3 <= n45743;
       VREG_29_4 <= n45776;
       VREG_29_5 <= n45809;
       VREG_29_6 <= n45842;
       VREG_29_7 <= n45875;
       VREG_29_8 <= n45908;
       VREG_29_9 <= n45941;
       VREG_2_0 <= n45974;
       VREG_2_1 <= n46007;
       VREG_2_10 <= n46040;
       VREG_2_11 <= n46073;
       VREG_2_12 <= n46106;
       VREG_2_13 <= n46139;
       VREG_2_14 <= n46172;
       VREG_2_15 <= n46205;
       VREG_2_2 <= n46238;
       VREG_2_3 <= n46271;
       VREG_2_4 <= n46304;
       VREG_2_5 <= n46337;
       VREG_2_6 <= n46370;
       VREG_2_7 <= n46403;
       VREG_2_8 <= n46436;
       VREG_2_9 <= n46469;
       VREG_30_0 <= n46502;
       VREG_30_1 <= n46535;
       VREG_30_10 <= n46568;
       VREG_30_11 <= n46601;
       VREG_30_12 <= n46634;
       VREG_30_13 <= n46667;
       VREG_30_14 <= n46700;
       VREG_30_15 <= n46733;
       VREG_30_2 <= n46766;
       VREG_30_3 <= n46799;
       VREG_30_4 <= n46832;
       VREG_30_5 <= n46865;
       VREG_30_6 <= n46898;
       VREG_30_7 <= n46931;
       VREG_30_8 <= n46964;
       VREG_30_9 <= n46997;
       VREG_31_0 <= n47030;
       VREG_31_1 <= n47063;
       VREG_31_10 <= n47096;
       VREG_31_11 <= n47129;
       VREG_31_12 <= n47162;
       VREG_31_13 <= n47195;
       VREG_31_14 <= n47228;
       VREG_31_15 <= n47261;
       VREG_31_2 <= n47294;
       VREG_31_3 <= n47327;
       VREG_31_4 <= n47360;
       VREG_31_5 <= n47393;
       VREG_31_6 <= n47426;
       VREG_31_7 <= n47459;
       VREG_31_8 <= n47492;
       VREG_31_9 <= n47525;
       VREG_3_0 <= n47558;
       VREG_3_1 <= n47591;
       VREG_3_10 <= n47624;
       VREG_3_11 <= n47657;
       VREG_3_12 <= n47690;
       VREG_3_13 <= n47723;
       VREG_3_14 <= n47756;
       VREG_3_15 <= n47789;
       VREG_3_2 <= n47822;
       VREG_3_3 <= n47855;
       VREG_3_4 <= n47888;
       VREG_3_5 <= n47921;
       VREG_3_6 <= n47954;
       VREG_3_7 <= n47987;
       VREG_3_8 <= n48020;
       VREG_3_9 <= n48053;
       VREG_4_0 <= n48086;
       VREG_4_1 <= n48119;
       VREG_4_10 <= n48152;
       VREG_4_11 <= n48185;
       VREG_4_12 <= n48218;
       VREG_4_13 <= n48251;
       VREG_4_14 <= n48284;
       VREG_4_15 <= n48317;
       VREG_4_2 <= n48350;
       VREG_4_3 <= n48383;
       VREG_4_4 <= n48416;
       VREG_4_5 <= n48449;
       VREG_4_6 <= n48482;
       VREG_4_7 <= n48515;
       VREG_4_8 <= n48548;
       VREG_4_9 <= n48581;
       VREG_5_0 <= n48614;
       VREG_5_1 <= n48647;
       VREG_5_10 <= n48680;
       VREG_5_11 <= n48713;
       VREG_5_12 <= n48746;
       VREG_5_13 <= n48779;
       VREG_5_14 <= n48812;
       VREG_5_15 <= n48845;
       VREG_5_2 <= n48878;
       VREG_5_3 <= n48911;
       VREG_5_4 <= n48944;
       VREG_5_5 <= n48977;
       VREG_5_6 <= n49010;
       VREG_5_7 <= n49043;
       VREG_5_8 <= n49076;
       VREG_5_9 <= n49109;
       VREG_6_0 <= n49142;
       VREG_6_1 <= n49175;
       VREG_6_10 <= n49208;
       VREG_6_11 <= n49241;
       VREG_6_12 <= n49274;
       VREG_6_13 <= n49307;
       VREG_6_14 <= n49340;
       VREG_6_15 <= n49373;
       VREG_6_2 <= n49406;
       VREG_6_3 <= n49439;
       VREG_6_4 <= n49472;
       VREG_6_5 <= n49505;
       VREG_6_6 <= n49538;
       VREG_6_7 <= n49571;
       VREG_6_8 <= n49604;
       VREG_6_9 <= n49637;
       VREG_7_0 <= n49670;
       VREG_7_1 <= n49703;
       VREG_7_10 <= n49736;
       VREG_7_11 <= n49769;
       VREG_7_12 <= n49802;
       VREG_7_13 <= n49835;
       VREG_7_14 <= n49868;
       VREG_7_15 <= n49901;
       VREG_7_2 <= n49934;
       VREG_7_3 <= n49967;
       VREG_7_4 <= n50000;
       VREG_7_5 <= n50033;
       VREG_7_6 <= n50066;
       VREG_7_7 <= n50099;
       VREG_7_8 <= n50132;
       VREG_7_9 <= n50165;
       VREG_8_0 <= n50198;
       VREG_8_1 <= n50231;
       VREG_8_10 <= n50264;
       VREG_8_11 <= n50297;
       VREG_8_12 <= n50330;
       VREG_8_13 <= n50363;
       VREG_8_14 <= n50396;
       VREG_8_15 <= n50429;
       VREG_8_2 <= n50462;
       VREG_8_3 <= n50495;
       VREG_8_4 <= n50528;
       VREG_8_5 <= n50561;
       VREG_8_6 <= n50594;
       VREG_8_7 <= n50627;
       VREG_8_8 <= n50660;
       VREG_8_9 <= n50693;
       VREG_9_0 <= n50726;
       VREG_9_1 <= n50759;
       VREG_9_10 <= n50792;
       VREG_9_11 <= n50825;
       VREG_9_12 <= n50858;
       VREG_9_13 <= n50891;
       VREG_9_14 <= n50924;
       VREG_9_15 <= n50957;
       VREG_9_2 <= n50990;
       VREG_9_3 <= n51023;
       VREG_9_4 <= n51056;
       VREG_9_5 <= n51089;
       VREG_9_6 <= n51122;
       VREG_9_7 <= n51155;
       VREG_9_8 <= n51188;
       VREG_9_9 <= n51221;
       pc <= n51222;
   end
end
endmodule
